module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041;
  assign n17 = x0 & x8;
  assign n18 = x1 & x8;
  assign n19 = x0 & x9;
  assign n20 = n18 & n19;
  assign n21 = n18 | n19;
  assign n22 = ~n20 & n21;
  assign n23 = x2 & x8;
  assign n24 = x1 & x9;
  assign n25 = n23 & n24;
  assign n26 = n23 | n24;
  assign n27 = ~n25 & n26;
  assign n28 = n20 & n27;
  assign n29 = n20 | n27;
  assign n30 = ~n28 & n29;
  assign n31 = x0 & x10;
  assign n32 = n30 & n31;
  assign n33 = n30 | n31;
  assign n34 = ~n32 & n33;
  assign n441 = n20 | n25;
  assign n442 = (n25 & n27) | (n25 & n441) | (n27 & n441);
  assign n36 = x3 & x8;
  assign n37 = x2 & x9;
  assign n38 = n36 & n37;
  assign n39 = n36 | n37;
  assign n40 = ~n38 & n39;
  assign n41 = n442 & n40;
  assign n42 = n442 | n40;
  assign n43 = ~n41 & n42;
  assign n44 = x1 & x10;
  assign n45 = n43 & n44;
  assign n46 = n43 | n44;
  assign n47 = ~n45 & n46;
  assign n48 = n32 & n47;
  assign n49 = n32 | n47;
  assign n50 = ~n48 & n49;
  assign n51 = x0 & x11;
  assign n52 = n50 & n51;
  assign n53 = n50 | n51;
  assign n54 = ~n52 & n53;
  assign n443 = n32 | n45;
  assign n444 = (n45 & n47) | (n45 & n443) | (n47 & n443);
  assign n445 = n38 | n40;
  assign n446 = (n38 & n442) | (n38 & n445) | (n442 & n445);
  assign n57 = x4 & x8;
  assign n58 = x3 & x9;
  assign n59 = n57 & n58;
  assign n60 = n57 | n58;
  assign n61 = ~n59 & n60;
  assign n62 = n446 & n61;
  assign n63 = n446 | n61;
  assign n64 = ~n62 & n63;
  assign n65 = x2 & x10;
  assign n66 = n64 & n65;
  assign n67 = n64 | n65;
  assign n68 = ~n66 & n67;
  assign n69 = n444 & n68;
  assign n70 = n444 | n68;
  assign n71 = ~n69 & n70;
  assign n72 = x1 & x11;
  assign n73 = n71 & n72;
  assign n74 = n71 | n72;
  assign n75 = ~n73 & n74;
  assign n76 = n52 & n75;
  assign n77 = n52 | n75;
  assign n78 = ~n76 & n77;
  assign n79 = x0 & x12;
  assign n80 = n78 & n79;
  assign n81 = n78 | n79;
  assign n82 = ~n80 & n81;
  assign n447 = n52 | n73;
  assign n448 = (n73 & n75) | (n73 & n447) | (n75 & n447);
  assign n86 = x5 & x8;
  assign n87 = x4 & x9;
  assign n88 = n86 & n87;
  assign n89 = n86 | n87;
  assign n90 = ~n88 & n89;
  assign n449 = n59 | n61;
  assign n451 = n90 & n449;
  assign n452 = n59 & n90;
  assign n453 = (n446 & n451) | (n446 & n452) | (n451 & n452);
  assign n454 = n90 | n449;
  assign n455 = n59 | n90;
  assign n456 = (n446 & n454) | (n446 & n455) | (n454 & n455);
  assign n93 = ~n453 & n456;
  assign n94 = x3 & x10;
  assign n95 = n93 & n94;
  assign n96 = n93 | n94;
  assign n97 = ~n95 & n96;
  assign n457 = n66 & n97;
  assign n458 = (n69 & n97) | (n69 & n457) | (n97 & n457);
  assign n459 = n66 | n97;
  assign n460 = n69 | n459;
  assign n100 = ~n458 & n460;
  assign n101 = x2 & x11;
  assign n102 = n100 & n101;
  assign n103 = n100 | n101;
  assign n104 = ~n102 & n103;
  assign n105 = n448 & n104;
  assign n106 = n448 | n104;
  assign n107 = ~n105 & n106;
  assign n108 = x1 & x12;
  assign n109 = n107 & n108;
  assign n110 = n107 | n108;
  assign n111 = ~n109 & n110;
  assign n112 = n80 & n111;
  assign n113 = n80 | n111;
  assign n114 = ~n112 & n113;
  assign n115 = x0 & x13;
  assign n116 = n114 & n115;
  assign n117 = n114 | n115;
  assign n118 = ~n116 & n117;
  assign n461 = n80 | n109;
  assign n462 = (n109 & n111) | (n109 & n461) | (n111 & n461);
  assign n120 = n102 | n105;
  assign n123 = x6 & x8;
  assign n124 = x5 & x9;
  assign n125 = n123 & n124;
  assign n126 = n123 | n124;
  assign n127 = ~n125 & n126;
  assign n463 = n88 & n127;
  assign n464 = (n127 & n453) | (n127 & n463) | (n453 & n463);
  assign n465 = n88 | n127;
  assign n466 = n453 | n465;
  assign n130 = ~n464 & n466;
  assign n131 = x4 & x10;
  assign n132 = n130 & n131;
  assign n133 = n130 | n131;
  assign n134 = ~n132 & n133;
  assign n467 = n95 & n134;
  assign n468 = (n134 & n458) | (n134 & n467) | (n458 & n467);
  assign n469 = n95 | n134;
  assign n470 = n458 | n469;
  assign n137 = ~n468 & n470;
  assign n138 = x3 & x11;
  assign n139 = n137 & n138;
  assign n140 = n137 | n138;
  assign n141 = ~n139 & n140;
  assign n142 = n120 & n141;
  assign n143 = n120 | n141;
  assign n144 = ~n142 & n143;
  assign n145 = x2 & x12;
  assign n146 = n144 & n145;
  assign n147 = n144 | n145;
  assign n148 = ~n146 & n147;
  assign n149 = n462 & n148;
  assign n150 = n462 | n148;
  assign n151 = ~n149 & n150;
  assign n152 = x1 & x13;
  assign n153 = n151 & n152;
  assign n154 = n151 | n152;
  assign n155 = ~n153 & n154;
  assign n156 = n116 & n155;
  assign n157 = n116 | n155;
  assign n158 = ~n156 & n157;
  assign n159 = x0 & x14;
  assign n160 = n158 & n159;
  assign n161 = n158 | n159;
  assign n162 = ~n160 & n161;
  assign n724 = n115 | n152;
  assign n725 = (n114 & n152) | (n114 & n724) | (n152 & n724);
  assign n598 = (n116 & n151) | (n116 & n725) | (n151 & n725);
  assign n472 = (n153 & n155) | (n153 & n598) | (n155 & n598);
  assign n473 = n146 | n462;
  assign n474 = (n146 & n148) | (n146 & n473) | (n148 & n473);
  assign n475 = n139 | n141;
  assign n476 = (n120 & n139) | (n120 & n475) | (n139 & n475);
  assign n168 = x7 & x8;
  assign n169 = x6 & x9;
  assign n170 = n168 & n169;
  assign n171 = n168 | n169;
  assign n172 = ~n170 & n171;
  assign n599 = n88 | n125;
  assign n600 = (n125 & n127) | (n125 & n599) | (n127 & n599);
  assign n480 = n172 & n600;
  assign n478 = n125 | n127;
  assign n481 = n172 & n478;
  assign n482 = (n453 & n480) | (n453 & n481) | (n480 & n481);
  assign n483 = n172 | n600;
  assign n484 = n172 | n478;
  assign n485 = (n453 & n483) | (n453 & n484) | (n483 & n484);
  assign n175 = ~n482 & n485;
  assign n176 = x5 & x10;
  assign n177 = n175 & n176;
  assign n178 = n175 | n176;
  assign n179 = ~n177 & n178;
  assign n486 = n132 & n179;
  assign n487 = (n179 & n468) | (n179 & n486) | (n468 & n486);
  assign n488 = n132 | n179;
  assign n489 = n468 | n488;
  assign n182 = ~n487 & n489;
  assign n183 = x4 & x11;
  assign n184 = n182 & n183;
  assign n185 = n182 | n183;
  assign n186 = ~n184 & n185;
  assign n187 = n476 & n186;
  assign n188 = n476 | n186;
  assign n189 = ~n187 & n188;
  assign n190 = x3 & x12;
  assign n191 = n189 & n190;
  assign n192 = n189 | n190;
  assign n193 = ~n191 & n192;
  assign n194 = n474 & n193;
  assign n195 = n474 | n193;
  assign n196 = ~n194 & n195;
  assign n197 = x2 & x13;
  assign n198 = n196 & n197;
  assign n199 = n196 | n197;
  assign n200 = ~n198 & n199;
  assign n201 = n472 & n200;
  assign n202 = n472 | n200;
  assign n203 = ~n201 & n202;
  assign n204 = x1 & x14;
  assign n205 = n203 & n204;
  assign n206 = n203 | n204;
  assign n207 = ~n205 & n206;
  assign n208 = n160 & n207;
  assign n209 = n160 | n207;
  assign n210 = ~n208 & n209;
  assign n211 = x0 & x15;
  assign n212 = n210 & n211;
  assign n213 = n210 | n211;
  assign n214 = ~n212 & n213;
  assign n490 = n160 | n205;
  assign n491 = (n205 & n207) | (n205 & n490) | (n207 & n490);
  assign n216 = n198 | n201;
  assign n217 = n191 | n194;
  assign n492 = n184 | n186;
  assign n493 = (n184 & n476) | (n184 & n492) | (n476 & n492);
  assign n221 = x7 & x9;
  assign n497 = n170 & n221;
  assign n726 = (n172 & n221) | (n172 & n497) | (n221 & n497);
  assign n728 = (n478 & n726) | (n478 & n497) | (n726 & n497);
  assign n729 = (n600 & n726) | (n600 & n497) | (n726 & n497);
  assign n605 = (n453 & n728) | (n453 & n729) | (n728 & n729);
  assign n499 = n170 | n221;
  assign n730 = n172 | n499;
  assign n731 = (n478 & n499) | (n478 & n730) | (n499 & n730);
  assign n732 = (n499 & n600) | (n499 & n730) | (n600 & n730);
  assign n608 = (n453 & n731) | (n453 & n732) | (n731 & n732);
  assign n224 = ~n605 & n608;
  assign n225 = x6 & x10;
  assign n226 = n224 & n225;
  assign n227 = n224 | n225;
  assign n228 = ~n226 & n227;
  assign n495 = n177 | n179;
  assign n609 = n228 & n495;
  assign n601 = n132 | n177;
  assign n602 = (n177 & n179) | (n177 & n601) | (n179 & n601);
  assign n610 = n228 & n602;
  assign n611 = (n468 & n609) | (n468 & n610) | (n609 & n610);
  assign n612 = n228 | n495;
  assign n613 = n228 | n602;
  assign n614 = (n468 & n612) | (n468 & n613) | (n612 & n613);
  assign n231 = ~n611 & n614;
  assign n232 = x5 & x11;
  assign n233 = n231 & n232;
  assign n234 = n231 | n232;
  assign n235 = ~n233 & n234;
  assign n236 = n493 & n235;
  assign n237 = n493 | n235;
  assign n238 = ~n236 & n237;
  assign n239 = x4 & x12;
  assign n240 = n238 & n239;
  assign n241 = n238 | n239;
  assign n242 = ~n240 & n241;
  assign n243 = n217 & n242;
  assign n244 = n217 | n242;
  assign n245 = ~n243 & n244;
  assign n246 = x3 & x13;
  assign n247 = n245 & n246;
  assign n248 = n245 | n246;
  assign n249 = ~n247 & n248;
  assign n250 = n216 & n249;
  assign n251 = n216 | n249;
  assign n252 = ~n250 & n251;
  assign n253 = x2 & x14;
  assign n254 = n252 & n253;
  assign n255 = n252 | n253;
  assign n256 = ~n254 & n255;
  assign n257 = n491 & n256;
  assign n258 = n491 | n256;
  assign n259 = ~n257 & n258;
  assign n260 = x1 & x15;
  assign n261 = n259 & n260;
  assign n262 = n259 | n260;
  assign n263 = ~n261 & n262;
  assign n264 = n212 & n263;
  assign n265 = n212 | n263;
  assign n266 = ~n264 & n265;
  assign n733 = n211 | n260;
  assign n734 = (n210 & n260) | (n210 & n733) | (n260 & n733);
  assign n616 = (n212 & n259) | (n212 & n734) | (n259 & n734);
  assign n502 = (n261 & n263) | (n261 & n616) | (n263 & n616);
  assign n503 = n254 | n491;
  assign n504 = (n254 & n256) | (n254 & n503) | (n256 & n503);
  assign n269 = n247 | n250;
  assign n505 = n240 | n242;
  assign n506 = (n217 & n240) | (n217 & n505) | (n240 & n505);
  assign n273 = x7 & x10;
  assign n512 = n221 & n273;
  assign n617 = n170 & n512;
  assign n735 = (n172 & n512) | (n172 & n617) | (n512 & n617);
  assign n736 = n512 & n617;
  assign n737 = (n478 & n735) | (n478 & n736) | (n735 & n736);
  assign n738 = (n600 & n735) | (n600 & n736) | (n735 & n736);
  assign n620 = (n453 & n737) | (n453 & n738) | (n737 & n738);
  assign n515 = n221 | n273;
  assign n621 = (n170 & n273) | (n170 & n515) | (n273 & n515);
  assign n739 = (n172 & n515) | (n172 & n621) | (n515 & n621);
  assign n740 = n515 & n621;
  assign n741 = (n478 & n739) | (n478 & n740) | (n739 & n740);
  assign n742 = (n600 & n739) | (n600 & n740) | (n739 & n740);
  assign n624 = (n453 & n741) | (n453 & n742) | (n741 & n742);
  assign n276 = ~n620 & n624;
  assign n518 = n226 & n276;
  assign n625 = (n228 & n276) | (n228 & n518) | (n276 & n518);
  assign n626 = (n495 & n518) | (n495 & n625) | (n518 & n625);
  assign n627 = (n518 & n602) | (n518 & n625) | (n602 & n625);
  assign n628 = (n468 & n626) | (n468 & n627) | (n626 & n627);
  assign n521 = n226 | n276;
  assign n629 = n228 | n521;
  assign n630 = (n495 & n521) | (n495 & n629) | (n521 & n629);
  assign n631 = (n521 & n602) | (n521 & n629) | (n602 & n629);
  assign n632 = (n468 & n630) | (n468 & n631) | (n630 & n631);
  assign n279 = ~n628 & n632;
  assign n280 = x6 & x11;
  assign n281 = n279 & n280;
  assign n282 = n279 | n280;
  assign n283 = ~n281 & n282;
  assign n507 = n233 | n235;
  assign n633 = n283 & n507;
  assign n634 = n233 & n283;
  assign n635 = (n493 & n633) | (n493 & n634) | (n633 & n634);
  assign n636 = n283 | n507;
  assign n637 = n233 | n283;
  assign n638 = (n493 & n636) | (n493 & n637) | (n636 & n637);
  assign n286 = ~n635 & n638;
  assign n287 = x5 & x12;
  assign n288 = n286 & n287;
  assign n289 = n286 | n287;
  assign n290 = ~n288 & n289;
  assign n291 = n506 & n290;
  assign n292 = n506 | n290;
  assign n293 = ~n291 & n292;
  assign n294 = x4 & x13;
  assign n295 = n293 & n294;
  assign n296 = n293 | n294;
  assign n297 = ~n295 & n296;
  assign n298 = n269 & n297;
  assign n299 = n269 | n297;
  assign n300 = ~n298 & n299;
  assign n301 = x3 & x14;
  assign n302 = n300 & n301;
  assign n303 = n300 | n301;
  assign n304 = ~n302 & n303;
  assign n305 = n504 & n304;
  assign n306 = n504 | n304;
  assign n307 = ~n305 & n306;
  assign n308 = x2 & x15;
  assign n309 = n307 & n308;
  assign n310 = n307 | n308;
  assign n311 = ~n309 & n310;
  assign n312 = n502 & n311;
  assign n313 = n502 | n311;
  assign n314 = ~n312 & n313;
  assign n523 = n309 | n502;
  assign n524 = (n309 & n311) | (n309 & n523) | (n311 & n523);
  assign n525 = n302 | n504;
  assign n526 = (n302 & n304) | (n302 & n525) | (n304 & n525);
  assign n527 = n295 | n297;
  assign n528 = (n269 & n295) | (n269 & n527) | (n295 & n527);
  assign n321 = x7 & x11;
  assign n743 = n321 & n738;
  assign n744 = n321 & n737;
  assign n745 = (n453 & n743) | (n453 & n744) | (n743 & n744);
  assign n534 = (n321 & n628) | (n321 & n745) | (n628 & n745);
  assign n746 = n321 | n738;
  assign n747 = n321 | n737;
  assign n748 = (n453 & n746) | (n453 & n747) | (n746 & n747);
  assign n536 = n628 | n748;
  assign n324 = ~n534 & n536;
  assign n538 = n281 & n324;
  assign n639 = (n283 & n324) | (n283 & n538) | (n324 & n538);
  assign n640 = (n507 & n538) | (n507 & n639) | (n538 & n639);
  assign n641 = (n233 & n538) | (n233 & n639) | (n538 & n639);
  assign n642 = (n493 & n640) | (n493 & n641) | (n640 & n641);
  assign n541 = n281 | n324;
  assign n643 = n283 | n541;
  assign n644 = (n507 & n541) | (n507 & n643) | (n541 & n643);
  assign n645 = (n233 & n541) | (n233 & n643) | (n541 & n643);
  assign n646 = (n493 & n644) | (n493 & n645) | (n644 & n645);
  assign n327 = ~n642 & n646;
  assign n328 = x6 & x12;
  assign n329 = n327 & n328;
  assign n330 = n327 | n328;
  assign n331 = ~n329 & n330;
  assign n529 = n288 | n290;
  assign n647 = n331 & n529;
  assign n648 = n288 & n331;
  assign n649 = (n506 & n647) | (n506 & n648) | (n647 & n648);
  assign n650 = n331 | n529;
  assign n651 = n288 | n331;
  assign n652 = (n506 & n650) | (n506 & n651) | (n650 & n651);
  assign n334 = ~n649 & n652;
  assign n335 = x5 & x13;
  assign n336 = n334 & n335;
  assign n337 = n334 | n335;
  assign n338 = ~n336 & n337;
  assign n339 = n528 & n338;
  assign n340 = n528 | n338;
  assign n341 = ~n339 & n340;
  assign n342 = x4 & x14;
  assign n343 = n341 & n342;
  assign n344 = n341 | n342;
  assign n345 = ~n343 & n344;
  assign n346 = n526 & n345;
  assign n347 = n526 | n345;
  assign n348 = ~n346 & n347;
  assign n349 = x3 & x15;
  assign n350 = n348 & n349;
  assign n351 = n348 | n349;
  assign n352 = ~n350 & n351;
  assign n353 = n524 & n352;
  assign n354 = n524 | n352;
  assign n355 = ~n353 & n354;
  assign n356 = n350 | n353;
  assign n361 = x7 & x12;
  assign n653 = n361 & n745;
  assign n654 = n321 & n361;
  assign n655 = (n628 & n653) | (n628 & n654) | (n653 & n654);
  assign n548 = (n361 & n642) | (n361 & n655) | (n642 & n655);
  assign n656 = n361 | n745;
  assign n657 = n321 | n361;
  assign n658 = (n628 & n656) | (n628 & n657) | (n656 & n657);
  assign n550 = n642 | n658;
  assign n364 = ~n548 & n550;
  assign n552 = n329 & n364;
  assign n659 = (n331 & n364) | (n331 & n552) | (n364 & n552);
  assign n660 = (n529 & n552) | (n529 & n659) | (n552 & n659);
  assign n661 = (n288 & n552) | (n288 & n659) | (n552 & n659);
  assign n662 = (n506 & n660) | (n506 & n661) | (n660 & n661);
  assign n555 = n329 | n364;
  assign n663 = n331 | n555;
  assign n664 = (n529 & n555) | (n529 & n663) | (n555 & n663);
  assign n665 = (n288 & n555) | (n288 & n663) | (n555 & n663);
  assign n666 = (n506 & n664) | (n506 & n665) | (n664 & n665);
  assign n367 = ~n662 & n666;
  assign n368 = x6 & x13;
  assign n369 = n367 & n368;
  assign n370 = n367 | n368;
  assign n371 = ~n369 & n370;
  assign n543 = n336 | n338;
  assign n667 = n371 & n543;
  assign n668 = n336 & n371;
  assign n669 = (n528 & n667) | (n528 & n668) | (n667 & n668);
  assign n670 = n371 | n543;
  assign n671 = n336 | n371;
  assign n672 = (n528 & n670) | (n528 & n671) | (n670 & n671);
  assign n374 = ~n669 & n672;
  assign n375 = x5 & x14;
  assign n376 = n374 & n375;
  assign n377 = n374 | n375;
  assign n378 = ~n376 & n377;
  assign n673 = n343 & n378;
  assign n674 = (n346 & n378) | (n346 & n673) | (n378 & n673);
  assign n675 = n343 | n378;
  assign n676 = n346 | n675;
  assign n381 = ~n674 & n676;
  assign n382 = x4 & x15;
  assign n383 = n381 & n382;
  assign n384 = n381 | n382;
  assign n385 = ~n383 & n384;
  assign n386 = n356 & n385;
  assign n387 = n356 | n385;
  assign n388 = ~n386 & n387;
  assign n677 = n383 | n385;
  assign n678 = (n356 & n383) | (n356 & n677) | (n383 & n677);
  assign n357 = n343 | n346;
  assign n393 = x7 & x13;
  assign n680 = n361 & n393;
  assign n2671 = n680 & n745;
  assign n750 = n393 & n654;
  assign n751 = (n628 & n2671) | (n628 & n750) | (n2671 & n750);
  assign n681 = (n642 & n751) | (n642 & n680) | (n751 & n680);
  assign n562 = (n393 & n662) | (n393 & n681) | (n662 & n681);
  assign n683 = n361 | n393;
  assign n2672 = (n393 & n683) | (n393 & n745) | (n683 & n745);
  assign n753 = n393 | n654;
  assign n754 = (n628 & n2672) | (n628 & n753) | (n2672 & n753);
  assign n684 = (n642 & n754) | (n642 & n683) | (n754 & n683);
  assign n564 = n662 | n684;
  assign n396 = ~n562 & n564;
  assign n566 = n369 & n396;
  assign n685 = (n371 & n396) | (n371 & n566) | (n396 & n566);
  assign n686 = (n543 & n566) | (n543 & n685) | (n566 & n685);
  assign n687 = (n336 & n566) | (n336 & n685) | (n566 & n685);
  assign n688 = (n528 & n686) | (n528 & n687) | (n686 & n687);
  assign n569 = n369 | n396;
  assign n689 = n371 | n569;
  assign n690 = (n543 & n569) | (n543 & n689) | (n569 & n689);
  assign n691 = (n336 & n569) | (n336 & n689) | (n569 & n689);
  assign n692 = (n528 & n690) | (n528 & n691) | (n690 & n691);
  assign n399 = ~n688 & n692;
  assign n400 = x6 & x14;
  assign n401 = n399 & n400;
  assign n402 = n399 | n400;
  assign n403 = ~n401 & n402;
  assign n557 = n376 | n378;
  assign n693 = n403 & n557;
  assign n694 = n376 & n403;
  assign n695 = (n357 & n693) | (n357 & n694) | (n693 & n694);
  assign n696 = n403 | n557;
  assign n697 = n376 | n403;
  assign n698 = (n357 & n696) | (n357 & n697) | (n696 & n697);
  assign n406 = ~n695 & n698;
  assign n407 = x5 & x15;
  assign n408 = n406 & n407;
  assign n409 = n406 | n407;
  assign n410 = ~n408 & n409;
  assign n411 = n678 & n410;
  assign n412 = n678 | n410;
  assign n413 = ~n411 & n412;
  assign n571 = n408 | n410;
  assign n572 = (n678 & n408) | (n678 & n571) | (n408 & n571);
  assign n417 = x7 & x14;
  assign n756 = n417 & n680;
  assign n3429 = n745 & n756;
  assign n700 = n393 & n417;
  assign n3430 = n654 & n700;
  assign n2675 = (n628 & n3429) | (n628 & n3430) | (n3429 & n3430);
  assign n757 = (n642 & n2675) | (n642 & n756) | (n2675 & n756);
  assign n701 = (n662 & n757) | (n662 & n700) | (n757 & n700);
  assign n576 = (n417 & n688) | (n417 & n701) | (n688 & n701);
  assign n759 = n417 | n680;
  assign n3431 = (n417 & n745) | (n417 & n759) | (n745 & n759);
  assign n703 = n393 | n417;
  assign n3432 = (n417 & n654) | (n417 & n703) | (n654 & n703);
  assign n2678 = (n628 & n3431) | (n628 & n3432) | (n3431 & n3432);
  assign n760 = (n642 & n2678) | (n642 & n759) | (n2678 & n759);
  assign n704 = (n662 & n760) | (n662 & n703) | (n760 & n703);
  assign n578 = n688 | n704;
  assign n420 = ~n576 & n578;
  assign n580 = n401 & n420;
  assign n705 = (n403 & n420) | (n403 & n580) | (n420 & n580);
  assign n706 = (n557 & n580) | (n557 & n705) | (n580 & n705);
  assign n707 = (n376 & n580) | (n376 & n705) | (n580 & n705);
  assign n708 = (n357 & n706) | (n357 & n707) | (n706 & n707);
  assign n583 = n401 | n420;
  assign n709 = n403 | n583;
  assign n710 = (n557 & n583) | (n557 & n709) | (n583 & n709);
  assign n711 = (n376 & n583) | (n376 & n709) | (n583 & n709);
  assign n712 = (n357 & n710) | (n357 & n711) | (n710 & n711);
  assign n423 = ~n708 & n712;
  assign n424 = x6 & x15;
  assign n425 = n423 & n424;
  assign n426 = n423 | n424;
  assign n427 = ~n425 & n426;
  assign n428 = n572 & n427;
  assign n429 = n572 | n427;
  assign n430 = ~n428 & n429;
  assign n433 = x7 & x15;
  assign n2680 = n433 & n756;
  assign n3895 = n745 & n2680;
  assign n3434 = n433 & n3430;
  assign n3435 = (n628 & n3895) | (n628 & n3434) | (n3895 & n3434);
  assign n714 = n417 & n433;
  assign n3436 = n680 & n714;
  assign n2681 = (n642 & n3435) | (n642 & n3436) | (n3435 & n3436);
  assign n762 = n433 & n700;
  assign n763 = (n662 & n2681) | (n662 & n762) | (n2681 & n762);
  assign n715 = (n688 & n763) | (n688 & n714) | (n763 & n714);
  assign n588 = (n433 & n708) | (n433 & n715) | (n708 & n715);
  assign n2683 = n433 | n756;
  assign n3896 = (n433 & n745) | (n433 & n2683) | (n745 & n2683);
  assign n3438 = n433 | n3430;
  assign n3439 = (n628 & n3896) | (n628 & n3438) | (n3896 & n3438);
  assign n717 = n417 | n433;
  assign n3440 = (n433 & n680) | (n433 & n717) | (n680 & n717);
  assign n2684 = (n642 & n3439) | (n642 & n3440) | (n3439 & n3440);
  assign n765 = n433 | n700;
  assign n766 = (n662 & n2684) | (n662 & n765) | (n2684 & n765);
  assign n718 = (n688 & n766) | (n688 & n717) | (n766 & n717);
  assign n590 = n708 | n718;
  assign n436 = ~n588 & n590;
  assign n592 = n425 & n436;
  assign n719 = (n427 & n436) | (n427 & n592) | (n436 & n592);
  assign n593 = (n572 & n719) | (n572 & n592) | (n719 & n592);
  assign n595 = n425 | n436;
  assign n720 = n427 | n595;
  assign n596 = (n572 & n720) | (n572 & n595) | (n720 & n595);
  assign n439 = ~n593 & n596;
  assign n721 = n588 | n719;
  assign n722 = n588 | n592;
  assign n723 = (n572 & n721) | (n572 & n722) | (n721 & n722);
  assign n799 = x16 & x32;
  assign n800 = x17 & x32;
  assign n801 = x16 & x33;
  assign n802 = n800 & n801;
  assign n803 = n800 | n801;
  assign n804 = ~n802 & n803;
  assign n805 = x18 & x32;
  assign n806 = x17 & x33;
  assign n807 = n805 & n806;
  assign n808 = n805 | n806;
  assign n809 = ~n807 & n808;
  assign n810 = n802 & n809;
  assign n811 = n802 | n809;
  assign n812 = ~n810 & n811;
  assign n813 = x16 & x34;
  assign n814 = n812 & n813;
  assign n815 = n812 | n813;
  assign n816 = ~n814 & n815;
  assign n2685 = n802 | n807;
  assign n2686 = (n807 & n809) | (n807 & n2685) | (n809 & n2685);
  assign n818 = x19 & x32;
  assign n819 = x18 & x33;
  assign n820 = n818 & n819;
  assign n821 = n818 | n819;
  assign n822 = ~n820 & n821;
  assign n823 = n2686 & n822;
  assign n824 = n2686 | n822;
  assign n825 = ~n823 & n824;
  assign n826 = x17 & x34;
  assign n827 = n825 & n826;
  assign n828 = n825 | n826;
  assign n829 = ~n827 & n828;
  assign n830 = n814 & n829;
  assign n831 = n814 | n829;
  assign n832 = ~n830 & n831;
  assign n833 = x16 & x35;
  assign n834 = n832 & n833;
  assign n835 = n832 | n833;
  assign n836 = ~n834 & n835;
  assign n2687 = n814 | n827;
  assign n2688 = (n827 & n829) | (n827 & n2687) | (n829 & n2687);
  assign n2689 = n820 | n822;
  assign n2690 = (n820 & n2686) | (n820 & n2689) | (n2686 & n2689);
  assign n839 = x20 & x32;
  assign n840 = x19 & x33;
  assign n841 = n839 & n840;
  assign n842 = n839 | n840;
  assign n843 = ~n841 & n842;
  assign n844 = n2690 & n843;
  assign n845 = n2690 | n843;
  assign n846 = ~n844 & n845;
  assign n847 = x18 & x34;
  assign n848 = n846 & n847;
  assign n849 = n846 | n847;
  assign n850 = ~n848 & n849;
  assign n851 = n2688 & n850;
  assign n852 = n2688 | n850;
  assign n853 = ~n851 & n852;
  assign n854 = x17 & x35;
  assign n855 = n853 & n854;
  assign n856 = n853 | n854;
  assign n857 = ~n855 & n856;
  assign n858 = n834 & n857;
  assign n859 = n834 | n857;
  assign n860 = ~n858 & n859;
  assign n861 = x16 & x36;
  assign n862 = n860 & n861;
  assign n863 = n860 | n861;
  assign n864 = ~n862 & n863;
  assign n2691 = n834 | n855;
  assign n2692 = (n855 & n857) | (n855 & n2691) | (n857 & n2691);
  assign n868 = x21 & x32;
  assign n869 = x20 & x33;
  assign n870 = n868 & n869;
  assign n871 = n868 | n869;
  assign n872 = ~n870 & n871;
  assign n2693 = n841 | n843;
  assign n2695 = n872 & n2693;
  assign n2696 = n841 & n872;
  assign n2697 = (n2690 & n2695) | (n2690 & n2696) | (n2695 & n2696);
  assign n2698 = n872 | n2693;
  assign n2699 = n841 | n872;
  assign n2700 = (n2690 & n2698) | (n2690 & n2699) | (n2698 & n2699);
  assign n875 = ~n2697 & n2700;
  assign n876 = x19 & x34;
  assign n877 = n875 & n876;
  assign n878 = n875 | n876;
  assign n879 = ~n877 & n878;
  assign n2701 = n848 & n879;
  assign n2702 = (n851 & n879) | (n851 & n2701) | (n879 & n2701);
  assign n2703 = n848 | n879;
  assign n2704 = n851 | n2703;
  assign n882 = ~n2702 & n2704;
  assign n883 = x18 & x35;
  assign n884 = n882 & n883;
  assign n885 = n882 | n883;
  assign n886 = ~n884 & n885;
  assign n887 = n2692 & n886;
  assign n888 = n2692 | n886;
  assign n889 = ~n887 & n888;
  assign n890 = x17 & x36;
  assign n891 = n889 & n890;
  assign n892 = n889 | n890;
  assign n893 = ~n891 & n892;
  assign n894 = n862 & n893;
  assign n895 = n862 | n893;
  assign n896 = ~n894 & n895;
  assign n897 = x16 & x37;
  assign n898 = n896 & n897;
  assign n899 = n896 | n897;
  assign n900 = ~n898 & n899;
  assign n2705 = n862 | n891;
  assign n2706 = (n891 & n893) | (n891 & n2705) | (n893 & n2705);
  assign n902 = n884 | n887;
  assign n905 = x22 & x32;
  assign n906 = x21 & x33;
  assign n907 = n905 & n906;
  assign n908 = n905 | n906;
  assign n909 = ~n907 & n908;
  assign n2707 = n870 & n909;
  assign n2708 = (n909 & n2697) | (n909 & n2707) | (n2697 & n2707);
  assign n2709 = n870 | n909;
  assign n2710 = n2697 | n2709;
  assign n912 = ~n2708 & n2710;
  assign n913 = x20 & x34;
  assign n914 = n912 & n913;
  assign n915 = n912 | n913;
  assign n916 = ~n914 & n915;
  assign n2711 = n877 & n916;
  assign n2712 = (n916 & n2702) | (n916 & n2711) | (n2702 & n2711);
  assign n2713 = n877 | n916;
  assign n2714 = n2702 | n2713;
  assign n919 = ~n2712 & n2714;
  assign n920 = x19 & x35;
  assign n921 = n919 & n920;
  assign n922 = n919 | n920;
  assign n923 = ~n921 & n922;
  assign n924 = n902 & n923;
  assign n925 = n902 | n923;
  assign n926 = ~n924 & n925;
  assign n927 = x18 & x36;
  assign n928 = n926 & n927;
  assign n929 = n926 | n927;
  assign n930 = ~n928 & n929;
  assign n931 = n2706 & n930;
  assign n932 = n2706 | n930;
  assign n933 = ~n931 & n932;
  assign n934 = x17 & x37;
  assign n935 = n933 & n934;
  assign n936 = n933 | n934;
  assign n937 = ~n935 & n936;
  assign n938 = n898 & n937;
  assign n939 = n898 | n937;
  assign n940 = ~n938 & n939;
  assign n941 = x16 & x38;
  assign n942 = n940 & n941;
  assign n943 = n940 | n941;
  assign n944 = ~n942 & n943;
  assign n3897 = n897 | n934;
  assign n3898 = (n896 & n934) | (n896 & n3897) | (n934 & n3897);
  assign n3442 = (n898 & n933) | (n898 & n3898) | (n933 & n3898);
  assign n2716 = (n935 & n937) | (n935 & n3442) | (n937 & n3442);
  assign n2717 = n928 | n2706;
  assign n2718 = (n928 & n930) | (n928 & n2717) | (n930 & n2717);
  assign n2719 = n921 | n923;
  assign n2720 = (n902 & n921) | (n902 & n2719) | (n921 & n2719);
  assign n950 = x23 & x32;
  assign n951 = x22 & x33;
  assign n952 = n950 & n951;
  assign n953 = n950 | n951;
  assign n954 = ~n952 & n953;
  assign n3443 = n870 | n907;
  assign n3444 = (n907 & n909) | (n907 & n3443) | (n909 & n3443);
  assign n2724 = n954 & n3444;
  assign n2722 = n907 | n909;
  assign n2725 = n954 & n2722;
  assign n2726 = (n2697 & n2724) | (n2697 & n2725) | (n2724 & n2725);
  assign n2727 = n954 | n3444;
  assign n2728 = n954 | n2722;
  assign n2729 = (n2697 & n2727) | (n2697 & n2728) | (n2727 & n2728);
  assign n957 = ~n2726 & n2729;
  assign n958 = x21 & x34;
  assign n959 = n957 & n958;
  assign n960 = n957 | n958;
  assign n961 = ~n959 & n960;
  assign n2730 = n914 & n961;
  assign n2731 = (n961 & n2712) | (n961 & n2730) | (n2712 & n2730);
  assign n2732 = n914 | n961;
  assign n2733 = n2712 | n2732;
  assign n964 = ~n2731 & n2733;
  assign n965 = x20 & x35;
  assign n966 = n964 & n965;
  assign n967 = n964 | n965;
  assign n968 = ~n966 & n967;
  assign n969 = n2720 & n968;
  assign n970 = n2720 | n968;
  assign n971 = ~n969 & n970;
  assign n972 = x19 & x36;
  assign n973 = n971 & n972;
  assign n974 = n971 | n972;
  assign n975 = ~n973 & n974;
  assign n976 = n2718 & n975;
  assign n977 = n2718 | n975;
  assign n978 = ~n976 & n977;
  assign n979 = x18 & x37;
  assign n980 = n978 & n979;
  assign n981 = n978 | n979;
  assign n982 = ~n980 & n981;
  assign n983 = n2716 & n982;
  assign n984 = n2716 | n982;
  assign n985 = ~n983 & n984;
  assign n986 = x17 & x38;
  assign n987 = n985 & n986;
  assign n988 = n985 | n986;
  assign n989 = ~n987 & n988;
  assign n990 = n942 & n989;
  assign n991 = n942 | n989;
  assign n992 = ~n990 & n991;
  assign n993 = x16 & x39;
  assign n994 = n992 & n993;
  assign n995 = n992 | n993;
  assign n996 = ~n994 & n995;
  assign n2734 = n942 | n987;
  assign n2735 = (n987 & n989) | (n987 & n2734) | (n989 & n2734);
  assign n998 = n980 | n983;
  assign n999 = n973 | n976;
  assign n2736 = n966 | n968;
  assign n2737 = (n966 & n2720) | (n966 & n2736) | (n2720 & n2736);
  assign n1003 = x24 & x32;
  assign n1004 = x23 & x33;
  assign n1005 = n1003 & n1004;
  assign n1006 = n1003 | n1004;
  assign n1007 = ~n1005 & n1006;
  assign n2741 = n952 & n1007;
  assign n3447 = (n1007 & n2725) | (n1007 & n2741) | (n2725 & n2741);
  assign n3448 = (n1007 & n2724) | (n1007 & n2741) | (n2724 & n2741);
  assign n3449 = (n2697 & n3447) | (n2697 & n3448) | (n3447 & n3448);
  assign n2743 = n952 | n1007;
  assign n3450 = n2725 | n2743;
  assign n3451 = n2724 | n2743;
  assign n3452 = (n2697 & n3450) | (n2697 & n3451) | (n3450 & n3451);
  assign n1010 = ~n3449 & n3452;
  assign n1011 = x22 & x34;
  assign n1012 = n1010 & n1011;
  assign n1013 = n1010 | n1011;
  assign n1014 = ~n1012 & n1013;
  assign n2739 = n959 | n961;
  assign n3453 = n1014 & n2739;
  assign n3445 = n914 | n959;
  assign n3446 = (n959 & n961) | (n959 & n3445) | (n961 & n3445);
  assign n3454 = n1014 & n3446;
  assign n3455 = (n2712 & n3453) | (n2712 & n3454) | (n3453 & n3454);
  assign n3456 = n1014 | n2739;
  assign n3457 = n1014 | n3446;
  assign n3458 = (n2712 & n3456) | (n2712 & n3457) | (n3456 & n3457);
  assign n1017 = ~n3455 & n3458;
  assign n1018 = x21 & x35;
  assign n1019 = n1017 & n1018;
  assign n1020 = n1017 | n1018;
  assign n1021 = ~n1019 & n1020;
  assign n1022 = n2737 & n1021;
  assign n1023 = n2737 | n1021;
  assign n1024 = ~n1022 & n1023;
  assign n1025 = x20 & x36;
  assign n1026 = n1024 & n1025;
  assign n1027 = n1024 | n1025;
  assign n1028 = ~n1026 & n1027;
  assign n1029 = n999 & n1028;
  assign n1030 = n999 | n1028;
  assign n1031 = ~n1029 & n1030;
  assign n1032 = x19 & x37;
  assign n1033 = n1031 & n1032;
  assign n1034 = n1031 | n1032;
  assign n1035 = ~n1033 & n1034;
  assign n1036 = n998 & n1035;
  assign n1037 = n998 | n1035;
  assign n1038 = ~n1036 & n1037;
  assign n1039 = x18 & x38;
  assign n1040 = n1038 & n1039;
  assign n1041 = n1038 | n1039;
  assign n1042 = ~n1040 & n1041;
  assign n1043 = n2735 & n1042;
  assign n1044 = n2735 | n1042;
  assign n1045 = ~n1043 & n1044;
  assign n1046 = x17 & x39;
  assign n1047 = n1045 & n1046;
  assign n1048 = n1045 | n1046;
  assign n1049 = ~n1047 & n1048;
  assign n1050 = n994 & n1049;
  assign n1051 = n994 | n1049;
  assign n1052 = ~n1050 & n1051;
  assign n1053 = x16 & x40;
  assign n1054 = n1052 & n1053;
  assign n1055 = n1052 | n1053;
  assign n1056 = ~n1054 & n1055;
  assign n3899 = n993 | n1046;
  assign n3900 = (n992 & n1046) | (n992 & n3899) | (n1046 & n3899);
  assign n3460 = (n994 & n1045) | (n994 & n3900) | (n1045 & n3900);
  assign n2746 = (n1047 & n1049) | (n1047 & n3460) | (n1049 & n3460);
  assign n2747 = n1040 | n2735;
  assign n2748 = (n1040 & n1042) | (n1040 & n2747) | (n1042 & n2747);
  assign n1059 = n1033 | n1036;
  assign n2749 = n1026 | n1028;
  assign n2750 = (n999 & n1026) | (n999 & n2749) | (n1026 & n2749);
  assign n2740 = (n2712 & n3446) | (n2712 & n2739) | (n3446 & n2739);
  assign n1064 = x25 & x32;
  assign n1065 = x24 & x33;
  assign n1066 = n1064 & n1065;
  assign n1067 = n1064 | n1065;
  assign n1068 = ~n1066 & n1067;
  assign n3461 = n952 | n1005;
  assign n3462 = (n1005 & n1007) | (n1005 & n3461) | (n1007 & n3461);
  assign n2758 = n1068 & n3462;
  assign n2756 = n1005 | n1007;
  assign n2759 = n1068 & n2756;
  assign n3463 = (n2725 & n2758) | (n2725 & n2759) | (n2758 & n2759);
  assign n3464 = (n2724 & n2758) | (n2724 & n2759) | (n2758 & n2759);
  assign n3465 = (n2697 & n3463) | (n2697 & n3464) | (n3463 & n3464);
  assign n2761 = n1068 | n3462;
  assign n2762 = n1068 | n2756;
  assign n3466 = (n2725 & n2761) | (n2725 & n2762) | (n2761 & n2762);
  assign n3467 = (n2724 & n2761) | (n2724 & n2762) | (n2761 & n2762);
  assign n3468 = (n2697 & n3466) | (n2697 & n3467) | (n3466 & n3467);
  assign n1071 = ~n3465 & n3468;
  assign n1072 = x23 & x34;
  assign n1073 = n1071 & n1072;
  assign n1074 = n1071 | n1072;
  assign n1075 = ~n1073 & n1074;
  assign n2753 = n1012 | n1014;
  assign n2764 = n1075 & n2753;
  assign n2765 = n1012 & n1075;
  assign n2766 = (n2740 & n2764) | (n2740 & n2765) | (n2764 & n2765);
  assign n2767 = n1075 | n2753;
  assign n2768 = n1012 | n1075;
  assign n2769 = (n2740 & n2767) | (n2740 & n2768) | (n2767 & n2768);
  assign n1078 = ~n2766 & n2769;
  assign n1079 = x22 & x35;
  assign n1080 = n1078 & n1079;
  assign n1081 = n1078 | n1079;
  assign n1082 = ~n1080 & n1081;
  assign n2751 = n1019 | n1021;
  assign n3469 = n1082 & n2751;
  assign n3470 = n1019 & n1082;
  assign n3471 = (n2737 & n3469) | (n2737 & n3470) | (n3469 & n3470);
  assign n3472 = n1082 | n2751;
  assign n3473 = n1019 | n1082;
  assign n3474 = (n2737 & n3472) | (n2737 & n3473) | (n3472 & n3473);
  assign n1085 = ~n3471 & n3474;
  assign n1086 = x21 & x36;
  assign n1087 = n1085 & n1086;
  assign n1088 = n1085 | n1086;
  assign n1089 = ~n1087 & n1088;
  assign n1090 = n2750 & n1089;
  assign n1091 = n2750 | n1089;
  assign n1092 = ~n1090 & n1091;
  assign n1093 = x20 & x37;
  assign n1094 = n1092 & n1093;
  assign n1095 = n1092 | n1093;
  assign n1096 = ~n1094 & n1095;
  assign n1097 = n1059 & n1096;
  assign n1098 = n1059 | n1096;
  assign n1099 = ~n1097 & n1098;
  assign n1100 = x19 & x38;
  assign n1101 = n1099 & n1100;
  assign n1102 = n1099 | n1100;
  assign n1103 = ~n1101 & n1102;
  assign n1104 = n2748 & n1103;
  assign n1105 = n2748 | n1103;
  assign n1106 = ~n1104 & n1105;
  assign n1107 = x18 & x39;
  assign n1108 = n1106 & n1107;
  assign n1109 = n1106 | n1107;
  assign n1110 = ~n1108 & n1109;
  assign n1111 = n2746 & n1110;
  assign n1112 = n2746 | n1110;
  assign n1113 = ~n1111 & n1112;
  assign n1114 = x17 & x40;
  assign n1115 = n1113 & n1114;
  assign n1116 = n1113 | n1114;
  assign n1117 = ~n1115 & n1116;
  assign n1118 = n1054 & n1117;
  assign n1119 = n1054 | n1117;
  assign n1120 = ~n1118 & n1119;
  assign n1121 = x16 & x41;
  assign n1122 = n1120 & n1121;
  assign n1123 = n1120 | n1121;
  assign n1124 = ~n1122 & n1123;
  assign n3901 = n1053 | n1114;
  assign n3902 = (n1052 & n1114) | (n1052 & n3901) | (n1114 & n3901);
  assign n3476 = (n1054 & n1113) | (n1054 & n3902) | (n1113 & n3902);
  assign n2771 = (n1115 & n1117) | (n1115 & n3476) | (n1117 & n3476);
  assign n2772 = n1108 | n2746;
  assign n2773 = (n1108 & n1110) | (n1108 & n2772) | (n1110 & n2772);
  assign n2774 = n1101 | n2748;
  assign n2775 = (n1101 & n1103) | (n1101 & n2774) | (n1103 & n2774);
  assign n2776 = n1094 | n1096;
  assign n2777 = (n1059 & n1094) | (n1059 & n2776) | (n1094 & n2776);
  assign n2752 = (n1019 & n2737) | (n1019 & n2751) | (n2737 & n2751);
  assign n3477 = n1066 | n1068;
  assign n3478 = (n1066 & n3462) | (n1066 & n3477) | (n3462 & n3477);
  assign n3479 = (n1066 & n2756) | (n1066 & n3477) | (n2756 & n3477);
  assign n3480 = (n2725 & n3478) | (n2725 & n3479) | (n3478 & n3479);
  assign n3481 = (n2724 & n3478) | (n2724 & n3479) | (n3478 & n3479);
  assign n3482 = (n2697 & n3480) | (n2697 & n3481) | (n3480 & n3481);
  assign n1133 = x26 & x32;
  assign n1134 = x25 & x33;
  assign n1135 = n1133 & n1134;
  assign n1136 = n1133 | n1134;
  assign n1137 = ~n1135 & n1136;
  assign n1138 = n3482 & n1137;
  assign n1139 = n3482 | n1137;
  assign n1140 = ~n1138 & n1139;
  assign n1141 = x24 & x34;
  assign n1142 = n1140 & n1141;
  assign n1143 = n1140 | n1141;
  assign n1144 = ~n1142 & n1143;
  assign n2785 = n1073 & n1144;
  assign n3483 = (n1144 & n2764) | (n1144 & n2785) | (n2764 & n2785);
  assign n3484 = (n1144 & n2765) | (n1144 & n2785) | (n2765 & n2785);
  assign n3485 = (n2740 & n3483) | (n2740 & n3484) | (n3483 & n3484);
  assign n2787 = n1073 | n1144;
  assign n3486 = n2764 | n2787;
  assign n3487 = n2765 | n2787;
  assign n3488 = (n2740 & n3486) | (n2740 & n3487) | (n3486 & n3487);
  assign n1147 = ~n3485 & n3488;
  assign n1148 = x23 & x35;
  assign n1149 = n1147 & n1148;
  assign n1150 = n1147 | n1148;
  assign n1151 = ~n1149 & n1150;
  assign n2780 = n1080 | n1082;
  assign n2789 = n1151 & n2780;
  assign n2790 = n1080 & n1151;
  assign n2791 = (n2752 & n2789) | (n2752 & n2790) | (n2789 & n2790);
  assign n2792 = n1151 | n2780;
  assign n2793 = n1080 | n1151;
  assign n2794 = (n2752 & n2792) | (n2752 & n2793) | (n2792 & n2793);
  assign n1154 = ~n2791 & n2794;
  assign n1155 = x22 & x36;
  assign n1156 = n1154 & n1155;
  assign n1157 = n1154 | n1155;
  assign n1158 = ~n1156 & n1157;
  assign n2778 = n1087 | n1089;
  assign n3489 = n1158 & n2778;
  assign n3490 = n1087 & n1158;
  assign n3491 = (n2750 & n3489) | (n2750 & n3490) | (n3489 & n3490);
  assign n3492 = n1158 | n2778;
  assign n3493 = n1087 | n1158;
  assign n3494 = (n2750 & n3492) | (n2750 & n3493) | (n3492 & n3493);
  assign n1161 = ~n3491 & n3494;
  assign n1162 = x21 & x37;
  assign n1163 = n1161 & n1162;
  assign n1164 = n1161 | n1162;
  assign n1165 = ~n1163 & n1164;
  assign n1166 = n2777 & n1165;
  assign n1167 = n2777 | n1165;
  assign n1168 = ~n1166 & n1167;
  assign n1169 = x20 & x38;
  assign n1170 = n1168 & n1169;
  assign n1171 = n1168 | n1169;
  assign n1172 = ~n1170 & n1171;
  assign n1173 = n2775 & n1172;
  assign n1174 = n2775 | n1172;
  assign n1175 = ~n1173 & n1174;
  assign n1176 = x19 & x39;
  assign n1177 = n1175 & n1176;
  assign n1178 = n1175 | n1176;
  assign n1179 = ~n1177 & n1178;
  assign n1180 = n2773 & n1179;
  assign n1181 = n2773 | n1179;
  assign n1182 = ~n1180 & n1181;
  assign n1183 = x18 & x40;
  assign n1184 = n1182 & n1183;
  assign n1185 = n1182 | n1183;
  assign n1186 = ~n1184 & n1185;
  assign n1187 = n2771 & n1186;
  assign n1188 = n2771 | n1186;
  assign n1189 = ~n1187 & n1188;
  assign n1190 = x17 & x41;
  assign n1191 = n1189 & n1190;
  assign n1192 = n1189 | n1190;
  assign n1193 = ~n1191 & n1192;
  assign n1194 = n1122 & n1193;
  assign n1195 = n1122 | n1193;
  assign n1196 = ~n1194 & n1195;
  assign n1197 = x16 & x42;
  assign n1198 = n1196 & n1197;
  assign n1199 = n1196 | n1197;
  assign n1200 = ~n1198 & n1199;
  assign n2795 = n1122 | n1191;
  assign n2796 = (n1191 & n1193) | (n1191 & n2795) | (n1193 & n2795);
  assign n1202 = n1184 | n1187;
  assign n1203 = n1177 | n1180;
  assign n2779 = (n1087 & n2750) | (n1087 & n2778) | (n2750 & n2778);
  assign n2802 = n1142 | n1144;
  assign n3495 = n1073 | n1142;
  assign n3496 = (n1142 & n1144) | (n1142 & n3495) | (n1144 & n3495);
  assign n3497 = (n2764 & n2802) | (n2764 & n3496) | (n2802 & n3496);
  assign n3498 = (n2765 & n2802) | (n2765 & n3496) | (n2802 & n3496);
  assign n3499 = (n2740 & n3497) | (n2740 & n3498) | (n3497 & n3498);
  assign n1210 = x27 & x32;
  assign n1211 = x26 & x33;
  assign n1212 = n1210 & n1211;
  assign n1213 = n1210 | n1211;
  assign n1214 = ~n1212 & n1213;
  assign n2804 = n1135 | n1137;
  assign n2806 = n1214 & n2804;
  assign n2807 = n1135 & n1214;
  assign n2808 = (n3482 & n2806) | (n3482 & n2807) | (n2806 & n2807);
  assign n2809 = n1214 | n2804;
  assign n2810 = n1135 | n1214;
  assign n2811 = (n3482 & n2809) | (n3482 & n2810) | (n2809 & n2810);
  assign n1217 = ~n2808 & n2811;
  assign n1218 = x25 & x34;
  assign n1219 = n1217 & n1218;
  assign n1220 = n1217 | n1218;
  assign n1221 = ~n1219 & n1220;
  assign n1222 = n3499 & n1221;
  assign n1223 = n3499 | n1221;
  assign n1224 = ~n1222 & n1223;
  assign n1225 = x24 & x35;
  assign n1226 = n1224 & n1225;
  assign n1227 = n1224 | n1225;
  assign n1228 = ~n1226 & n1227;
  assign n2812 = n1149 & n1228;
  assign n2813 = (n1228 & n2791) | (n1228 & n2812) | (n2791 & n2812);
  assign n2814 = n1149 | n1228;
  assign n2815 = n2791 | n2814;
  assign n1231 = ~n2813 & n2815;
  assign n1232 = x23 & x36;
  assign n1233 = n1231 & n1232;
  assign n1234 = n1231 | n1232;
  assign n1235 = ~n1233 & n1234;
  assign n2799 = n1156 | n1158;
  assign n2816 = n1235 & n2799;
  assign n2817 = n1156 & n1235;
  assign n2818 = (n2779 & n2816) | (n2779 & n2817) | (n2816 & n2817);
  assign n2819 = n1235 | n2799;
  assign n2820 = n1156 | n1235;
  assign n2821 = (n2779 & n2819) | (n2779 & n2820) | (n2819 & n2820);
  assign n1238 = ~n2818 & n2821;
  assign n1239 = x22 & x37;
  assign n1240 = n1238 & n1239;
  assign n1241 = n1238 | n1239;
  assign n1242 = ~n1240 & n1241;
  assign n2797 = n1163 | n1165;
  assign n3500 = n1242 & n2797;
  assign n3501 = n1163 & n1242;
  assign n3502 = (n2777 & n3500) | (n2777 & n3501) | (n3500 & n3501);
  assign n3503 = n1242 | n2797;
  assign n3504 = n1163 | n1242;
  assign n3505 = (n2777 & n3503) | (n2777 & n3504) | (n3503 & n3504);
  assign n1245 = ~n3502 & n3505;
  assign n1246 = x21 & x38;
  assign n1247 = n1245 & n1246;
  assign n1248 = n1245 | n1246;
  assign n1249 = ~n1247 & n1248;
  assign n3506 = n1170 & n1249;
  assign n3507 = (n1173 & n1249) | (n1173 & n3506) | (n1249 & n3506);
  assign n3508 = n1170 | n1249;
  assign n3509 = n1173 | n3508;
  assign n1252 = ~n3507 & n3509;
  assign n1253 = x20 & x39;
  assign n1254 = n1252 & n1253;
  assign n1255 = n1252 | n1253;
  assign n1256 = ~n1254 & n1255;
  assign n1257 = n1203 & n1256;
  assign n1258 = n1203 | n1256;
  assign n1259 = ~n1257 & n1258;
  assign n1260 = x19 & x40;
  assign n1261 = n1259 & n1260;
  assign n1262 = n1259 | n1260;
  assign n1263 = ~n1261 & n1262;
  assign n1264 = n1202 & n1263;
  assign n1265 = n1202 | n1263;
  assign n1266 = ~n1264 & n1265;
  assign n1267 = x18 & x41;
  assign n1268 = n1266 & n1267;
  assign n1269 = n1266 | n1267;
  assign n1270 = ~n1268 & n1269;
  assign n1271 = n2796 & n1270;
  assign n1272 = n2796 | n1270;
  assign n1273 = ~n1271 & n1272;
  assign n1274 = x17 & x42;
  assign n1275 = n1273 & n1274;
  assign n1276 = n1273 | n1274;
  assign n1277 = ~n1275 & n1276;
  assign n1278 = n1198 & n1277;
  assign n1279 = n1198 | n1277;
  assign n1280 = ~n1278 & n1279;
  assign n1281 = x16 & x43;
  assign n1282 = n1280 & n1281;
  assign n1283 = n1280 | n1281;
  assign n1284 = ~n1282 & n1283;
  assign n3903 = n1197 | n1274;
  assign n3904 = (n1196 & n1274) | (n1196 & n3903) | (n1274 & n3903);
  assign n3511 = (n1198 & n1273) | (n1198 & n3904) | (n1273 & n3904);
  assign n2823 = (n1275 & n1277) | (n1275 & n3511) | (n1277 & n3511);
  assign n2824 = n1268 | n2796;
  assign n2825 = (n1268 & n1270) | (n1268 & n2824) | (n1270 & n2824);
  assign n1287 = n1261 | n1264;
  assign n3512 = n1254 | n1256;
  assign n3513 = (n1203 & n1254) | (n1203 & n3512) | (n1254 & n3512);
  assign n1204 = n1170 | n1173;
  assign n2798 = (n1163 & n2777) | (n1163 & n2797) | (n2777 & n2797);
  assign n1295 = x28 & x32;
  assign n1296 = x27 & x33;
  assign n1297 = n1295 & n1296;
  assign n1298 = n1295 | n1296;
  assign n1299 = ~n1297 & n1298;
  assign n3514 = n1212 | n1214;
  assign n3515 = (n1212 & n2804) | (n1212 & n3514) | (n2804 & n3514);
  assign n2835 = n1299 & n3515;
  assign n3516 = n1135 | n1212;
  assign n3517 = (n1212 & n1214) | (n1212 & n3516) | (n1214 & n3516);
  assign n2836 = n1299 & n3517;
  assign n2837 = (n3482 & n2835) | (n3482 & n2836) | (n2835 & n2836);
  assign n2838 = n1299 | n3515;
  assign n2839 = n1299 | n3517;
  assign n2840 = (n3482 & n2838) | (n3482 & n2839) | (n2838 & n2839);
  assign n1302 = ~n2837 & n2840;
  assign n1303 = x26 & x34;
  assign n1304 = n1302 & n1303;
  assign n1305 = n1302 | n1303;
  assign n1306 = ~n1304 & n1305;
  assign n2830 = n1219 | n1221;
  assign n2841 = n1306 & n2830;
  assign n2842 = n1219 & n1306;
  assign n2843 = (n3499 & n2841) | (n3499 & n2842) | (n2841 & n2842);
  assign n2844 = n1306 | n2830;
  assign n2845 = n1219 | n1306;
  assign n2846 = (n3499 & n2844) | (n3499 & n2845) | (n2844 & n2845);
  assign n1309 = ~n2843 & n2846;
  assign n1310 = x25 & x35;
  assign n1311 = n1309 & n1310;
  assign n1312 = n1309 | n1310;
  assign n1313 = ~n1311 & n1312;
  assign n2847 = n1226 & n1313;
  assign n3518 = (n1313 & n2812) | (n1313 & n2847) | (n2812 & n2847);
  assign n3519 = (n1228 & n1313) | (n1228 & n2847) | (n1313 & n2847);
  assign n3520 = (n2791 & n3518) | (n2791 & n3519) | (n3518 & n3519);
  assign n2849 = n1226 | n1313;
  assign n3521 = n2812 | n2849;
  assign n3522 = n1228 | n2849;
  assign n3523 = (n2791 & n3521) | (n2791 & n3522) | (n3521 & n3522);
  assign n1316 = ~n3520 & n3523;
  assign n1317 = x24 & x36;
  assign n1318 = n1316 & n1317;
  assign n1319 = n1316 | n1317;
  assign n1320 = ~n1318 & n1319;
  assign n2851 = n1233 & n1320;
  assign n2852 = (n1320 & n2818) | (n1320 & n2851) | (n2818 & n2851);
  assign n2853 = n1233 | n1320;
  assign n2854 = n2818 | n2853;
  assign n1323 = ~n2852 & n2854;
  assign n1324 = x23 & x37;
  assign n1325 = n1323 & n1324;
  assign n1326 = n1323 | n1324;
  assign n1327 = ~n1325 & n1326;
  assign n2828 = n1240 | n1242;
  assign n2855 = n1327 & n2828;
  assign n2856 = n1240 & n1327;
  assign n2857 = (n2798 & n2855) | (n2798 & n2856) | (n2855 & n2856);
  assign n2858 = n1327 | n2828;
  assign n2859 = n1240 | n1327;
  assign n2860 = (n2798 & n2858) | (n2798 & n2859) | (n2858 & n2859);
  assign n1330 = ~n2857 & n2860;
  assign n1331 = x22 & x38;
  assign n1332 = n1330 & n1331;
  assign n1333 = n1330 | n1331;
  assign n1334 = ~n1332 & n1333;
  assign n2826 = n1247 | n1249;
  assign n3524 = n1334 & n2826;
  assign n3525 = n1247 & n1334;
  assign n3526 = (n1204 & n3524) | (n1204 & n3525) | (n3524 & n3525);
  assign n3527 = n1334 | n2826;
  assign n3528 = n1247 | n1334;
  assign n3529 = (n1204 & n3527) | (n1204 & n3528) | (n3527 & n3528);
  assign n1337 = ~n3526 & n3529;
  assign n1338 = x21 & x39;
  assign n1339 = n1337 & n1338;
  assign n1340 = n1337 | n1338;
  assign n1341 = ~n1339 & n1340;
  assign n1342 = n3513 & n1341;
  assign n1343 = n3513 | n1341;
  assign n1344 = ~n1342 & n1343;
  assign n1345 = x20 & x40;
  assign n1346 = n1344 & n1345;
  assign n1347 = n1344 | n1345;
  assign n1348 = ~n1346 & n1347;
  assign n1349 = n1287 & n1348;
  assign n1350 = n1287 | n1348;
  assign n1351 = ~n1349 & n1350;
  assign n1352 = x19 & x41;
  assign n1353 = n1351 & n1352;
  assign n1354 = n1351 | n1352;
  assign n1355 = ~n1353 & n1354;
  assign n1356 = n2825 & n1355;
  assign n1357 = n2825 | n1355;
  assign n1358 = ~n1356 & n1357;
  assign n1359 = x18 & x42;
  assign n1360 = n1358 & n1359;
  assign n1361 = n1358 | n1359;
  assign n1362 = ~n1360 & n1361;
  assign n1363 = n2823 & n1362;
  assign n1364 = n2823 | n1362;
  assign n1365 = ~n1363 & n1364;
  assign n1366 = x17 & x43;
  assign n1367 = n1365 & n1366;
  assign n1368 = n1365 | n1366;
  assign n1369 = ~n1367 & n1368;
  assign n1370 = n1282 & n1369;
  assign n1371 = n1282 | n1369;
  assign n1372 = ~n1370 & n1371;
  assign n1373 = x16 & x44;
  assign n1374 = n1372 & n1373;
  assign n1375 = n1372 | n1373;
  assign n1376 = ~n1374 & n1375;
  assign n3905 = n1281 | n1366;
  assign n3906 = (n1280 & n1366) | (n1280 & n3905) | (n1366 & n3905);
  assign n3531 = (n1282 & n1365) | (n1282 & n3906) | (n1365 & n3906);
  assign n2862 = (n1367 & n1369) | (n1367 & n3531) | (n1369 & n3531);
  assign n2863 = n1360 | n2823;
  assign n2864 = (n1360 & n1362) | (n1360 & n2863) | (n1362 & n2863);
  assign n2865 = n1353 | n2825;
  assign n2866 = (n1353 & n1355) | (n1353 & n2865) | (n1355 & n2865);
  assign n3532 = n1346 | n1348;
  assign n3533 = (n1287 & n1346) | (n1287 & n3532) | (n1346 & n3532);
  assign n2867 = n1339 | n1341;
  assign n2868 = (n3513 & n1339) | (n3513 & n2867) | (n1339 & n2867);
  assign n2827 = (n1204 & n1247) | (n1204 & n2826) | (n1247 & n2826);
  assign n2872 = n1311 | n1313;
  assign n3534 = n1226 | n1311;
  assign n3535 = (n1311 & n1313) | (n1311 & n3534) | (n1313 & n3534);
  assign n3536 = (n2812 & n2872) | (n2812 & n3535) | (n2872 & n3535);
  assign n3537 = (n1228 & n2872) | (n1228 & n3535) | (n2872 & n3535);
  assign n3538 = (n2791 & n3536) | (n2791 & n3537) | (n3536 & n3537);
  assign n1388 = x29 & x32;
  assign n1389 = x28 & x33;
  assign n1390 = n1388 & n1389;
  assign n1391 = n1388 | n1389;
  assign n1392 = ~n1390 & n1391;
  assign n3543 = n1297 | n1299;
  assign n3907 = n1392 & n3543;
  assign n3908 = n1297 & n1392;
  assign n3909 = (n3515 & n3907) | (n3515 & n3908) | (n3907 & n3908);
  assign n3545 = (n1297 & n3517) | (n1297 & n3543) | (n3517 & n3543);
  assign n3547 = n1392 & n3545;
  assign n3548 = (n3482 & n3909) | (n3482 & n3547) | (n3909 & n3547);
  assign n3910 = n1392 | n3543;
  assign n3911 = n1297 | n1392;
  assign n3912 = (n3515 & n3910) | (n3515 & n3911) | (n3910 & n3911);
  assign n3550 = n1392 | n3545;
  assign n3551 = (n3482 & n3912) | (n3482 & n3550) | (n3912 & n3550);
  assign n1395 = ~n3548 & n3551;
  assign n1396 = x27 & x34;
  assign n1397 = n1395 & n1396;
  assign n1398 = n1395 | n1396;
  assign n1399 = ~n1397 & n1398;
  assign n3539 = n1304 | n1306;
  assign n3540 = (n1304 & n2830) | (n1304 & n3539) | (n2830 & n3539);
  assign n3552 = n1399 & n3540;
  assign n3541 = n1219 | n1304;
  assign n3542 = (n1304 & n1306) | (n1304 & n3541) | (n1306 & n3541);
  assign n3553 = n1399 & n3542;
  assign n3554 = (n3499 & n3552) | (n3499 & n3553) | (n3552 & n3553);
  assign n3555 = n1399 | n3540;
  assign n3556 = n1399 | n3542;
  assign n3557 = (n3499 & n3555) | (n3499 & n3556) | (n3555 & n3556);
  assign n1402 = ~n3554 & n3557;
  assign n1403 = x26 & x35;
  assign n1404 = n1402 & n1403;
  assign n1405 = n1402 | n1403;
  assign n1406 = ~n1404 & n1405;
  assign n1407 = n3538 & n1406;
  assign n1408 = n3538 | n1406;
  assign n1409 = ~n1407 & n1408;
  assign n1410 = x25 & x36;
  assign n1411 = n1409 & n1410;
  assign n1412 = n1409 | n1410;
  assign n1413 = ~n1411 & n1412;
  assign n2880 = n1318 & n1413;
  assign n2881 = (n1413 & n2852) | (n1413 & n2880) | (n2852 & n2880);
  assign n2882 = n1318 | n1413;
  assign n2883 = n2852 | n2882;
  assign n1416 = ~n2881 & n2883;
  assign n1417 = x24 & x37;
  assign n1418 = n1416 & n1417;
  assign n1419 = n1416 | n1417;
  assign n1420 = ~n1418 & n1419;
  assign n2884 = n1325 & n1420;
  assign n2885 = (n1420 & n2857) | (n1420 & n2884) | (n2857 & n2884);
  assign n2886 = n1325 | n1420;
  assign n2887 = n2857 | n2886;
  assign n1423 = ~n2885 & n2887;
  assign n1424 = x23 & x38;
  assign n1425 = n1423 & n1424;
  assign n1426 = n1423 | n1424;
  assign n1427 = ~n1425 & n1426;
  assign n2869 = n1332 | n1334;
  assign n2888 = n1427 & n2869;
  assign n2889 = n1332 & n1427;
  assign n2890 = (n2827 & n2888) | (n2827 & n2889) | (n2888 & n2889);
  assign n2891 = n1427 | n2869;
  assign n2892 = n1332 | n1427;
  assign n2893 = (n2827 & n2891) | (n2827 & n2892) | (n2891 & n2892);
  assign n1430 = ~n2890 & n2893;
  assign n1431 = x22 & x39;
  assign n1432 = n1430 & n1431;
  assign n1433 = n1430 | n1431;
  assign n1434 = ~n1432 & n1433;
  assign n1435 = n2868 & n1434;
  assign n1436 = n2868 | n1434;
  assign n1437 = ~n1435 & n1436;
  assign n1438 = x21 & x40;
  assign n1439 = n1437 & n1438;
  assign n1440 = n1437 | n1438;
  assign n1441 = ~n1439 & n1440;
  assign n1442 = n3533 & n1441;
  assign n1443 = n3533 | n1441;
  assign n1444 = ~n1442 & n1443;
  assign n1445 = x20 & x41;
  assign n1446 = n1444 & n1445;
  assign n1447 = n1444 | n1445;
  assign n1448 = ~n1446 & n1447;
  assign n1449 = n2866 & n1448;
  assign n1450 = n2866 | n1448;
  assign n1451 = ~n1449 & n1450;
  assign n1452 = x19 & x42;
  assign n1453 = n1451 & n1452;
  assign n1454 = n1451 | n1452;
  assign n1455 = ~n1453 & n1454;
  assign n1456 = n2864 & n1455;
  assign n1457 = n2864 | n1455;
  assign n1458 = ~n1456 & n1457;
  assign n1459 = x18 & x43;
  assign n1460 = n1458 & n1459;
  assign n1461 = n1458 | n1459;
  assign n1462 = ~n1460 & n1461;
  assign n1463 = n2862 & n1462;
  assign n1464 = n2862 | n1462;
  assign n1465 = ~n1463 & n1464;
  assign n1466 = x17 & x44;
  assign n1467 = n1465 & n1466;
  assign n1468 = n1465 | n1466;
  assign n1469 = ~n1467 & n1468;
  assign n1470 = n1374 & n1469;
  assign n1471 = n1374 | n1469;
  assign n1472 = ~n1470 & n1471;
  assign n1473 = x16 & x45;
  assign n1474 = n1472 & n1473;
  assign n1475 = n1472 | n1473;
  assign n1476 = ~n1474 & n1475;
  assign n2894 = n1374 | n1467;
  assign n2895 = (n1467 & n1469) | (n1467 & n2894) | (n1469 & n2894);
  assign n2896 = n1460 | n2862;
  assign n2897 = (n1460 & n1462) | (n1460 & n2896) | (n1462 & n2896);
  assign n2898 = n1453 | n2864;
  assign n2899 = (n1453 & n1455) | (n1453 & n2898) | (n1455 & n2898);
  assign n2900 = n1446 | n2866;
  assign n2901 = (n1446 & n1448) | (n1446 & n2900) | (n1448 & n2900);
  assign n2902 = n1439 | n1441;
  assign n2903 = (n3533 & n1439) | (n3533 & n2902) | (n1439 & n2902);
  assign n1489 = x30 & x32;
  assign n1490 = x29 & x33;
  assign n1491 = n1489 & n1490;
  assign n1492 = n1489 | n1490;
  assign n1493 = ~n1491 & n1492;
  assign n2910 = n1390 | n1392;
  assign n2912 = n1493 & n2910;
  assign n2913 = n1390 & n1493;
  assign n3544 = (n1297 & n3515) | (n1297 & n3543) | (n3515 & n3543);
  assign n3558 = (n2912 & n2913) | (n2912 & n3544) | (n2913 & n3544);
  assign n3559 = (n2912 & n2913) | (n2912 & n3545) | (n2913 & n3545);
  assign n3560 = (n3482 & n3558) | (n3482 & n3559) | (n3558 & n3559);
  assign n2915 = n1493 | n2910;
  assign n2916 = n1390 | n1493;
  assign n3561 = (n2915 & n2916) | (n2915 & n3544) | (n2916 & n3544);
  assign n3562 = (n2915 & n2916) | (n2915 & n3545) | (n2916 & n3545);
  assign n3563 = (n3482 & n3561) | (n3482 & n3562) | (n3561 & n3562);
  assign n1496 = ~n3560 & n3563;
  assign n1497 = x28 & x34;
  assign n1498 = n1496 & n1497;
  assign n1499 = n1496 | n1497;
  assign n1500 = ~n1498 & n1499;
  assign n2908 = n1397 | n1399;
  assign n2918 = n1500 & n2908;
  assign n2919 = n1397 & n1500;
  assign n3564 = (n2918 & n2919) | (n2918 & n3540) | (n2919 & n3540);
  assign n3565 = (n2918 & n2919) | (n2918 & n3542) | (n2919 & n3542);
  assign n3566 = (n3499 & n3564) | (n3499 & n3565) | (n3564 & n3565);
  assign n2921 = n1500 | n2908;
  assign n2922 = n1397 | n1500;
  assign n3567 = (n2921 & n2922) | (n2921 & n3540) | (n2922 & n3540);
  assign n3568 = (n2921 & n2922) | (n2921 & n3542) | (n2922 & n3542);
  assign n3569 = (n3499 & n3567) | (n3499 & n3568) | (n3567 & n3568);
  assign n1503 = ~n3566 & n3569;
  assign n1504 = x27 & x35;
  assign n1505 = n1503 & n1504;
  assign n1506 = n1503 | n1504;
  assign n1507 = ~n1505 & n1506;
  assign n2906 = n1404 | n1406;
  assign n2924 = n1507 & n2906;
  assign n2925 = n1404 & n1507;
  assign n2926 = (n3538 & n2924) | (n3538 & n2925) | (n2924 & n2925);
  assign n2927 = n1507 | n2906;
  assign n2928 = n1404 | n1507;
  assign n2929 = (n3538 & n2927) | (n3538 & n2928) | (n2927 & n2928);
  assign n1510 = ~n2926 & n2929;
  assign n1511 = x26 & x36;
  assign n1512 = n1510 & n1511;
  assign n1513 = n1510 | n1511;
  assign n1514 = ~n1512 & n1513;
  assign n2930 = n1411 & n1514;
  assign n3570 = (n1514 & n2880) | (n1514 & n2930) | (n2880 & n2930);
  assign n3571 = (n1413 & n1514) | (n1413 & n2930) | (n1514 & n2930);
  assign n3572 = (n2852 & n3570) | (n2852 & n3571) | (n3570 & n3571);
  assign n2932 = n1411 | n1514;
  assign n3573 = n2880 | n2932;
  assign n3574 = n1413 | n2932;
  assign n3575 = (n2852 & n3573) | (n2852 & n3574) | (n3573 & n3574);
  assign n1517 = ~n3572 & n3575;
  assign n1518 = x25 & x37;
  assign n1519 = n1517 & n1518;
  assign n1520 = n1517 | n1518;
  assign n1521 = ~n1519 & n1520;
  assign n2934 = n1418 & n1521;
  assign n2935 = (n1521 & n2885) | (n1521 & n2934) | (n2885 & n2934);
  assign n2936 = n1418 | n1521;
  assign n2937 = n2885 | n2936;
  assign n1524 = ~n2935 & n2937;
  assign n1525 = x24 & x38;
  assign n1526 = n1524 & n1525;
  assign n1527 = n1524 | n1525;
  assign n1528 = ~n1526 & n1527;
  assign n2938 = n1425 & n1528;
  assign n2939 = (n1528 & n2890) | (n1528 & n2938) | (n2890 & n2938);
  assign n2940 = n1425 | n1528;
  assign n2941 = n2890 | n2940;
  assign n1531 = ~n2939 & n2941;
  assign n1532 = x23 & x39;
  assign n1533 = n1531 & n1532;
  assign n1534 = n1531 | n1532;
  assign n1535 = ~n1533 & n1534;
  assign n2904 = n1432 | n1434;
  assign n2942 = n1535 & n2904;
  assign n2943 = n1432 & n1535;
  assign n2944 = (n2868 & n2942) | (n2868 & n2943) | (n2942 & n2943);
  assign n2945 = n1535 | n2904;
  assign n2946 = n1432 | n1535;
  assign n2947 = (n2868 & n2945) | (n2868 & n2946) | (n2945 & n2946);
  assign n1538 = ~n2944 & n2947;
  assign n1539 = x22 & x40;
  assign n1540 = n1538 & n1539;
  assign n1541 = n1538 | n1539;
  assign n1542 = ~n1540 & n1541;
  assign n1543 = n2903 & n1542;
  assign n1544 = n2903 | n1542;
  assign n1545 = ~n1543 & n1544;
  assign n1546 = x21 & x41;
  assign n1547 = n1545 & n1546;
  assign n1548 = n1545 | n1546;
  assign n1549 = ~n1547 & n1548;
  assign n1550 = n2901 & n1549;
  assign n1551 = n2901 | n1549;
  assign n1552 = ~n1550 & n1551;
  assign n1553 = x20 & x42;
  assign n1554 = n1552 & n1553;
  assign n1555 = n1552 | n1553;
  assign n1556 = ~n1554 & n1555;
  assign n1557 = n2899 & n1556;
  assign n1558 = n2899 | n1556;
  assign n1559 = ~n1557 & n1558;
  assign n1560 = x19 & x43;
  assign n1561 = n1559 & n1560;
  assign n1562 = n1559 | n1560;
  assign n1563 = ~n1561 & n1562;
  assign n1564 = n2897 & n1563;
  assign n1565 = n2897 | n1563;
  assign n1566 = ~n1564 & n1565;
  assign n1567 = x18 & x44;
  assign n1568 = n1566 & n1567;
  assign n1569 = n1566 | n1567;
  assign n1570 = ~n1568 & n1569;
  assign n1571 = n2895 & n1570;
  assign n1572 = n2895 | n1570;
  assign n1573 = ~n1571 & n1572;
  assign n1574 = x17 & x45;
  assign n1575 = n1573 & n1574;
  assign n1576 = n1573 | n1574;
  assign n1577 = ~n1575 & n1576;
  assign n1578 = n1474 & n1577;
  assign n1579 = n1474 | n1577;
  assign n1580 = ~n1578 & n1579;
  assign n1581 = x16 & x46;
  assign n1582 = n1580 & n1581;
  assign n1583 = n1580 | n1581;
  assign n1584 = ~n1582 & n1583;
  assign n3913 = n1473 | n1574;
  assign n3914 = (n1472 & n1574) | (n1472 & n3913) | (n1574 & n3913);
  assign n3577 = (n1474 & n1573) | (n1474 & n3914) | (n1573 & n3914);
  assign n2949 = (n1575 & n1577) | (n1575 & n3577) | (n1577 & n3577);
  assign n3578 = n1568 | n2895;
  assign n3579 = (n1568 & n1570) | (n1568 & n3578) | (n1570 & n3578);
  assign n1587 = n1561 | n1564;
  assign n1588 = n1554 | n1557;
  assign n2953 = n1512 | n1514;
  assign n3580 = n1411 | n1512;
  assign n3581 = (n1512 & n1514) | (n1512 & n3580) | (n1514 & n3580);
  assign n3582 = (n2880 & n2953) | (n2880 & n3581) | (n2953 & n3581);
  assign n3583 = (n1413 & n2953) | (n1413 & n3581) | (n2953 & n3581);
  assign n3584 = (n2852 & n3582) | (n2852 & n3583) | (n3582 & n3583);
  assign n3585 = n1498 | n1500;
  assign n3586 = (n1498 & n2908) | (n1498 & n3585) | (n2908 & n3585);
  assign n3587 = n1397 | n1498;
  assign n3588 = (n1498 & n1500) | (n1498 & n3587) | (n1500 & n3587);
  assign n3589 = (n3540 & n3586) | (n3540 & n3588) | (n3586 & n3588);
  assign n3590 = (n3542 & n3586) | (n3542 & n3588) | (n3586 & n3588);
  assign n3591 = (n3499 & n3589) | (n3499 & n3590) | (n3589 & n3590);
  assign n1598 = x31 & x32;
  assign n1599 = x30 & x33;
  assign n1600 = n1598 & n1599;
  assign n1601 = n1598 | n1599;
  assign n1602 = ~n1600 & n1601;
  assign n3592 = n1491 | n1493;
  assign n3593 = (n1491 & n2910) | (n1491 & n3592) | (n2910 & n3592);
  assign n2961 = n1602 & n3593;
  assign n3594 = n1390 | n1491;
  assign n3595 = (n1491 & n1493) | (n1491 & n3594) | (n1493 & n3594);
  assign n2962 = n1602 & n3595;
  assign n3596 = (n2961 & n2962) | (n2961 & n3544) | (n2962 & n3544);
  assign n3597 = (n2961 & n2962) | (n2961 & n3545) | (n2962 & n3545);
  assign n3598 = (n3482 & n3596) | (n3482 & n3597) | (n3596 & n3597);
  assign n2964 = n1602 | n3593;
  assign n2965 = n1602 | n3595;
  assign n3599 = (n2964 & n2965) | (n2964 & n3544) | (n2965 & n3544);
  assign n3600 = (n2964 & n2965) | (n2964 & n3545) | (n2965 & n3545);
  assign n3601 = (n3482 & n3599) | (n3482 & n3600) | (n3599 & n3600);
  assign n1605 = ~n3598 & n3601;
  assign n1606 = x29 & x34;
  assign n1607 = n1605 & n1606;
  assign n1608 = n1605 | n1606;
  assign n1609 = ~n1607 & n1608;
  assign n1610 = n3591 & n1609;
  assign n1611 = n3591 | n1609;
  assign n1612 = ~n1610 & n1611;
  assign n1613 = x28 & x35;
  assign n1614 = n1612 & n1613;
  assign n1615 = n1612 | n1613;
  assign n1616 = ~n1614 & n1615;
  assign n2967 = n1505 & n1616;
  assign n3602 = (n1616 & n2924) | (n1616 & n2967) | (n2924 & n2967);
  assign n3603 = (n1616 & n2925) | (n1616 & n2967) | (n2925 & n2967);
  assign n3604 = (n3538 & n3602) | (n3538 & n3603) | (n3602 & n3603);
  assign n2969 = n1505 | n1616;
  assign n3605 = n2924 | n2969;
  assign n3606 = n2925 | n2969;
  assign n3607 = (n3538 & n3605) | (n3538 & n3606) | (n3605 & n3606);
  assign n1619 = ~n3604 & n3607;
  assign n1620 = x27 & x36;
  assign n1621 = n1619 & n1620;
  assign n1622 = n1619 | n1620;
  assign n1623 = ~n1621 & n1622;
  assign n1624 = n3584 & n1623;
  assign n1625 = n3584 | n1623;
  assign n1626 = ~n1624 & n1625;
  assign n1627 = x26 & x37;
  assign n1628 = n1626 & n1627;
  assign n1629 = n1626 | n1627;
  assign n1630 = ~n1628 & n1629;
  assign n2971 = n1519 & n1630;
  assign n2972 = (n1630 & n2935) | (n1630 & n2971) | (n2935 & n2971);
  assign n2973 = n1519 | n1630;
  assign n2974 = n2935 | n2973;
  assign n1633 = ~n2972 & n2974;
  assign n1634 = x25 & x38;
  assign n1635 = n1633 & n1634;
  assign n1636 = n1633 | n1634;
  assign n1637 = ~n1635 & n1636;
  assign n2975 = n1526 & n1637;
  assign n2976 = (n1637 & n2939) | (n1637 & n2975) | (n2939 & n2975);
  assign n2977 = n1526 | n1637;
  assign n2978 = n2939 | n2977;
  assign n1640 = ~n2976 & n2978;
  assign n1641 = x24 & x39;
  assign n1642 = n1640 & n1641;
  assign n1643 = n1640 | n1641;
  assign n1644 = ~n1642 & n1643;
  assign n2979 = n1533 & n1644;
  assign n2980 = (n1644 & n2944) | (n1644 & n2979) | (n2944 & n2979);
  assign n2981 = n1533 | n1644;
  assign n2982 = n2944 | n2981;
  assign n1647 = ~n2980 & n2982;
  assign n1648 = x23 & x40;
  assign n1649 = n1647 & n1648;
  assign n1650 = n1647 | n1648;
  assign n1651 = ~n1649 & n1650;
  assign n2950 = n1540 | n1542;
  assign n2983 = n1651 & n2950;
  assign n2984 = n1540 & n1651;
  assign n2985 = (n2903 & n2983) | (n2903 & n2984) | (n2983 & n2984);
  assign n2986 = n1651 | n2950;
  assign n2987 = n1540 | n1651;
  assign n2988 = (n2903 & n2986) | (n2903 & n2987) | (n2986 & n2987);
  assign n1654 = ~n2985 & n2988;
  assign n1655 = x22 & x41;
  assign n1656 = n1654 & n1655;
  assign n1657 = n1654 | n1655;
  assign n1658 = ~n1656 & n1657;
  assign n2989 = n1547 & n1658;
  assign n2990 = (n1550 & n1658) | (n1550 & n2989) | (n1658 & n2989);
  assign n2991 = n1547 | n1658;
  assign n2992 = n1550 | n2991;
  assign n1661 = ~n2990 & n2992;
  assign n1662 = x21 & x42;
  assign n1663 = n1661 & n1662;
  assign n1664 = n1661 | n1662;
  assign n1665 = ~n1663 & n1664;
  assign n1666 = n1588 & n1665;
  assign n1667 = n1588 | n1665;
  assign n1668 = ~n1666 & n1667;
  assign n1669 = x20 & x43;
  assign n1670 = n1668 & n1669;
  assign n1671 = n1668 | n1669;
  assign n1672 = ~n1670 & n1671;
  assign n1673 = n1587 & n1672;
  assign n1674 = n1587 | n1672;
  assign n1675 = ~n1673 & n1674;
  assign n1676 = x19 & x44;
  assign n1677 = n1675 & n1676;
  assign n1678 = n1675 | n1676;
  assign n1679 = ~n1677 & n1678;
  assign n1680 = n3579 & n1679;
  assign n1681 = n3579 | n1679;
  assign n1682 = ~n1680 & n1681;
  assign n1683 = x18 & x45;
  assign n1684 = n1682 & n1683;
  assign n1685 = n1682 | n1683;
  assign n1686 = ~n1684 & n1685;
  assign n1687 = n2949 & n1686;
  assign n1688 = n2949 | n1686;
  assign n1689 = ~n1687 & n1688;
  assign n1690 = x17 & x46;
  assign n1691 = n1689 & n1690;
  assign n1692 = n1689 | n1690;
  assign n1693 = ~n1691 & n1692;
  assign n1694 = n1582 & n1693;
  assign n1695 = n1582 | n1693;
  assign n1696 = ~n1694 & n1695;
  assign n1697 = x16 & x47;
  assign n1698 = n1696 & n1697;
  assign n1699 = n1696 | n1697;
  assign n1700 = ~n1698 & n1699;
  assign n3915 = n1581 | n1690;
  assign n3916 = (n1580 & n1690) | (n1580 & n3915) | (n1690 & n3915);
  assign n3609 = (n1582 & n1689) | (n1582 & n3916) | (n1689 & n3916);
  assign n2994 = (n1691 & n1693) | (n1691 & n3609) | (n1693 & n3609);
  assign n2995 = n1684 | n2949;
  assign n2996 = (n1684 & n1686) | (n1684 & n2995) | (n1686 & n2995);
  assign n3610 = n1677 | n3579;
  assign n3611 = (n1677 & n1679) | (n1677 & n3610) | (n1679 & n3610);
  assign n1704 = n1670 | n1673;
  assign n2997 = n1663 | n1665;
  assign n2998 = (n1588 & n1663) | (n1588 & n2997) | (n1663 & n2997);
  assign n3002 = n1614 | n1616;
  assign n3612 = n1505 | n1614;
  assign n3613 = (n1614 & n1616) | (n1614 & n3612) | (n1616 & n3612);
  assign n3614 = (n2924 & n3002) | (n2924 & n3613) | (n3002 & n3613);
  assign n3615 = (n2925 & n3002) | (n2925 & n3613) | (n3002 & n3613);
  assign n3616 = (n3538 & n3614) | (n3538 & n3615) | (n3614 & n3615);
  assign n1715 = x31 & x33;
  assign n3617 = n1600 | n1602;
  assign n3622 = (n1600 & n3595) | (n1600 & n3617) | (n3595 & n3617);
  assign n3010 = n1715 & n3622;
  assign n3620 = n1600 & n1715;
  assign n3917 = (n1602 & n1715) | (n1602 & n3620) | (n1715 & n3620);
  assign n3621 = (n3593 & n3917) | (n3593 & n3620) | (n3917 & n3620);
  assign n3623 = (n3010 & n3544) | (n3010 & n3621) | (n3544 & n3621);
  assign n3624 = (n3010 & n3545) | (n3010 & n3621) | (n3545 & n3621);
  assign n3625 = (n3482 & n3623) | (n3482 & n3624) | (n3623 & n3624);
  assign n3013 = n1715 | n3622;
  assign n3627 = n1600 | n1715;
  assign n3918 = n1602 | n3627;
  assign n3628 = (n3593 & n3918) | (n3593 & n3627) | (n3918 & n3627);
  assign n3629 = (n3013 & n3544) | (n3013 & n3628) | (n3544 & n3628);
  assign n3630 = (n3013 & n3545) | (n3013 & n3628) | (n3545 & n3628);
  assign n3631 = (n3482 & n3629) | (n3482 & n3630) | (n3629 & n3630);
  assign n1718 = ~n3625 & n3631;
  assign n1719 = x30 & x34;
  assign n1720 = n1718 & n1719;
  assign n1721 = n1718 | n1719;
  assign n1722 = ~n1720 & n1721;
  assign n3004 = n1607 | n1609;
  assign n3015 = n1722 & n3004;
  assign n3016 = n1607 & n1722;
  assign n3017 = (n3591 & n3015) | (n3591 & n3016) | (n3015 & n3016);
  assign n3018 = n1722 | n3004;
  assign n3019 = n1607 | n1722;
  assign n3020 = (n3591 & n3018) | (n3591 & n3019) | (n3018 & n3019);
  assign n1725 = ~n3017 & n3020;
  assign n1726 = x29 & x35;
  assign n1727 = n1725 & n1726;
  assign n1728 = n1725 | n1726;
  assign n1729 = ~n1727 & n1728;
  assign n1730 = n3616 & n1729;
  assign n1731 = n3616 | n1729;
  assign n1732 = ~n1730 & n1731;
  assign n1733 = x28 & x36;
  assign n1734 = n1732 & n1733;
  assign n1735 = n1732 | n1733;
  assign n1736 = ~n1734 & n1735;
  assign n2999 = n1621 | n1623;
  assign n3021 = n1736 & n2999;
  assign n3022 = n1621 & n1736;
  assign n3023 = (n3584 & n3021) | (n3584 & n3022) | (n3021 & n3022);
  assign n3024 = n1736 | n2999;
  assign n3025 = n1621 | n1736;
  assign n3026 = (n3584 & n3024) | (n3584 & n3025) | (n3024 & n3025);
  assign n1739 = ~n3023 & n3026;
  assign n1740 = x27 & x37;
  assign n1741 = n1739 & n1740;
  assign n1742 = n1739 | n1740;
  assign n1743 = ~n1741 & n1742;
  assign n3027 = n1628 & n1743;
  assign n3632 = (n1743 & n2971) | (n1743 & n3027) | (n2971 & n3027);
  assign n3633 = (n1630 & n1743) | (n1630 & n3027) | (n1743 & n3027);
  assign n3634 = (n2935 & n3632) | (n2935 & n3633) | (n3632 & n3633);
  assign n3029 = n1628 | n1743;
  assign n3635 = n2971 | n3029;
  assign n3636 = n1630 | n3029;
  assign n3637 = (n2935 & n3635) | (n2935 & n3636) | (n3635 & n3636);
  assign n1746 = ~n3634 & n3637;
  assign n1747 = x26 & x38;
  assign n1748 = n1746 & n1747;
  assign n1749 = n1746 | n1747;
  assign n1750 = ~n1748 & n1749;
  assign n3031 = n1635 & n1750;
  assign n3032 = (n1750 & n2976) | (n1750 & n3031) | (n2976 & n3031);
  assign n3033 = n1635 | n1750;
  assign n3034 = n2976 | n3033;
  assign n1753 = ~n3032 & n3034;
  assign n1754 = x25 & x39;
  assign n1755 = n1753 & n1754;
  assign n1756 = n1753 | n1754;
  assign n1757 = ~n1755 & n1756;
  assign n3035 = n1642 & n1757;
  assign n3036 = (n1757 & n2980) | (n1757 & n3035) | (n2980 & n3035);
  assign n3037 = n1642 | n1757;
  assign n3038 = n2980 | n3037;
  assign n1760 = ~n3036 & n3038;
  assign n1761 = x24 & x40;
  assign n1762 = n1760 & n1761;
  assign n1763 = n1760 | n1761;
  assign n1764 = ~n1762 & n1763;
  assign n3039 = n1649 & n1764;
  assign n3040 = (n1764 & n2985) | (n1764 & n3039) | (n2985 & n3039);
  assign n3041 = n1649 | n1764;
  assign n3042 = n2985 | n3041;
  assign n1767 = ~n3040 & n3042;
  assign n1768 = x23 & x41;
  assign n1769 = n1767 & n1768;
  assign n1770 = n1767 | n1768;
  assign n1771 = ~n1769 & n1770;
  assign n3043 = n1656 & n1771;
  assign n3044 = (n1771 & n2990) | (n1771 & n3043) | (n2990 & n3043);
  assign n3045 = n1656 | n1771;
  assign n3046 = n2990 | n3045;
  assign n1774 = ~n3044 & n3046;
  assign n1775 = x22 & x42;
  assign n1776 = n1774 & n1775;
  assign n1777 = n1774 | n1775;
  assign n1778 = ~n1776 & n1777;
  assign n1779 = n2998 & n1778;
  assign n1780 = n2998 | n1778;
  assign n1781 = ~n1779 & n1780;
  assign n1782 = x21 & x43;
  assign n1783 = n1781 & n1782;
  assign n1784 = n1781 | n1782;
  assign n1785 = ~n1783 & n1784;
  assign n1786 = n1704 & n1785;
  assign n1787 = n1704 | n1785;
  assign n1788 = ~n1786 & n1787;
  assign n1789 = x20 & x44;
  assign n1790 = n1788 & n1789;
  assign n1791 = n1788 | n1789;
  assign n1792 = ~n1790 & n1791;
  assign n1793 = n3611 & n1792;
  assign n1794 = n3611 | n1792;
  assign n1795 = ~n1793 & n1794;
  assign n1796 = x19 & x45;
  assign n1797 = n1795 & n1796;
  assign n1798 = n1795 | n1796;
  assign n1799 = ~n1797 & n1798;
  assign n1800 = n2996 & n1799;
  assign n1801 = n2996 | n1799;
  assign n1802 = ~n1800 & n1801;
  assign n1803 = x18 & x46;
  assign n1804 = n1802 & n1803;
  assign n1805 = n1802 | n1803;
  assign n1806 = ~n1804 & n1805;
  assign n1807 = n2994 & n1806;
  assign n1808 = n2994 | n1806;
  assign n1809 = ~n1807 & n1808;
  assign n1810 = x17 & x47;
  assign n1811 = n1809 & n1810;
  assign n1812 = n1809 | n1810;
  assign n1813 = ~n1811 & n1812;
  assign n1814 = n1698 & n1813;
  assign n1815 = n1698 | n1813;
  assign n1816 = ~n1814 & n1815;
  assign n3919 = n1697 | n1810;
  assign n3920 = (n1696 & n1810) | (n1696 & n3919) | (n1810 & n3919);
  assign n3639 = (n1698 & n1809) | (n1698 & n3920) | (n1809 & n3920);
  assign n3048 = (n1811 & n1813) | (n1811 & n3639) | (n1813 & n3639);
  assign n3049 = n1804 | n2994;
  assign n3050 = (n1804 & n1806) | (n1804 & n3049) | (n1806 & n3049);
  assign n3051 = n1797 | n2996;
  assign n3052 = (n1797 & n1799) | (n1797 & n3051) | (n1799 & n3051);
  assign n3640 = n1790 | n3611;
  assign n3641 = (n1790 & n1792) | (n1790 & n3640) | (n1792 & n3640);
  assign n3053 = n1783 | n1785;
  assign n3054 = (n1704 & n1783) | (n1704 & n3053) | (n1783 & n3053);
  assign n3055 = n1776 | n1778;
  assign n3056 = (n1776 & n2998) | (n1776 & n3055) | (n2998 & n3055);
  assign n3058 = n1741 | n1743;
  assign n3642 = n1628 | n1741;
  assign n3643 = (n1741 & n1743) | (n1741 & n3642) | (n1743 & n3642);
  assign n3644 = (n2971 & n3058) | (n2971 & n3643) | (n3058 & n3643);
  assign n3645 = (n1630 & n3058) | (n1630 & n3643) | (n3058 & n3643);
  assign n3646 = (n2935 & n3644) | (n2935 & n3645) | (n3644 & n3645);
  assign n1831 = x31 & x34;
  assign n1832 = n3625 & n1831;
  assign n1833 = n3625 | n1831;
  assign n1834 = ~n1832 & n1833;
  assign n3647 = n1720 | n1722;
  assign n3648 = (n1720 & n3004) | (n1720 & n3647) | (n3004 & n3647);
  assign n3065 = n1834 & n3648;
  assign n3649 = n1607 | n1720;
  assign n3650 = (n1720 & n1722) | (n1720 & n3649) | (n1722 & n3649);
  assign n3066 = n1834 & n3650;
  assign n3067 = (n3591 & n3065) | (n3591 & n3066) | (n3065 & n3066);
  assign n3068 = n1834 | n3648;
  assign n3069 = n1834 | n3650;
  assign n3070 = (n3591 & n3068) | (n3591 & n3069) | (n3068 & n3069);
  assign n1837 = ~n3067 & n3070;
  assign n1838 = x30 & x35;
  assign n1839 = n1837 & n1838;
  assign n1840 = n1837 | n1838;
  assign n1841 = ~n1839 & n1840;
  assign n3060 = n1727 | n1729;
  assign n3071 = n1841 & n3060;
  assign n3072 = n1727 & n1841;
  assign n3073 = (n3616 & n3071) | (n3616 & n3072) | (n3071 & n3072);
  assign n3074 = n1841 | n3060;
  assign n3075 = n1727 | n1841;
  assign n3076 = (n3616 & n3074) | (n3616 & n3075) | (n3074 & n3075);
  assign n1844 = ~n3073 & n3076;
  assign n1845 = x29 & x36;
  assign n1846 = n1844 & n1845;
  assign n1847 = n1844 | n1845;
  assign n1848 = ~n1846 & n1847;
  assign n3077 = n1734 & n1848;
  assign n3651 = (n1848 & n3022) | (n1848 & n3077) | (n3022 & n3077);
  assign n3652 = (n1848 & n3021) | (n1848 & n3077) | (n3021 & n3077);
  assign n3653 = (n3584 & n3651) | (n3584 & n3652) | (n3651 & n3652);
  assign n3079 = n1734 | n1848;
  assign n3654 = n3022 | n3079;
  assign n3655 = n3021 | n3079;
  assign n3656 = (n3584 & n3654) | (n3584 & n3655) | (n3654 & n3655);
  assign n1851 = ~n3653 & n3656;
  assign n1852 = x28 & x37;
  assign n1853 = n1851 & n1852;
  assign n1854 = n1851 | n1852;
  assign n1855 = ~n1853 & n1854;
  assign n1856 = n3646 & n1855;
  assign n1857 = n3646 | n1855;
  assign n1858 = ~n1856 & n1857;
  assign n1859 = x27 & x38;
  assign n1860 = n1858 & n1859;
  assign n1861 = n1858 | n1859;
  assign n1862 = ~n1860 & n1861;
  assign n3081 = n1748 & n1862;
  assign n3082 = (n1862 & n3032) | (n1862 & n3081) | (n3032 & n3081);
  assign n3083 = n1748 | n1862;
  assign n3084 = n3032 | n3083;
  assign n1865 = ~n3082 & n3084;
  assign n1866 = x26 & x39;
  assign n1867 = n1865 & n1866;
  assign n1868 = n1865 | n1866;
  assign n1869 = ~n1867 & n1868;
  assign n3085 = n1755 & n1869;
  assign n3086 = (n1869 & n3036) | (n1869 & n3085) | (n3036 & n3085);
  assign n3087 = n1755 | n1869;
  assign n3088 = n3036 | n3087;
  assign n1872 = ~n3086 & n3088;
  assign n1873 = x25 & x40;
  assign n1874 = n1872 & n1873;
  assign n1875 = n1872 | n1873;
  assign n1876 = ~n1874 & n1875;
  assign n3089 = n1762 & n1876;
  assign n3090 = (n1876 & n3040) | (n1876 & n3089) | (n3040 & n3089);
  assign n3091 = n1762 | n1876;
  assign n3092 = n3040 | n3091;
  assign n1879 = ~n3090 & n3092;
  assign n1880 = x24 & x41;
  assign n1881 = n1879 & n1880;
  assign n1882 = n1879 | n1880;
  assign n1883 = ~n1881 & n1882;
  assign n3093 = n1769 & n1883;
  assign n3094 = (n1883 & n3044) | (n1883 & n3093) | (n3044 & n3093);
  assign n3095 = n1769 | n1883;
  assign n3096 = n3044 | n3095;
  assign n1886 = ~n3094 & n3096;
  assign n1887 = x23 & x42;
  assign n1888 = n1886 & n1887;
  assign n1889 = n1886 | n1887;
  assign n1890 = ~n1888 & n1889;
  assign n1891 = n3056 & n1890;
  assign n1892 = n3056 | n1890;
  assign n1893 = ~n1891 & n1892;
  assign n1894 = x22 & x43;
  assign n1895 = n1893 & n1894;
  assign n1896 = n1893 | n1894;
  assign n1897 = ~n1895 & n1896;
  assign n1898 = n3054 & n1897;
  assign n1899 = n3054 | n1897;
  assign n1900 = ~n1898 & n1899;
  assign n1901 = x21 & x44;
  assign n1902 = n1900 & n1901;
  assign n1903 = n1900 | n1901;
  assign n1904 = ~n1902 & n1903;
  assign n1905 = n3641 & n1904;
  assign n1906 = n3641 | n1904;
  assign n1907 = ~n1905 & n1906;
  assign n1908 = x20 & x45;
  assign n1909 = n1907 & n1908;
  assign n1910 = n1907 | n1908;
  assign n1911 = ~n1909 & n1910;
  assign n1912 = n3052 & n1911;
  assign n1913 = n3052 | n1911;
  assign n1914 = ~n1912 & n1913;
  assign n1915 = x19 & x46;
  assign n1916 = n1914 & n1915;
  assign n1917 = n1914 | n1915;
  assign n1918 = ~n1916 & n1917;
  assign n1919 = n3050 & n1918;
  assign n1920 = n3050 | n1918;
  assign n1921 = ~n1919 & n1920;
  assign n1922 = x18 & x47;
  assign n1923 = n1921 & n1922;
  assign n1924 = n1921 | n1922;
  assign n1925 = ~n1923 & n1924;
  assign n1926 = n3048 & n1925;
  assign n1927 = n3048 | n1925;
  assign n1928 = ~n1926 & n1927;
  assign n3097 = n1923 | n3048;
  assign n3098 = (n1923 & n1925) | (n1923 & n3097) | (n1925 & n3097);
  assign n3099 = n1916 | n3050;
  assign n3100 = (n1916 & n1918) | (n1916 & n3099) | (n1918 & n3099);
  assign n3101 = n1909 | n3052;
  assign n3102 = (n1909 & n1911) | (n1909 & n3101) | (n1911 & n3101);
  assign n3103 = n1902 | n1904;
  assign n3104 = (n3641 & n1902) | (n3641 & n3103) | (n1902 & n3103);
  assign n3105 = n1895 | n1897;
  assign n3106 = (n1895 & n3054) | (n1895 & n3105) | (n3054 & n3105);
  assign n3107 = n1888 | n1890;
  assign n3108 = (n1888 & n3056) | (n1888 & n3107) | (n3056 & n3107);
  assign n3112 = n1846 | n1848;
  assign n3657 = n1734 | n1846;
  assign n3658 = (n1846 & n1848) | (n1846 & n3657) | (n1848 & n3657);
  assign n3659 = (n3022 & n3112) | (n3022 & n3658) | (n3112 & n3658);
  assign n3660 = (n3021 & n3112) | (n3021 & n3658) | (n3112 & n3658);
  assign n3661 = (n3584 & n3659) | (n3584 & n3660) | (n3659 & n3660);
  assign n1943 = x31 & x35;
  assign n3666 = n1831 & n1943;
  assign n3667 = n3625 & n3666;
  assign n3921 = (n1834 & n1943) | (n1834 & n3667) | (n1943 & n3667);
  assign n3922 = n1943 & n3667;
  assign n3923 = (n3648 & n3921) | (n3648 & n3922) | (n3921 & n3922);
  assign n3924 = (n3650 & n3921) | (n3650 & n3922) | (n3921 & n3922);
  assign n3670 = (n3591 & n3923) | (n3591 & n3924) | (n3923 & n3924);
  assign n3671 = n1831 | n1943;
  assign n3672 = (n1943 & n3625) | (n1943 & n3671) | (n3625 & n3671);
  assign n3925 = n1834 | n3672;
  assign n3926 = (n3648 & n3672) | (n3648 & n3925) | (n3672 & n3925);
  assign n3927 = (n3650 & n3672) | (n3650 & n3925) | (n3672 & n3925);
  assign n3675 = (n3591 & n3926) | (n3591 & n3927) | (n3926 & n3927);
  assign n1946 = ~n3670 & n3675;
  assign n3662 = n1839 | n1841;
  assign n3663 = (n1839 & n3060) | (n1839 & n3662) | (n3060 & n3662);
  assign n3676 = n1946 & n3663;
  assign n3664 = n1727 | n1839;
  assign n3665 = (n1839 & n1841) | (n1839 & n3664) | (n1841 & n3664);
  assign n3677 = n1946 & n3665;
  assign n3678 = (n3616 & n3676) | (n3616 & n3677) | (n3676 & n3677);
  assign n3679 = n1946 | n3663;
  assign n3680 = n1946 | n3665;
  assign n3681 = (n3616 & n3679) | (n3616 & n3680) | (n3679 & n3680);
  assign n1949 = ~n3678 & n3681;
  assign n1950 = x30 & x36;
  assign n1951 = n1949 & n1950;
  assign n1952 = n1949 | n1950;
  assign n1953 = ~n1951 & n1952;
  assign n1954 = n3661 & n1953;
  assign n1955 = n3661 | n1953;
  assign n1956 = ~n1954 & n1955;
  assign n1957 = x29 & x37;
  assign n1958 = n1956 & n1957;
  assign n1959 = n1956 | n1957;
  assign n1960 = ~n1958 & n1959;
  assign n3109 = n1853 | n1855;
  assign n3121 = n1960 & n3109;
  assign n3122 = n1853 & n1960;
  assign n3123 = (n3646 & n3121) | (n3646 & n3122) | (n3121 & n3122);
  assign n3124 = n1960 | n3109;
  assign n3125 = n1853 | n1960;
  assign n3126 = (n3646 & n3124) | (n3646 & n3125) | (n3124 & n3125);
  assign n1963 = ~n3123 & n3126;
  assign n1964 = x28 & x38;
  assign n1965 = n1963 & n1964;
  assign n1966 = n1963 | n1964;
  assign n1967 = ~n1965 & n1966;
  assign n3127 = n1860 & n1967;
  assign n3682 = (n1967 & n3081) | (n1967 & n3127) | (n3081 & n3127);
  assign n3683 = (n1862 & n1967) | (n1862 & n3127) | (n1967 & n3127);
  assign n3684 = (n3032 & n3682) | (n3032 & n3683) | (n3682 & n3683);
  assign n3129 = n1860 | n1967;
  assign n3685 = n3081 | n3129;
  assign n3686 = n1862 | n3129;
  assign n3687 = (n3032 & n3685) | (n3032 & n3686) | (n3685 & n3686);
  assign n1970 = ~n3684 & n3687;
  assign n1971 = x27 & x39;
  assign n1972 = n1970 & n1971;
  assign n1973 = n1970 | n1971;
  assign n1974 = ~n1972 & n1973;
  assign n3131 = n1867 & n1974;
  assign n3132 = (n1974 & n3086) | (n1974 & n3131) | (n3086 & n3131);
  assign n3133 = n1867 | n1974;
  assign n3134 = n3086 | n3133;
  assign n1977 = ~n3132 & n3134;
  assign n1978 = x26 & x40;
  assign n1979 = n1977 & n1978;
  assign n1980 = n1977 | n1978;
  assign n1981 = ~n1979 & n1980;
  assign n3135 = n1874 & n1981;
  assign n3136 = (n1981 & n3090) | (n1981 & n3135) | (n3090 & n3135);
  assign n3137 = n1874 | n1981;
  assign n3138 = n3090 | n3137;
  assign n1984 = ~n3136 & n3138;
  assign n1985 = x25 & x41;
  assign n1986 = n1984 & n1985;
  assign n1987 = n1984 | n1985;
  assign n1988 = ~n1986 & n1987;
  assign n3139 = n1881 & n1988;
  assign n3140 = (n1988 & n3094) | (n1988 & n3139) | (n3094 & n3139);
  assign n3141 = n1881 | n1988;
  assign n3142 = n3094 | n3141;
  assign n1991 = ~n3140 & n3142;
  assign n1992 = x24 & x42;
  assign n1993 = n1991 & n1992;
  assign n1994 = n1991 | n1992;
  assign n1995 = ~n1993 & n1994;
  assign n1996 = n3108 & n1995;
  assign n1997 = n3108 | n1995;
  assign n1998 = ~n1996 & n1997;
  assign n1999 = x23 & x43;
  assign n2000 = n1998 & n1999;
  assign n2001 = n1998 | n1999;
  assign n2002 = ~n2000 & n2001;
  assign n2003 = n3106 & n2002;
  assign n2004 = n3106 | n2002;
  assign n2005 = ~n2003 & n2004;
  assign n2006 = x22 & x44;
  assign n2007 = n2005 & n2006;
  assign n2008 = n2005 | n2006;
  assign n2009 = ~n2007 & n2008;
  assign n2010 = n3104 & n2009;
  assign n2011 = n3104 | n2009;
  assign n2012 = ~n2010 & n2011;
  assign n2013 = x21 & x45;
  assign n2014 = n2012 & n2013;
  assign n2015 = n2012 | n2013;
  assign n2016 = ~n2014 & n2015;
  assign n2017 = n3102 & n2016;
  assign n2018 = n3102 | n2016;
  assign n2019 = ~n2017 & n2018;
  assign n2020 = x20 & x46;
  assign n2021 = n2019 & n2020;
  assign n2022 = n2019 | n2020;
  assign n2023 = ~n2021 & n2022;
  assign n2024 = n3100 & n2023;
  assign n2025 = n3100 | n2023;
  assign n2026 = ~n2024 & n2025;
  assign n2027 = x19 & x47;
  assign n2028 = n2026 & n2027;
  assign n2029 = n2026 | n2027;
  assign n2030 = ~n2028 & n2029;
  assign n2031 = n3098 & n2030;
  assign n2032 = n3098 | n2030;
  assign n2033 = ~n2031 & n2032;
  assign n2034 = n2028 | n2031;
  assign n2035 = n2021 | n2024;
  assign n2036 = n2014 | n2017;
  assign n3143 = n2007 | n2009;
  assign n3144 = (n2007 & n3104) | (n2007 & n3143) | (n3104 & n3143);
  assign n3145 = n2000 | n2002;
  assign n3146 = (n2000 & n3106) | (n2000 & n3145) | (n3106 & n3145);
  assign n3147 = n1993 | n1995;
  assign n3148 = (n1993 & n3108) | (n1993 & n3147) | (n3108 & n3147);
  assign n3150 = n1965 | n1967;
  assign n3688 = n1860 | n1965;
  assign n3689 = (n1965 & n1967) | (n1965 & n3688) | (n1967 & n3688);
  assign n3690 = (n3081 & n3150) | (n3081 & n3689) | (n3150 & n3689);
  assign n3691 = (n1862 & n3150) | (n1862 & n3689) | (n3150 & n3689);
  assign n3692 = (n3032 & n3690) | (n3032 & n3691) | (n3690 & n3691);
  assign n2047 = x31 & x36;
  assign n3928 = n2047 & n3923;
  assign n3929 = n2047 & n3924;
  assign n3930 = (n3591 & n3928) | (n3591 & n3929) | (n3928 & n3929);
  assign n3694 = (n1946 & n2047) | (n1946 & n3930) | (n2047 & n3930);
  assign n3695 = (n3930 & n3663) | (n3930 & n3694) | (n3663 & n3694);
  assign n3696 = (n3930 & n3665) | (n3930 & n3694) | (n3665 & n3694);
  assign n3697 = (n3616 & n3695) | (n3616 & n3696) | (n3695 & n3696);
  assign n3931 = n2047 | n3923;
  assign n3932 = n2047 | n3924;
  assign n3933 = (n3591 & n3931) | (n3591 & n3932) | (n3931 & n3932);
  assign n3699 = n1946 | n3933;
  assign n3700 = (n3933 & n3663) | (n3933 & n3699) | (n3663 & n3699);
  assign n3701 = (n3933 & n3665) | (n3933 & n3699) | (n3665 & n3699);
  assign n3702 = (n3616 & n3700) | (n3616 & n3701) | (n3700 & n3701);
  assign n2050 = ~n3697 & n3702;
  assign n3163 = n1951 & n2050;
  assign n3703 = (n1953 & n2050) | (n1953 & n3163) | (n2050 & n3163);
  assign n3164 = (n3661 & n3703) | (n3661 & n3163) | (n3703 & n3163);
  assign n3166 = n1951 | n2050;
  assign n3704 = n1953 | n3166;
  assign n3167 = (n3661 & n3704) | (n3661 & n3166) | (n3704 & n3166);
  assign n2053 = ~n3164 & n3167;
  assign n2054 = x30 & x37;
  assign n2055 = n2053 & n2054;
  assign n2056 = n2053 | n2054;
  assign n2057 = ~n2055 & n2056;
  assign n3168 = n1958 & n2057;
  assign n3705 = (n2057 & n3122) | (n2057 & n3168) | (n3122 & n3168);
  assign n3706 = (n2057 & n3121) | (n2057 & n3168) | (n3121 & n3168);
  assign n3707 = (n3646 & n3705) | (n3646 & n3706) | (n3705 & n3706);
  assign n3170 = n1958 | n2057;
  assign n3708 = n3122 | n3170;
  assign n3709 = n3121 | n3170;
  assign n3710 = (n3646 & n3708) | (n3646 & n3709) | (n3708 & n3709);
  assign n2060 = ~n3707 & n3710;
  assign n2061 = x29 & x38;
  assign n2062 = n2060 & n2061;
  assign n2063 = n2060 | n2061;
  assign n2064 = ~n2062 & n2063;
  assign n2065 = n3692 & n2064;
  assign n2066 = n3692 | n2064;
  assign n2067 = ~n2065 & n2066;
  assign n2068 = x28 & x39;
  assign n2069 = n2067 & n2068;
  assign n2070 = n2067 | n2068;
  assign n2071 = ~n2069 & n2070;
  assign n3172 = n1972 & n2071;
  assign n3173 = (n2071 & n3132) | (n2071 & n3172) | (n3132 & n3172);
  assign n3174 = n1972 | n2071;
  assign n3175 = n3132 | n3174;
  assign n2074 = ~n3173 & n3175;
  assign n2075 = x27 & x40;
  assign n2076 = n2074 & n2075;
  assign n2077 = n2074 | n2075;
  assign n2078 = ~n2076 & n2077;
  assign n3176 = n1979 & n2078;
  assign n3177 = (n2078 & n3136) | (n2078 & n3176) | (n3136 & n3176);
  assign n3178 = n1979 | n2078;
  assign n3179 = n3136 | n3178;
  assign n2081 = ~n3177 & n3179;
  assign n2082 = x26 & x41;
  assign n2083 = n2081 & n2082;
  assign n2084 = n2081 | n2082;
  assign n2085 = ~n2083 & n2084;
  assign n3180 = n1986 & n2085;
  assign n3181 = (n2085 & n3140) | (n2085 & n3180) | (n3140 & n3180);
  assign n3182 = n1986 | n2085;
  assign n3183 = n3140 | n3182;
  assign n2088 = ~n3181 & n3183;
  assign n2089 = x25 & x42;
  assign n2090 = n2088 & n2089;
  assign n2091 = n2088 | n2089;
  assign n2092 = ~n2090 & n2091;
  assign n2093 = n3148 & n2092;
  assign n2094 = n3148 | n2092;
  assign n2095 = ~n2093 & n2094;
  assign n2096 = x24 & x43;
  assign n2097 = n2095 & n2096;
  assign n2098 = n2095 | n2096;
  assign n2099 = ~n2097 & n2098;
  assign n2100 = n3146 & n2099;
  assign n2101 = n3146 | n2099;
  assign n2102 = ~n2100 & n2101;
  assign n2103 = x23 & x44;
  assign n2104 = n2102 & n2103;
  assign n2105 = n2102 | n2103;
  assign n2106 = ~n2104 & n2105;
  assign n2107 = n3144 & n2106;
  assign n2108 = n3144 | n2106;
  assign n2109 = ~n2107 & n2108;
  assign n2110 = x22 & x45;
  assign n2111 = n2109 & n2110;
  assign n2112 = n2109 | n2110;
  assign n2113 = ~n2111 & n2112;
  assign n2114 = n2036 & n2113;
  assign n2115 = n2036 | n2113;
  assign n2116 = ~n2114 & n2115;
  assign n2117 = x21 & x46;
  assign n2118 = n2116 & n2117;
  assign n2119 = n2116 | n2117;
  assign n2120 = ~n2118 & n2119;
  assign n2121 = n2035 & n2120;
  assign n2122 = n2035 | n2120;
  assign n2123 = ~n2121 & n2122;
  assign n2124 = x20 & x47;
  assign n2125 = n2123 & n2124;
  assign n2126 = n2123 | n2124;
  assign n2127 = ~n2125 & n2126;
  assign n2128 = n2034 & n2127;
  assign n2129 = n2034 | n2127;
  assign n2130 = ~n2128 & n2129;
  assign n2131 = n2125 | n2128;
  assign n2132 = n2118 | n2121;
  assign n3184 = n2111 | n2113;
  assign n3185 = (n2036 & n2111) | (n2036 & n3184) | (n2111 & n3184);
  assign n3186 = n2104 | n2106;
  assign n3187 = (n2104 & n3144) | (n2104 & n3186) | (n3144 & n3186);
  assign n3188 = n2097 | n2099;
  assign n3189 = (n2097 & n3146) | (n2097 & n3188) | (n3146 & n3188);
  assign n3190 = n2090 | n2092;
  assign n3191 = (n2090 & n3148) | (n2090 & n3190) | (n3148 & n3190);
  assign n3195 = n2055 | n2057;
  assign n3711 = n1958 | n2055;
  assign n3712 = (n2055 & n2057) | (n2055 & n3711) | (n2057 & n3711);
  assign n3713 = (n3122 & n3195) | (n3122 & n3712) | (n3195 & n3712);
  assign n3714 = (n3121 & n3195) | (n3121 & n3712) | (n3195 & n3712);
  assign n3715 = (n3646 & n3713) | (n3646 & n3714) | (n3713 & n3714);
  assign n2143 = x31 & x37;
  assign n3197 = n2143 & n3697;
  assign n3716 = (n2143 & n3197) | (n2143 & n3703) | (n3197 & n3703);
  assign n3934 = (n2050 & n2143) | (n2050 & n3197) | (n2143 & n3197);
  assign n3935 = n2143 & n3197;
  assign n3936 = (n1951 & n3934) | (n1951 & n3935) | (n3934 & n3935);
  assign n3718 = (n3661 & n3716) | (n3661 & n3936) | (n3716 & n3936);
  assign n3199 = n2143 | n3697;
  assign n3719 = n3199 | n3703;
  assign n3937 = n2050 | n3199;
  assign n3938 = (n1951 & n3199) | (n1951 & n3937) | (n3199 & n3937);
  assign n3721 = (n3661 & n3719) | (n3661 & n3938) | (n3719 & n3938);
  assign n2146 = ~n3718 & n3721;
  assign n2147 = n3715 & n2146;
  assign n2148 = n3715 | n2146;
  assign n2149 = ~n2147 & n2148;
  assign n2150 = x30 & x38;
  assign n2151 = n2149 & n2150;
  assign n2152 = n2149 | n2150;
  assign n2153 = ~n2151 & n2152;
  assign n3192 = n2062 | n2064;
  assign n3201 = n2153 & n3192;
  assign n3202 = n2062 & n2153;
  assign n3203 = (n3692 & n3201) | (n3692 & n3202) | (n3201 & n3202);
  assign n3204 = n2153 | n3192;
  assign n3205 = n2062 | n2153;
  assign n3206 = (n3692 & n3204) | (n3692 & n3205) | (n3204 & n3205);
  assign n2156 = ~n3203 & n3206;
  assign n2157 = x29 & x39;
  assign n2158 = n2156 & n2157;
  assign n2159 = n2156 | n2157;
  assign n2160 = ~n2158 & n2159;
  assign n3207 = n2069 & n2160;
  assign n3722 = (n2160 & n3172) | (n2160 & n3207) | (n3172 & n3207);
  assign n3723 = (n2071 & n2160) | (n2071 & n3207) | (n2160 & n3207);
  assign n3724 = (n3132 & n3722) | (n3132 & n3723) | (n3722 & n3723);
  assign n3209 = n2069 | n2160;
  assign n3725 = n3172 | n3209;
  assign n3726 = n2071 | n3209;
  assign n3727 = (n3132 & n3725) | (n3132 & n3726) | (n3725 & n3726);
  assign n2163 = ~n3724 & n3727;
  assign n2164 = x28 & x40;
  assign n2165 = n2163 & n2164;
  assign n2166 = n2163 | n2164;
  assign n2167 = ~n2165 & n2166;
  assign n3211 = n2076 & n2167;
  assign n3212 = (n2167 & n3177) | (n2167 & n3211) | (n3177 & n3211);
  assign n3213 = n2076 | n2167;
  assign n3214 = n3177 | n3213;
  assign n2170 = ~n3212 & n3214;
  assign n2171 = x27 & x41;
  assign n2172 = n2170 & n2171;
  assign n2173 = n2170 | n2171;
  assign n2174 = ~n2172 & n2173;
  assign n3215 = n2083 & n2174;
  assign n3216 = (n2174 & n3181) | (n2174 & n3215) | (n3181 & n3215);
  assign n3217 = n2083 | n2174;
  assign n3218 = n3181 | n3217;
  assign n2177 = ~n3216 & n3218;
  assign n2178 = x26 & x42;
  assign n2179 = n2177 & n2178;
  assign n2180 = n2177 | n2178;
  assign n2181 = ~n2179 & n2180;
  assign n2182 = n3191 & n2181;
  assign n2183 = n3191 | n2181;
  assign n2184 = ~n2182 & n2183;
  assign n2185 = x25 & x43;
  assign n2186 = n2184 & n2185;
  assign n2187 = n2184 | n2185;
  assign n2188 = ~n2186 & n2187;
  assign n2189 = n3189 & n2188;
  assign n2190 = n3189 | n2188;
  assign n2191 = ~n2189 & n2190;
  assign n2192 = x24 & x44;
  assign n2193 = n2191 & n2192;
  assign n2194 = n2191 | n2192;
  assign n2195 = ~n2193 & n2194;
  assign n2196 = n3187 & n2195;
  assign n2197 = n3187 | n2195;
  assign n2198 = ~n2196 & n2197;
  assign n2199 = x23 & x45;
  assign n2200 = n2198 & n2199;
  assign n2201 = n2198 | n2199;
  assign n2202 = ~n2200 & n2201;
  assign n2203 = n3185 & n2202;
  assign n2204 = n3185 | n2202;
  assign n2205 = ~n2203 & n2204;
  assign n2206 = x22 & x46;
  assign n2207 = n2205 & n2206;
  assign n2208 = n2205 | n2206;
  assign n2209 = ~n2207 & n2208;
  assign n2210 = n2132 & n2209;
  assign n2211 = n2132 | n2209;
  assign n2212 = ~n2210 & n2211;
  assign n2213 = x21 & x47;
  assign n2214 = n2212 & n2213;
  assign n2215 = n2212 | n2213;
  assign n2216 = ~n2214 & n2215;
  assign n2217 = n2131 & n2216;
  assign n2218 = n2131 | n2216;
  assign n2219 = ~n2217 & n2218;
  assign n2220 = n2214 | n2217;
  assign n3219 = n2207 | n2209;
  assign n3220 = (n2132 & n2207) | (n2132 & n3219) | (n2207 & n3219);
  assign n3221 = n2200 | n2202;
  assign n3222 = (n2200 & n3185) | (n2200 & n3221) | (n3185 & n3221);
  assign n3223 = n2193 | n2195;
  assign n3224 = (n2193 & n3187) | (n2193 & n3223) | (n3187 & n3223);
  assign n3225 = n2186 | n2188;
  assign n3226 = (n2186 & n3189) | (n2186 & n3225) | (n3189 & n3225);
  assign n3227 = n2179 | n2181;
  assign n3228 = (n2179 & n3191) | (n2179 & n3227) | (n3191 & n3227);
  assign n3230 = n2158 | n2160;
  assign n3728 = n2069 | n2158;
  assign n3729 = (n2158 & n2160) | (n2158 & n3728) | (n2160 & n3728);
  assign n3730 = (n3172 & n3230) | (n3172 & n3729) | (n3230 & n3729);
  assign n3731 = (n2071 & n3230) | (n2071 & n3729) | (n3230 & n3729);
  assign n3732 = (n3132 & n3730) | (n3132 & n3731) | (n3730 & n3731);
  assign n2231 = x31 & x38;
  assign n3941 = n2231 & n3197;
  assign n3942 = n2143 & n2231;
  assign n3943 = (n3703 & n3941) | (n3703 & n3942) | (n3941 & n3942);
  assign n3939 = n2231 & n3936;
  assign n3940 = (n3661 & n3943) | (n3661 & n3939) | (n3943 & n3939);
  assign n3734 = (n2146 & n2231) | (n2146 & n3940) | (n2231 & n3940);
  assign n3736 = n2231 & n3936;
  assign n3737 = (n3661 & n3943) | (n3661 & n3736) | (n3943 & n3736);
  assign n3236 = (n3715 & n3734) | (n3715 & n3737) | (n3734 & n3737);
  assign n3946 = n2231 | n3197;
  assign n3947 = n2143 | n2231;
  assign n3948 = (n3703 & n3946) | (n3703 & n3947) | (n3946 & n3947);
  assign n3944 = n2231 | n3936;
  assign n3945 = (n3661 & n3948) | (n3661 & n3944) | (n3948 & n3944);
  assign n3739 = n2146 | n3945;
  assign n3741 = n2231 | n3936;
  assign n3742 = (n3661 & n3948) | (n3661 & n3741) | (n3948 & n3741);
  assign n3239 = (n3715 & n3739) | (n3715 & n3742) | (n3739 & n3742);
  assign n2234 = ~n3236 & n3239;
  assign n3240 = n2151 & n2234;
  assign n3743 = (n2234 & n3202) | (n2234 & n3240) | (n3202 & n3240);
  assign n3744 = (n2234 & n3201) | (n2234 & n3240) | (n3201 & n3240);
  assign n3745 = (n3692 & n3743) | (n3692 & n3744) | (n3743 & n3744);
  assign n3242 = n2151 | n2234;
  assign n3746 = n3202 | n3242;
  assign n3747 = n3201 | n3242;
  assign n3748 = (n3692 & n3746) | (n3692 & n3747) | (n3746 & n3747);
  assign n2237 = ~n3745 & n3748;
  assign n2238 = x30 & x39;
  assign n2239 = n2237 & n2238;
  assign n2240 = n2237 | n2238;
  assign n2241 = ~n2239 & n2240;
  assign n2242 = n3732 & n2241;
  assign n2243 = n3732 | n2241;
  assign n2244 = ~n2242 & n2243;
  assign n2245 = x29 & x40;
  assign n2246 = n2244 & n2245;
  assign n2247 = n2244 | n2245;
  assign n2248 = ~n2246 & n2247;
  assign n3244 = n2165 & n2248;
  assign n3245 = (n2248 & n3212) | (n2248 & n3244) | (n3212 & n3244);
  assign n3246 = n2165 | n2248;
  assign n3247 = n3212 | n3246;
  assign n2251 = ~n3245 & n3247;
  assign n2252 = x28 & x41;
  assign n2253 = n2251 & n2252;
  assign n2254 = n2251 | n2252;
  assign n2255 = ~n2253 & n2254;
  assign n3248 = n2172 & n2255;
  assign n3249 = (n2255 & n3216) | (n2255 & n3248) | (n3216 & n3248);
  assign n3250 = n2172 | n2255;
  assign n3251 = n3216 | n3250;
  assign n2258 = ~n3249 & n3251;
  assign n2259 = x27 & x42;
  assign n2260 = n2258 & n2259;
  assign n2261 = n2258 | n2259;
  assign n2262 = ~n2260 & n2261;
  assign n2263 = n3228 & n2262;
  assign n2264 = n3228 | n2262;
  assign n2265 = ~n2263 & n2264;
  assign n2266 = x26 & x43;
  assign n2267 = n2265 & n2266;
  assign n2268 = n2265 | n2266;
  assign n2269 = ~n2267 & n2268;
  assign n2270 = n3226 & n2269;
  assign n2271 = n3226 | n2269;
  assign n2272 = ~n2270 & n2271;
  assign n2273 = x25 & x44;
  assign n2274 = n2272 & n2273;
  assign n2275 = n2272 | n2273;
  assign n2276 = ~n2274 & n2275;
  assign n2277 = n3224 & n2276;
  assign n2278 = n3224 | n2276;
  assign n2279 = ~n2277 & n2278;
  assign n2280 = x24 & x45;
  assign n2281 = n2279 & n2280;
  assign n2282 = n2279 | n2280;
  assign n2283 = ~n2281 & n2282;
  assign n2284 = n3222 & n2283;
  assign n2285 = n3222 | n2283;
  assign n2286 = ~n2284 & n2285;
  assign n2287 = x23 & x46;
  assign n2288 = n2286 & n2287;
  assign n2289 = n2286 | n2287;
  assign n2290 = ~n2288 & n2289;
  assign n2291 = n3220 & n2290;
  assign n2292 = n3220 | n2290;
  assign n2293 = ~n2291 & n2292;
  assign n2294 = x22 & x47;
  assign n2295 = n2293 & n2294;
  assign n2296 = n2293 | n2294;
  assign n2297 = ~n2295 & n2296;
  assign n2298 = n2220 & n2297;
  assign n2299 = n2220 | n2297;
  assign n2300 = ~n2298 & n2299;
  assign n3252 = n2295 | n2297;
  assign n3253 = (n2220 & n2295) | (n2220 & n3252) | (n2295 & n3252);
  assign n3254 = n2288 | n2290;
  assign n3255 = (n2288 & n3220) | (n2288 & n3254) | (n3220 & n3254);
  assign n3256 = n2281 | n2283;
  assign n3257 = (n2281 & n3222) | (n2281 & n3256) | (n3222 & n3256);
  assign n3258 = n2274 | n2276;
  assign n3259 = (n2274 & n3224) | (n2274 & n3258) | (n3224 & n3258);
  assign n3260 = n2267 | n2269;
  assign n3261 = (n2267 & n3226) | (n2267 & n3260) | (n3226 & n3260);
  assign n3262 = n2260 | n2262;
  assign n3263 = (n2260 & n3228) | (n2260 & n3262) | (n3228 & n3262);
  assign n2311 = x31 & x39;
  assign n3267 = n2234 | n3236;
  assign n3749 = (n2151 & n3236) | (n2151 & n3267) | (n3236 & n3267);
  assign n3269 = n2311 & n3749;
  assign n3949 = n2311 & n3734;
  assign n3950 = n2311 & n3737;
  assign n3951 = (n3715 & n3949) | (n3715 & n3950) | (n3949 & n3950);
  assign n3751 = (n2234 & n2311) | (n2234 & n3951) | (n2311 & n3951);
  assign n3752 = (n3202 & n3269) | (n3202 & n3751) | (n3269 & n3751);
  assign n3753 = (n3201 & n3269) | (n3201 & n3751) | (n3269 & n3751);
  assign n3754 = (n3692 & n3752) | (n3692 & n3753) | (n3752 & n3753);
  assign n3272 = n2311 | n3749;
  assign n3952 = n2311 | n3734;
  assign n3953 = n2311 | n3737;
  assign n3954 = (n3715 & n3952) | (n3715 & n3953) | (n3952 & n3953);
  assign n3756 = n2234 | n3954;
  assign n3757 = (n3202 & n3272) | (n3202 & n3756) | (n3272 & n3756);
  assign n3758 = (n3201 & n3272) | (n3201 & n3756) | (n3272 & n3756);
  assign n3759 = (n3692 & n3757) | (n3692 & n3758) | (n3757 & n3758);
  assign n2314 = ~n3754 & n3759;
  assign n3276 = n2239 & n2314;
  assign n3760 = (n2241 & n2314) | (n2241 & n3276) | (n2314 & n3276);
  assign n3277 = (n3732 & n3760) | (n3732 & n3276) | (n3760 & n3276);
  assign n3279 = n2239 | n2314;
  assign n3761 = n2241 | n3279;
  assign n3280 = (n3732 & n3761) | (n3732 & n3279) | (n3761 & n3279);
  assign n2317 = ~n3277 & n3280;
  assign n2318 = x30 & x40;
  assign n2319 = n2317 & n2318;
  assign n2320 = n2317 | n2318;
  assign n2321 = ~n2319 & n2320;
  assign n3281 = n2246 & n2321;
  assign n3762 = (n2321 & n3244) | (n2321 & n3281) | (n3244 & n3281);
  assign n3763 = (n2248 & n2321) | (n2248 & n3281) | (n2321 & n3281);
  assign n3764 = (n3212 & n3762) | (n3212 & n3763) | (n3762 & n3763);
  assign n3283 = n2246 | n2321;
  assign n3765 = n3244 | n3283;
  assign n3766 = n2248 | n3283;
  assign n3767 = (n3212 & n3765) | (n3212 & n3766) | (n3765 & n3766);
  assign n2324 = ~n3764 & n3767;
  assign n2325 = x29 & x41;
  assign n2326 = n2324 & n2325;
  assign n2327 = n2324 | n2325;
  assign n2328 = ~n2326 & n2327;
  assign n3285 = n2253 & n2328;
  assign n3286 = (n2328 & n3249) | (n2328 & n3285) | (n3249 & n3285);
  assign n3287 = n2253 | n2328;
  assign n3288 = n3249 | n3287;
  assign n2331 = ~n3286 & n3288;
  assign n2332 = x28 & x42;
  assign n2333 = n2331 & n2332;
  assign n2334 = n2331 | n2332;
  assign n2335 = ~n2333 & n2334;
  assign n2336 = n3263 & n2335;
  assign n2337 = n3263 | n2335;
  assign n2338 = ~n2336 & n2337;
  assign n2339 = x27 & x43;
  assign n2340 = n2338 & n2339;
  assign n2341 = n2338 | n2339;
  assign n2342 = ~n2340 & n2341;
  assign n2343 = n3261 & n2342;
  assign n2344 = n3261 | n2342;
  assign n2345 = ~n2343 & n2344;
  assign n2346 = x26 & x44;
  assign n2347 = n2345 & n2346;
  assign n2348 = n2345 | n2346;
  assign n2349 = ~n2347 & n2348;
  assign n2350 = n3259 & n2349;
  assign n2351 = n3259 | n2349;
  assign n2352 = ~n2350 & n2351;
  assign n2353 = x25 & x45;
  assign n2354 = n2352 & n2353;
  assign n2355 = n2352 | n2353;
  assign n2356 = ~n2354 & n2355;
  assign n2357 = n3257 & n2356;
  assign n2358 = n3257 | n2356;
  assign n2359 = ~n2357 & n2358;
  assign n2360 = x24 & x46;
  assign n2361 = n2359 & n2360;
  assign n2362 = n2359 | n2360;
  assign n2363 = ~n2361 & n2362;
  assign n2364 = n3255 & n2363;
  assign n2365 = n3255 | n2363;
  assign n2366 = ~n2364 & n2365;
  assign n2367 = x23 & x47;
  assign n2368 = n2366 & n2367;
  assign n2369 = n2366 | n2367;
  assign n2370 = ~n2368 & n2369;
  assign n2371 = n3253 & n2370;
  assign n2372 = n3253 | n2370;
  assign n2373 = ~n2371 & n2372;
  assign n3289 = n2368 | n2370;
  assign n3290 = (n2368 & n3253) | (n2368 & n3289) | (n3253 & n3289);
  assign n3291 = n2361 | n2363;
  assign n3292 = (n2361 & n3255) | (n2361 & n3291) | (n3255 & n3291);
  assign n3293 = n2354 | n2356;
  assign n3294 = (n2354 & n3257) | (n2354 & n3293) | (n3257 & n3293);
  assign n3295 = n2347 | n2349;
  assign n3296 = (n2347 & n3259) | (n2347 & n3295) | (n3259 & n3295);
  assign n3297 = n2340 | n2342;
  assign n3298 = (n2340 & n3261) | (n2340 & n3297) | (n3261 & n3297);
  assign n3299 = n2333 | n2335;
  assign n3300 = (n2333 & n3263) | (n2333 & n3299) | (n3263 & n3299);
  assign n3302 = n2319 | n2321;
  assign n3768 = n2246 | n2319;
  assign n3769 = (n2319 & n2321) | (n2319 & n3768) | (n2321 & n3768);
  assign n3770 = (n3244 & n3302) | (n3244 & n3769) | (n3302 & n3769);
  assign n3771 = (n2248 & n3302) | (n2248 & n3769) | (n3302 & n3769);
  assign n3772 = (n3212 & n3770) | (n3212 & n3771) | (n3770 & n3771);
  assign n2383 = x31 & x40;
  assign n3304 = n2383 & n3754;
  assign n3773 = (n2383 & n3304) | (n2383 & n3760) | (n3304 & n3760);
  assign n3955 = (n2314 & n2383) | (n2314 & n3304) | (n2383 & n3304);
  assign n3956 = n2383 & n3304;
  assign n3957 = (n2239 & n3955) | (n2239 & n3956) | (n3955 & n3956);
  assign n3775 = (n3732 & n3773) | (n3732 & n3957) | (n3773 & n3957);
  assign n3306 = n2383 | n3754;
  assign n3776 = n3306 | n3760;
  assign n3958 = n2314 | n3306;
  assign n3959 = (n2239 & n3306) | (n2239 & n3958) | (n3306 & n3958);
  assign n3778 = (n3732 & n3776) | (n3732 & n3959) | (n3776 & n3959);
  assign n2386 = ~n3775 & n3778;
  assign n2387 = n3772 & n2386;
  assign n2388 = n3772 | n2386;
  assign n2389 = ~n2387 & n2388;
  assign n2390 = x30 & x41;
  assign n2391 = n2389 & n2390;
  assign n2392 = n2389 | n2390;
  assign n2393 = ~n2391 & n2392;
  assign n3308 = n2326 & n2393;
  assign n3309 = (n2393 & n3286) | (n2393 & n3308) | (n3286 & n3308);
  assign n3310 = n2326 | n2393;
  assign n3311 = n3286 | n3310;
  assign n2396 = ~n3309 & n3311;
  assign n2397 = x29 & x42;
  assign n2398 = n2396 & n2397;
  assign n2399 = n2396 | n2397;
  assign n2400 = ~n2398 & n2399;
  assign n2401 = n3300 & n2400;
  assign n2402 = n3300 | n2400;
  assign n2403 = ~n2401 & n2402;
  assign n2404 = x28 & x43;
  assign n2405 = n2403 & n2404;
  assign n2406 = n2403 | n2404;
  assign n2407 = ~n2405 & n2406;
  assign n2408 = n3298 & n2407;
  assign n2409 = n3298 | n2407;
  assign n2410 = ~n2408 & n2409;
  assign n2411 = x27 & x44;
  assign n2412 = n2410 & n2411;
  assign n2413 = n2410 | n2411;
  assign n2414 = ~n2412 & n2413;
  assign n2415 = n3296 & n2414;
  assign n2416 = n3296 | n2414;
  assign n2417 = ~n2415 & n2416;
  assign n2418 = x26 & x45;
  assign n2419 = n2417 & n2418;
  assign n2420 = n2417 | n2418;
  assign n2421 = ~n2419 & n2420;
  assign n2422 = n3294 & n2421;
  assign n2423 = n3294 | n2421;
  assign n2424 = ~n2422 & n2423;
  assign n2425 = x25 & x46;
  assign n2426 = n2424 & n2425;
  assign n2427 = n2424 | n2425;
  assign n2428 = ~n2426 & n2427;
  assign n2429 = n3292 & n2428;
  assign n2430 = n3292 | n2428;
  assign n2431 = ~n2429 & n2430;
  assign n2432 = x24 & x47;
  assign n2433 = n2431 & n2432;
  assign n2434 = n2431 | n2432;
  assign n2435 = ~n2433 & n2434;
  assign n2436 = n3290 & n2435;
  assign n2437 = n3290 | n2435;
  assign n2438 = ~n2436 & n2437;
  assign n3312 = n2433 | n2435;
  assign n3313 = (n2433 & n3290) | (n2433 & n3312) | (n3290 & n3312);
  assign n3314 = n2426 | n2428;
  assign n3315 = (n2426 & n3292) | (n2426 & n3314) | (n3292 & n3314);
  assign n3316 = n2419 | n2421;
  assign n3317 = (n2419 & n3294) | (n2419 & n3316) | (n3294 & n3316);
  assign n3318 = n2412 | n2414;
  assign n3319 = (n2412 & n3296) | (n2412 & n3318) | (n3296 & n3318);
  assign n3320 = n2405 | n2407;
  assign n3321 = (n2405 & n3298) | (n2405 & n3320) | (n3298 & n3320);
  assign n3322 = n2398 | n2400;
  assign n3323 = (n2398 & n3300) | (n2398 & n3322) | (n3300 & n3322);
  assign n2447 = x31 & x41;
  assign n3962 = n2447 & n3304;
  assign n3963 = n2383 & n2447;
  assign n3964 = (n3760 & n3962) | (n3760 & n3963) | (n3962 & n3963);
  assign n3960 = n2447 & n3957;
  assign n3961 = (n3732 & n3964) | (n3732 & n3960) | (n3964 & n3960);
  assign n3780 = (n2386 & n2447) | (n2386 & n3961) | (n2447 & n3961);
  assign n3782 = n2447 & n3957;
  assign n3783 = (n3732 & n3964) | (n3732 & n3782) | (n3964 & n3782);
  assign n3328 = (n3772 & n3780) | (n3772 & n3783) | (n3780 & n3783);
  assign n3967 = n2447 | n3304;
  assign n3968 = n2383 | n2447;
  assign n3969 = (n3760 & n3967) | (n3760 & n3968) | (n3967 & n3968);
  assign n3965 = n2447 | n3957;
  assign n3966 = (n3732 & n3969) | (n3732 & n3965) | (n3969 & n3965);
  assign n3785 = n2386 | n3966;
  assign n3787 = n2447 | n3957;
  assign n3788 = (n3732 & n3969) | (n3732 & n3787) | (n3969 & n3787);
  assign n3331 = (n3772 & n3785) | (n3772 & n3788) | (n3785 & n3788);
  assign n2450 = ~n3328 & n3331;
  assign n3332 = n2391 & n2450;
  assign n3789 = (n2450 & n3308) | (n2450 & n3332) | (n3308 & n3332);
  assign n3790 = (n2393 & n2450) | (n2393 & n3332) | (n2450 & n3332);
  assign n3791 = (n3286 & n3789) | (n3286 & n3790) | (n3789 & n3790);
  assign n3334 = n2391 | n2450;
  assign n3792 = n3308 | n3334;
  assign n3793 = n2393 | n3334;
  assign n3794 = (n3286 & n3792) | (n3286 & n3793) | (n3792 & n3793);
  assign n2453 = ~n3791 & n3794;
  assign n2454 = x30 & x42;
  assign n2455 = n2453 & n2454;
  assign n2456 = n2453 | n2454;
  assign n2457 = ~n2455 & n2456;
  assign n2458 = n3323 & n2457;
  assign n2459 = n3323 | n2457;
  assign n2460 = ~n2458 & n2459;
  assign n2461 = x29 & x43;
  assign n2462 = n2460 & n2461;
  assign n2463 = n2460 | n2461;
  assign n2464 = ~n2462 & n2463;
  assign n2465 = n3321 & n2464;
  assign n2466 = n3321 | n2464;
  assign n2467 = ~n2465 & n2466;
  assign n2468 = x28 & x44;
  assign n2469 = n2467 & n2468;
  assign n2470 = n2467 | n2468;
  assign n2471 = ~n2469 & n2470;
  assign n2472 = n3319 & n2471;
  assign n2473 = n3319 | n2471;
  assign n2474 = ~n2472 & n2473;
  assign n2475 = x27 & x45;
  assign n2476 = n2474 & n2475;
  assign n2477 = n2474 | n2475;
  assign n2478 = ~n2476 & n2477;
  assign n2479 = n3317 & n2478;
  assign n2480 = n3317 | n2478;
  assign n2481 = ~n2479 & n2480;
  assign n2482 = x26 & x46;
  assign n2483 = n2481 & n2482;
  assign n2484 = n2481 | n2482;
  assign n2485 = ~n2483 & n2484;
  assign n2486 = n3315 & n2485;
  assign n2487 = n3315 | n2485;
  assign n2488 = ~n2486 & n2487;
  assign n2489 = x25 & x47;
  assign n2490 = n2488 & n2489;
  assign n2491 = n2488 | n2489;
  assign n2492 = ~n2490 & n2491;
  assign n2493 = n3313 & n2492;
  assign n2494 = n3313 | n2492;
  assign n2495 = ~n2493 & n2494;
  assign n3336 = n2490 | n2492;
  assign n3337 = (n2490 & n3313) | (n2490 & n3336) | (n3313 & n3336);
  assign n3338 = n2483 | n2485;
  assign n3339 = (n2483 & n3315) | (n2483 & n3338) | (n3315 & n3338);
  assign n3340 = n2476 | n2478;
  assign n3341 = (n2476 & n3317) | (n2476 & n3340) | (n3317 & n3340);
  assign n3342 = n2469 | n2471;
  assign n3343 = (n2469 & n3319) | (n2469 & n3342) | (n3319 & n3342);
  assign n3344 = n2462 | n2464;
  assign n3345 = (n2462 & n3321) | (n2462 & n3344) | (n3321 & n3344);
  assign n2503 = x31 & x42;
  assign n3349 = n2450 | n3328;
  assign n3795 = (n2391 & n3328) | (n2391 & n3349) | (n3328 & n3349);
  assign n3351 = n2503 & n3795;
  assign n3970 = n2503 & n3780;
  assign n3971 = n2503 & n3783;
  assign n3972 = (n3772 & n3970) | (n3772 & n3971) | (n3970 & n3971);
  assign n3797 = (n2450 & n2503) | (n2450 & n3972) | (n2503 & n3972);
  assign n3798 = (n3308 & n3351) | (n3308 & n3797) | (n3351 & n3797);
  assign n3799 = (n2393 & n3351) | (n2393 & n3797) | (n3351 & n3797);
  assign n3800 = (n3286 & n3798) | (n3286 & n3799) | (n3798 & n3799);
  assign n3354 = n2503 | n3795;
  assign n3973 = n2503 | n3780;
  assign n3974 = n2503 | n3783;
  assign n3975 = (n3772 & n3973) | (n3772 & n3974) | (n3973 & n3974);
  assign n3802 = n2450 | n3975;
  assign n3803 = (n3308 & n3354) | (n3308 & n3802) | (n3354 & n3802);
  assign n3804 = (n2393 & n3354) | (n2393 & n3802) | (n3354 & n3802);
  assign n3805 = (n3286 & n3803) | (n3286 & n3804) | (n3803 & n3804);
  assign n2506 = ~n3800 & n3805;
  assign n3807 = n2455 & n2506;
  assign n3976 = (n2457 & n2506) | (n2457 & n3807) | (n2506 & n3807);
  assign n3808 = (n3323 & n3976) | (n3323 & n3807) | (n3976 & n3807);
  assign n3810 = n2455 | n2506;
  assign n3977 = n2457 | n3810;
  assign n3811 = (n3323 & n3977) | (n3323 & n3810) | (n3977 & n3810);
  assign n2509 = ~n3808 & n3811;
  assign n2510 = x30 & x43;
  assign n2511 = n2509 & n2510;
  assign n2512 = n2509 | n2510;
  assign n2513 = ~n2511 & n2512;
  assign n2514 = n3345 & n2513;
  assign n2515 = n3345 | n2513;
  assign n2516 = ~n2514 & n2515;
  assign n2517 = x29 & x44;
  assign n2518 = n2516 & n2517;
  assign n2519 = n2516 | n2517;
  assign n2520 = ~n2518 & n2519;
  assign n2521 = n3343 & n2520;
  assign n2522 = n3343 | n2520;
  assign n2523 = ~n2521 & n2522;
  assign n2524 = x28 & x45;
  assign n2525 = n2523 & n2524;
  assign n2526 = n2523 | n2524;
  assign n2527 = ~n2525 & n2526;
  assign n2528 = n3341 & n2527;
  assign n2529 = n3341 | n2527;
  assign n2530 = ~n2528 & n2529;
  assign n2531 = x27 & x46;
  assign n2532 = n2530 & n2531;
  assign n2533 = n2530 | n2531;
  assign n2534 = ~n2532 & n2533;
  assign n2535 = n3339 & n2534;
  assign n2536 = n3339 | n2534;
  assign n2537 = ~n2535 & n2536;
  assign n2538 = x26 & x47;
  assign n2539 = n2537 & n2538;
  assign n2540 = n2537 | n2538;
  assign n2541 = ~n2539 & n2540;
  assign n2542 = n3337 & n2541;
  assign n2543 = n3337 | n2541;
  assign n2544 = ~n2542 & n2543;
  assign n3357 = n2539 | n2541;
  assign n3358 = (n2539 & n3337) | (n2539 & n3357) | (n3337 & n3357);
  assign n3359 = n2532 | n2534;
  assign n3360 = (n2532 & n3339) | (n2532 & n3359) | (n3339 & n3359);
  assign n3361 = n2525 | n2527;
  assign n3362 = (n2525 & n3341) | (n2525 & n3361) | (n3341 & n3361);
  assign n3363 = n2518 | n2520;
  assign n3364 = (n2518 & n3343) | (n2518 & n3363) | (n3343 & n3363);
  assign n2551 = x31 & x43;
  assign n3370 = n2551 & n3800;
  assign n3812 = n2551 & n3800;
  assign n3813 = (n2506 & n2551) | (n2506 & n3812) | (n2551 & n3812);
  assign n3815 = (n2455 & n3370) | (n2455 & n3813) | (n3370 & n3813);
  assign n3978 = n3370 | n3813;
  assign n3979 = (n2457 & n3815) | (n2457 & n3978) | (n3815 & n3978);
  assign n3816 = (n3323 & n3979) | (n3323 & n3815) | (n3979 & n3815);
  assign n3373 = n2551 | n3800;
  assign n3817 = n2551 | n3800;
  assign n3818 = n2506 | n3817;
  assign n3820 = (n2455 & n3373) | (n2455 & n3818) | (n3373 & n3818);
  assign n3980 = n3373 | n3818;
  assign n3981 = (n2457 & n3820) | (n2457 & n3980) | (n3820 & n3980);
  assign n3821 = (n3323 & n3981) | (n3323 & n3820) | (n3981 & n3820);
  assign n2554 = ~n3816 & n3821;
  assign n3823 = n2511 & n2554;
  assign n3982 = (n2513 & n2554) | (n2513 & n3823) | (n2554 & n3823);
  assign n3824 = (n3345 & n3982) | (n3345 & n3823) | (n3982 & n3823);
  assign n3826 = n2511 | n2554;
  assign n3983 = n2513 | n3826;
  assign n3827 = (n3345 & n3983) | (n3345 & n3826) | (n3983 & n3826);
  assign n2557 = ~n3824 & n3827;
  assign n2558 = x30 & x44;
  assign n2559 = n2557 & n2558;
  assign n2560 = n2557 | n2558;
  assign n2561 = ~n2559 & n2560;
  assign n2562 = n3364 & n2561;
  assign n2563 = n3364 | n2561;
  assign n2564 = ~n2562 & n2563;
  assign n2565 = x29 & x45;
  assign n2566 = n2564 & n2565;
  assign n2567 = n2564 | n2565;
  assign n2568 = ~n2566 & n2567;
  assign n2569 = n3362 & n2568;
  assign n2570 = n3362 | n2568;
  assign n2571 = ~n2569 & n2570;
  assign n2572 = x28 & x46;
  assign n2573 = n2571 & n2572;
  assign n2574 = n2571 | n2572;
  assign n2575 = ~n2573 & n2574;
  assign n2576 = n3360 & n2575;
  assign n2577 = n3360 | n2575;
  assign n2578 = ~n2576 & n2577;
  assign n2579 = x27 & x47;
  assign n2580 = n2578 & n2579;
  assign n2581 = n2578 | n2579;
  assign n2582 = ~n2580 & n2581;
  assign n2583 = n3358 & n2582;
  assign n2584 = n3358 | n2582;
  assign n2585 = ~n2583 & n2584;
  assign n3375 = n2580 | n2582;
  assign n3376 = (n2580 & n3358) | (n2580 & n3375) | (n3358 & n3375);
  assign n3377 = n2573 | n2575;
  assign n3378 = (n2573 & n3360) | (n2573 & n3377) | (n3360 & n3377);
  assign n3379 = n2566 | n2568;
  assign n3380 = (n2566 & n3362) | (n2566 & n3379) | (n3362 & n3379);
  assign n2591 = x31 & x44;
  assign n3984 = n2591 & n3979;
  assign n3985 = n2591 & n3815;
  assign n3986 = (n3323 & n3984) | (n3323 & n3985) | (n3984 & n3985);
  assign n3829 = (n2554 & n2591) | (n2554 & n3986) | (n2591 & n3986);
  assign n3987 = (n2511 & n3829) | (n2511 & n3986) | (n3829 & n3986);
  assign n3988 = n3829 | n3986;
  assign n3989 = (n2513 & n3987) | (n2513 & n3988) | (n3987 & n3988);
  assign n3831 = (n2511 & n3986) | (n2511 & n3829) | (n3986 & n3829);
  assign n3832 = (n3345 & n3989) | (n3345 & n3831) | (n3989 & n3831);
  assign n3990 = n2591 | n3979;
  assign n3991 = n2591 | n3815;
  assign n3992 = (n3323 & n3990) | (n3323 & n3991) | (n3990 & n3991);
  assign n3834 = n2554 | n3992;
  assign n3993 = (n2511 & n3834) | (n2511 & n3992) | (n3834 & n3992);
  assign n3994 = n3834 | n3992;
  assign n3995 = (n2513 & n3993) | (n2513 & n3994) | (n3993 & n3994);
  assign n3836 = (n2511 & n3992) | (n2511 & n3834) | (n3992 & n3834);
  assign n3837 = (n3345 & n3995) | (n3345 & n3836) | (n3995 & n3836);
  assign n2594 = ~n3832 & n3837;
  assign n3839 = n2559 & n2594;
  assign n3996 = (n2561 & n2594) | (n2561 & n3839) | (n2594 & n3839);
  assign n3840 = (n3364 & n3996) | (n3364 & n3839) | (n3996 & n3839);
  assign n3842 = n2559 | n2594;
  assign n3997 = n2561 | n3842;
  assign n3843 = (n3364 & n3997) | (n3364 & n3842) | (n3997 & n3842);
  assign n2597 = ~n3840 & n3843;
  assign n2598 = x30 & x45;
  assign n2599 = n2597 & n2598;
  assign n2600 = n2597 | n2598;
  assign n2601 = ~n2599 & n2600;
  assign n2602 = n3380 & n2601;
  assign n2603 = n3380 | n2601;
  assign n2604 = ~n2602 & n2603;
  assign n2605 = x29 & x46;
  assign n2606 = n2604 & n2605;
  assign n2607 = n2604 | n2605;
  assign n2608 = ~n2606 & n2607;
  assign n2609 = n3378 & n2608;
  assign n2610 = n3378 | n2608;
  assign n2611 = ~n2609 & n2610;
  assign n2612 = x28 & x47;
  assign n2613 = n2611 & n2612;
  assign n2614 = n2611 | n2612;
  assign n2615 = ~n2613 & n2614;
  assign n2616 = n3376 & n2615;
  assign n2617 = n3376 | n2615;
  assign n2618 = ~n2616 & n2617;
  assign n3391 = n2613 | n2615;
  assign n3392 = (n2613 & n3376) | (n2613 & n3391) | (n3376 & n3391);
  assign n3393 = n2606 | n2608;
  assign n3394 = (n2606 & n3378) | (n2606 & n3393) | (n3378 & n3393);
  assign n2623 = x31 & x45;
  assign n3998 = n2623 & n3989;
  assign n3999 = n2623 & n3831;
  assign n4000 = (n3345 & n3998) | (n3345 & n3999) | (n3998 & n3999);
  assign n3845 = (n2594 & n2623) | (n2594 & n4000) | (n2623 & n4000);
  assign n4001 = (n2559 & n3845) | (n2559 & n4000) | (n3845 & n4000);
  assign n4002 = n3845 | n4000;
  assign n4003 = (n2561 & n4001) | (n2561 & n4002) | (n4001 & n4002);
  assign n3847 = (n2559 & n4000) | (n2559 & n3845) | (n4000 & n3845);
  assign n3848 = (n3364 & n4003) | (n3364 & n3847) | (n4003 & n3847);
  assign n4004 = n2623 | n3989;
  assign n4005 = n2623 | n3831;
  assign n4006 = (n3345 & n4004) | (n3345 & n4005) | (n4004 & n4005);
  assign n3850 = n2594 | n4006;
  assign n4007 = (n2559 & n3850) | (n2559 & n4006) | (n3850 & n4006);
  assign n4008 = n3850 | n4006;
  assign n4009 = (n2561 & n4007) | (n2561 & n4008) | (n4007 & n4008);
  assign n3852 = (n2559 & n4006) | (n2559 & n3850) | (n4006 & n3850);
  assign n3853 = (n3364 & n4009) | (n3364 & n3852) | (n4009 & n3852);
  assign n2626 = ~n3848 & n3853;
  assign n3855 = n2599 & n2626;
  assign n4010 = (n2601 & n2626) | (n2601 & n3855) | (n2626 & n3855);
  assign n3856 = (n3380 & n4010) | (n3380 & n3855) | (n4010 & n3855);
  assign n3858 = n2599 | n2626;
  assign n4011 = n2601 | n3858;
  assign n3859 = (n3380 & n4011) | (n3380 & n3858) | (n4011 & n3858);
  assign n2629 = ~n3856 & n3859;
  assign n2630 = x30 & x46;
  assign n2631 = n2629 & n2630;
  assign n2632 = n2629 | n2630;
  assign n2633 = ~n2631 & n2632;
  assign n2634 = n3394 & n2633;
  assign n2635 = n3394 | n2633;
  assign n2636 = ~n2634 & n2635;
  assign n2637 = x29 & x47;
  assign n2638 = n2636 & n2637;
  assign n2639 = n2636 | n2637;
  assign n2640 = ~n2638 & n2639;
  assign n2641 = n3392 & n2640;
  assign n2642 = n3392 | n2640;
  assign n2643 = ~n2641 & n2642;
  assign n3405 = n2638 | n2640;
  assign n3406 = (n2638 & n3392) | (n2638 & n3405) | (n3392 & n3405);
  assign n2647 = x31 & x46;
  assign n4012 = n2647 & n4003;
  assign n4013 = n2647 & n3847;
  assign n4014 = (n3364 & n4012) | (n3364 & n4013) | (n4012 & n4013);
  assign n3861 = (n2626 & n2647) | (n2626 & n4014) | (n2647 & n4014);
  assign n4015 = (n2599 & n3861) | (n2599 & n4014) | (n3861 & n4014);
  assign n4016 = n3861 | n4014;
  assign n4017 = (n2601 & n4015) | (n2601 & n4016) | (n4015 & n4016);
  assign n3863 = (n2599 & n4014) | (n2599 & n3861) | (n4014 & n3861);
  assign n3864 = (n3380 & n4017) | (n3380 & n3863) | (n4017 & n3863);
  assign n4018 = n2647 | n4003;
  assign n4019 = n2647 | n3847;
  assign n4020 = (n3364 & n4018) | (n3364 & n4019) | (n4018 & n4019);
  assign n3866 = n2626 | n4020;
  assign n4021 = (n2599 & n3866) | (n2599 & n4020) | (n3866 & n4020);
  assign n4022 = n3866 | n4020;
  assign n4023 = (n2601 & n4021) | (n2601 & n4022) | (n4021 & n4022);
  assign n3868 = (n2599 & n4020) | (n2599 & n3866) | (n4020 & n3866);
  assign n3869 = (n3380 & n4023) | (n3380 & n3868) | (n4023 & n3868);
  assign n2650 = ~n3864 & n3869;
  assign n3871 = n2631 & n2650;
  assign n4024 = (n2633 & n2650) | (n2633 & n3871) | (n2650 & n3871);
  assign n3872 = (n3394 & n4024) | (n3394 & n3871) | (n4024 & n3871);
  assign n3874 = n2631 | n2650;
  assign n4025 = n2633 | n3874;
  assign n3875 = (n3394 & n4025) | (n3394 & n3874) | (n4025 & n3874);
  assign n2653 = ~n3872 & n3875;
  assign n2654 = x30 & x47;
  assign n2655 = n2653 & n2654;
  assign n2656 = n2653 | n2654;
  assign n2657 = ~n2655 & n2656;
  assign n2658 = n3406 & n2657;
  assign n2659 = n3406 | n2657;
  assign n2660 = ~n2658 & n2659;
  assign n2663 = x31 & x47;
  assign n4026 = n2663 & n4017;
  assign n4027 = n2663 & n3863;
  assign n4028 = (n3380 & n4026) | (n3380 & n4027) | (n4026 & n4027);
  assign n3877 = (n2650 & n2663) | (n2650 & n4028) | (n2663 & n4028);
  assign n4029 = (n2631 & n3877) | (n2631 & n4028) | (n3877 & n4028);
  assign n4030 = n3877 | n4028;
  assign n4031 = (n2633 & n4029) | (n2633 & n4030) | (n4029 & n4030);
  assign n3879 = (n2631 & n4028) | (n2631 & n3877) | (n4028 & n3877);
  assign n3880 = (n3394 & n4031) | (n3394 & n3879) | (n4031 & n3879);
  assign n4032 = n2663 | n4017;
  assign n4033 = n2663 | n3863;
  assign n4034 = (n3380 & n4032) | (n3380 & n4033) | (n4032 & n4033);
  assign n3882 = n2650 | n4034;
  assign n4035 = (n2631 & n3882) | (n2631 & n4034) | (n3882 & n4034);
  assign n4036 = n3882 | n4034;
  assign n4037 = (n2633 & n4035) | (n2633 & n4036) | (n4035 & n4036);
  assign n3884 = (n2631 & n4034) | (n2631 & n3882) | (n4034 & n3882);
  assign n3885 = (n3394 & n4037) | (n3394 & n3884) | (n4037 & n3884);
  assign n2666 = ~n3880 & n3885;
  assign n3887 = n2655 & n2666;
  assign n4038 = (n2657 & n2666) | (n2657 & n3887) | (n2666 & n3887);
  assign n3888 = (n3406 & n4038) | (n3406 & n3887) | (n4038 & n3887);
  assign n3890 = n2655 | n2666;
  assign n4039 = n2657 | n3890;
  assign n3891 = (n3406 & n4039) | (n3406 & n3890) | (n4039 & n3890);
  assign n2669 = ~n3888 & n3891;
  assign n3427 = n2666 | n3880;
  assign n3893 = (n2655 & n3427) | (n2655 & n3880) | (n3427 & n3880);
  assign n4040 = n3427 | n3880;
  assign n4041 = (n2657 & n3893) | (n2657 & n4040) | (n3893 & n4040);
  assign n3894 = (n3406 & n4041) | (n3406 & n3893) | (n4041 & n3893);
  assign y0 = n17;
  assign y1 = n22;
  assign y2 = n34;
  assign y3 = n54;
  assign y4 = n82;
  assign y5 = n118;
  assign y6 = n162;
  assign y7 = n214;
  assign y8 = n266;
  assign y9 = n314;
  assign y10 = n355;
  assign y11 = n388;
  assign y12 = n413;
  assign y13 = n430;
  assign y14 = n439;
  assign y15 = n723;
  assign y16 = n799;
  assign y17 = n804;
  assign y18 = n816;
  assign y19 = n836;
  assign y20 = n864;
  assign y21 = n900;
  assign y22 = n944;
  assign y23 = n996;
  assign y24 = n1056;
  assign y25 = n1124;
  assign y26 = n1200;
  assign y27 = n1284;
  assign y28 = n1376;
  assign y29 = n1476;
  assign y30 = n1584;
  assign y31 = n1700;
  assign y32 = n1816;
  assign y33 = n1928;
  assign y34 = n2033;
  assign y35 = n2130;
  assign y36 = n2219;
  assign y37 = n2300;
  assign y38 = n2373;
  assign y39 = n2438;
  assign y40 = n2495;
  assign y41 = n2544;
  assign y42 = n2585;
  assign y43 = n2618;
  assign y44 = n2643;
  assign y45 = n2660;
  assign y46 = n2669;
  assign y47 = n3894;
endmodule

