module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766;
  assign n17 = x0 & x8;
  assign n18 = x1 & x8;
  assign n19 = x0 & x9;
  assign n20 = n18 & n19;
  assign n21 = n18 | n19;
  assign n22 = ~n20 & n21;
  assign n23 = x2 & x8;
  assign n24 = x1 & x9;
  assign n25 = n23 & n24;
  assign n26 = n23 | n24;
  assign n27 = ~n25 & n26;
  assign n28 = n20 & n27;
  assign n29 = n20 | n27;
  assign n30 = ~n28 & n29;
  assign n31 = x0 & x10;
  assign n32 = n30 & n31;
  assign n33 = n30 | n31;
  assign n34 = ~n32 & n33;
  assign n441 = n20 | n25;
  assign n442 = (n25 & n27) | (n25 & n441) | (n27 & n441);
  assign n36 = x3 & x8;
  assign n37 = x2 & x9;
  assign n38 = n36 & n37;
  assign n39 = n36 | n37;
  assign n40 = ~n38 & n39;
  assign n41 = n442 & n40;
  assign n42 = n442 | n40;
  assign n43 = ~n41 & n42;
  assign n44 = x1 & x10;
  assign n45 = n43 & n44;
  assign n46 = n43 | n44;
  assign n47 = ~n45 & n46;
  assign n48 = n32 & n47;
  assign n49 = n32 | n47;
  assign n50 = ~n48 & n49;
  assign n51 = x0 & x11;
  assign n52 = n50 & n51;
  assign n53 = n50 | n51;
  assign n54 = ~n52 & n53;
  assign n443 = n32 | n45;
  assign n444 = (n45 & n47) | (n45 & n443) | (n47 & n443);
  assign n445 = n38 | n40;
  assign n446 = (n38 & n442) | (n38 & n445) | (n442 & n445);
  assign n57 = x4 & x8;
  assign n58 = x3 & x9;
  assign n59 = n57 & n58;
  assign n60 = n57 | n58;
  assign n61 = ~n59 & n60;
  assign n62 = n446 & n61;
  assign n63 = n446 | n61;
  assign n64 = ~n62 & n63;
  assign n65 = x2 & x10;
  assign n66 = n64 & n65;
  assign n67 = n64 | n65;
  assign n68 = ~n66 & n67;
  assign n69 = n444 & n68;
  assign n70 = n444 | n68;
  assign n71 = ~n69 & n70;
  assign n72 = x1 & x11;
  assign n73 = n71 & n72;
  assign n74 = n71 | n72;
  assign n75 = ~n73 & n74;
  assign n76 = n52 & n75;
  assign n77 = n52 | n75;
  assign n78 = ~n76 & n77;
  assign n79 = x0 & x12;
  assign n80 = n78 & n79;
  assign n81 = n78 | n79;
  assign n82 = ~n80 & n81;
  assign n447 = n52 | n73;
  assign n448 = (n73 & n75) | (n73 & n447) | (n75 & n447);
  assign n86 = x5 & x8;
  assign n87 = x4 & x9;
  assign n88 = n86 & n87;
  assign n89 = n86 | n87;
  assign n90 = ~n88 & n89;
  assign n449 = n59 | n61;
  assign n451 = n90 & n449;
  assign n452 = n59 & n90;
  assign n453 = (n446 & n451) | (n446 & n452) | (n451 & n452);
  assign n454 = n90 | n449;
  assign n455 = n59 | n90;
  assign n456 = (n446 & n454) | (n446 & n455) | (n454 & n455);
  assign n93 = ~n453 & n456;
  assign n94 = x3 & x10;
  assign n95 = n93 & n94;
  assign n96 = n93 | n94;
  assign n97 = ~n95 & n96;
  assign n457 = n66 & n97;
  assign n458 = (n69 & n97) | (n69 & n457) | (n97 & n457);
  assign n459 = n66 | n97;
  assign n460 = n69 | n459;
  assign n100 = ~n458 & n460;
  assign n101 = x2 & x11;
  assign n102 = n100 & n101;
  assign n103 = n100 | n101;
  assign n104 = ~n102 & n103;
  assign n105 = n448 & n104;
  assign n106 = n448 | n104;
  assign n107 = ~n105 & n106;
  assign n108 = x1 & x12;
  assign n109 = n107 & n108;
  assign n110 = n107 | n108;
  assign n111 = ~n109 & n110;
  assign n112 = n80 & n111;
  assign n113 = n80 | n111;
  assign n114 = ~n112 & n113;
  assign n115 = x0 & x13;
  assign n116 = n114 & n115;
  assign n117 = n114 | n115;
  assign n118 = ~n116 & n117;
  assign n461 = n80 | n109;
  assign n462 = (n109 & n111) | (n109 & n461) | (n111 & n461);
  assign n120 = n102 | n105;
  assign n123 = x6 & x8;
  assign n124 = x5 & x9;
  assign n125 = n123 & n124;
  assign n126 = n123 | n124;
  assign n127 = ~n125 & n126;
  assign n463 = n88 & n127;
  assign n464 = (n127 & n453) | (n127 & n463) | (n453 & n463);
  assign n465 = n88 | n127;
  assign n466 = n453 | n465;
  assign n130 = ~n464 & n466;
  assign n131 = x4 & x10;
  assign n132 = n130 & n131;
  assign n133 = n130 | n131;
  assign n134 = ~n132 & n133;
  assign n467 = n95 & n134;
  assign n468 = (n134 & n458) | (n134 & n467) | (n458 & n467);
  assign n469 = n95 | n134;
  assign n470 = n458 | n469;
  assign n137 = ~n468 & n470;
  assign n138 = x3 & x11;
  assign n139 = n137 & n138;
  assign n140 = n137 | n138;
  assign n141 = ~n139 & n140;
  assign n142 = n120 & n141;
  assign n143 = n120 | n141;
  assign n144 = ~n142 & n143;
  assign n145 = x2 & x12;
  assign n146 = n144 & n145;
  assign n147 = n144 | n145;
  assign n148 = ~n146 & n147;
  assign n149 = n462 & n148;
  assign n150 = n462 | n148;
  assign n151 = ~n149 & n150;
  assign n152 = x1 & x13;
  assign n153 = n151 & n152;
  assign n154 = n151 | n152;
  assign n155 = ~n153 & n154;
  assign n156 = n116 & n155;
  assign n157 = n116 | n155;
  assign n158 = ~n156 & n157;
  assign n159 = x0 & x14;
  assign n160 = n158 & n159;
  assign n161 = n158 | n159;
  assign n162 = ~n160 & n161;
  assign n724 = n115 | n152;
  assign n725 = (n114 & n152) | (n114 & n724) | (n152 & n724);
  assign n598 = (n116 & n151) | (n116 & n725) | (n151 & n725);
  assign n472 = (n153 & n155) | (n153 & n598) | (n155 & n598);
  assign n473 = n146 | n462;
  assign n474 = (n146 & n148) | (n146 & n473) | (n148 & n473);
  assign n475 = n139 | n141;
  assign n476 = (n120 & n139) | (n120 & n475) | (n139 & n475);
  assign n168 = x7 & x8;
  assign n169 = x6 & x9;
  assign n170 = n168 & n169;
  assign n171 = n168 | n169;
  assign n172 = ~n170 & n171;
  assign n599 = n88 | n125;
  assign n600 = (n125 & n127) | (n125 & n599) | (n127 & n599);
  assign n480 = n172 & n600;
  assign n478 = n125 | n127;
  assign n481 = n172 & n478;
  assign n482 = (n453 & n480) | (n453 & n481) | (n480 & n481);
  assign n483 = n172 | n600;
  assign n484 = n172 | n478;
  assign n485 = (n453 & n483) | (n453 & n484) | (n483 & n484);
  assign n175 = ~n482 & n485;
  assign n176 = x5 & x10;
  assign n177 = n175 & n176;
  assign n178 = n175 | n176;
  assign n179 = ~n177 & n178;
  assign n486 = n132 & n179;
  assign n487 = (n179 & n468) | (n179 & n486) | (n468 & n486);
  assign n488 = n132 | n179;
  assign n489 = n468 | n488;
  assign n182 = ~n487 & n489;
  assign n183 = x4 & x11;
  assign n184 = n182 & n183;
  assign n185 = n182 | n183;
  assign n186 = ~n184 & n185;
  assign n187 = n476 & n186;
  assign n188 = n476 | n186;
  assign n189 = ~n187 & n188;
  assign n190 = x3 & x12;
  assign n191 = n189 & n190;
  assign n192 = n189 | n190;
  assign n193 = ~n191 & n192;
  assign n194 = n474 & n193;
  assign n195 = n474 | n193;
  assign n196 = ~n194 & n195;
  assign n197 = x2 & x13;
  assign n198 = n196 & n197;
  assign n199 = n196 | n197;
  assign n200 = ~n198 & n199;
  assign n201 = n472 & n200;
  assign n202 = n472 | n200;
  assign n203 = ~n201 & n202;
  assign n204 = x1 & x14;
  assign n205 = n203 & n204;
  assign n206 = n203 | n204;
  assign n207 = ~n205 & n206;
  assign n208 = n160 & n207;
  assign n209 = n160 | n207;
  assign n210 = ~n208 & n209;
  assign n211 = x0 & x15;
  assign n212 = n210 & n211;
  assign n213 = n210 | n211;
  assign n214 = ~n212 & n213;
  assign n490 = n160 | n205;
  assign n491 = (n205 & n207) | (n205 & n490) | (n207 & n490);
  assign n216 = n198 | n201;
  assign n217 = n191 | n194;
  assign n492 = n184 | n186;
  assign n493 = (n184 & n476) | (n184 & n492) | (n476 & n492);
  assign n221 = x7 & x9;
  assign n497 = n170 & n221;
  assign n726 = (n172 & n221) | (n172 & n497) | (n221 & n497);
  assign n727 = n221 & n497;
  assign n728 = (n478 & n726) | (n478 & n727) | (n726 & n727);
  assign n729 = (n600 & n726) | (n600 & n727) | (n726 & n727);
  assign n605 = (n453 & n728) | (n453 & n729) | (n728 & n729);
  assign n499 = n170 | n221;
  assign n730 = n172 | n499;
  assign n731 = (n478 & n499) | (n478 & n730) | (n499 & n730);
  assign n732 = (n499 & n600) | (n499 & n730) | (n600 & n730);
  assign n608 = (n453 & n731) | (n453 & n732) | (n731 & n732);
  assign n224 = ~n605 & n608;
  assign n225 = x6 & x10;
  assign n226 = n224 & n225;
  assign n227 = n224 | n225;
  assign n228 = ~n226 & n227;
  assign n495 = n177 | n179;
  assign n609 = n228 & n495;
  assign n601 = n132 | n177;
  assign n602 = (n177 & n179) | (n177 & n601) | (n179 & n601);
  assign n610 = n228 & n602;
  assign n611 = (n468 & n609) | (n468 & n610) | (n609 & n610);
  assign n612 = n228 | n495;
  assign n613 = n228 | n602;
  assign n614 = (n468 & n612) | (n468 & n613) | (n612 & n613);
  assign n231 = ~n611 & n614;
  assign n232 = x5 & x11;
  assign n233 = n231 & n232;
  assign n234 = n231 | n232;
  assign n235 = ~n233 & n234;
  assign n236 = n493 & n235;
  assign n237 = n493 | n235;
  assign n238 = ~n236 & n237;
  assign n239 = x4 & x12;
  assign n240 = n238 & n239;
  assign n241 = n238 | n239;
  assign n242 = ~n240 & n241;
  assign n243 = n217 & n242;
  assign n244 = n217 | n242;
  assign n245 = ~n243 & n244;
  assign n246 = x3 & x13;
  assign n247 = n245 & n246;
  assign n248 = n245 | n246;
  assign n249 = ~n247 & n248;
  assign n250 = n216 & n249;
  assign n251 = n216 | n249;
  assign n252 = ~n250 & n251;
  assign n253 = x2 & x14;
  assign n254 = n252 & n253;
  assign n255 = n252 | n253;
  assign n256 = ~n254 & n255;
  assign n257 = n491 & n256;
  assign n258 = n491 | n256;
  assign n259 = ~n257 & n258;
  assign n260 = x1 & x15;
  assign n261 = n259 & n260;
  assign n262 = n259 | n260;
  assign n263 = ~n261 & n262;
  assign n264 = n212 & n263;
  assign n265 = n212 | n263;
  assign n266 = ~n264 & n265;
  assign n733 = n211 | n260;
  assign n734 = (n210 & n260) | (n210 & n733) | (n260 & n733);
  assign n616 = (n212 & n259) | (n212 & n734) | (n259 & n734);
  assign n502 = (n261 & n263) | (n261 & n616) | (n263 & n616);
  assign n503 = n254 | n491;
  assign n504 = (n254 & n256) | (n254 & n503) | (n256 & n503);
  assign n269 = n247 | n250;
  assign n505 = n240 | n242;
  assign n506 = (n217 & n240) | (n217 & n505) | (n240 & n505);
  assign n273 = x7 & x10;
  assign n512 = n221 & n273;
  assign n617 = n170 & n512;
  assign n735 = (n172 & n512) | (n172 & n617) | (n512 & n617);
  assign n736 = n512 & n617;
  assign n737 = (n478 & n735) | (n478 & n736) | (n735 & n736);
  assign n738 = (n600 & n735) | (n600 & n736) | (n735 & n736);
  assign n620 = (n453 & n737) | (n453 & n738) | (n737 & n738);
  assign n515 = n221 | n273;
  assign n621 = (n170 & n273) | (n170 & n515) | (n273 & n515);
  assign n739 = (n172 & n515) | (n172 & n621) | (n515 & n621);
  assign n740 = n515 & n621;
  assign n741 = (n478 & n739) | (n478 & n740) | (n739 & n740);
  assign n742 = (n600 & n739) | (n600 & n740) | (n739 & n740);
  assign n624 = (n453 & n741) | (n453 & n742) | (n741 & n742);
  assign n276 = ~n620 & n624;
  assign n518 = n226 & n276;
  assign n625 = (n228 & n276) | (n228 & n518) | (n276 & n518);
  assign n626 = (n495 & n518) | (n495 & n625) | (n518 & n625);
  assign n627 = (n518 & n602) | (n518 & n625) | (n602 & n625);
  assign n628 = (n468 & n626) | (n468 & n627) | (n626 & n627);
  assign n521 = n226 | n276;
  assign n629 = n228 | n521;
  assign n630 = (n495 & n521) | (n495 & n629) | (n521 & n629);
  assign n631 = (n521 & n602) | (n521 & n629) | (n602 & n629);
  assign n632 = (n468 & n630) | (n468 & n631) | (n630 & n631);
  assign n279 = ~n628 & n632;
  assign n280 = x6 & x11;
  assign n281 = n279 & n280;
  assign n282 = n279 | n280;
  assign n283 = ~n281 & n282;
  assign n507 = n233 | n235;
  assign n633 = n283 & n507;
  assign n634 = n233 & n283;
  assign n635 = (n493 & n633) | (n493 & n634) | (n633 & n634);
  assign n636 = n283 | n507;
  assign n637 = n233 | n283;
  assign n638 = (n493 & n636) | (n493 & n637) | (n636 & n637);
  assign n286 = ~n635 & n638;
  assign n287 = x5 & x12;
  assign n288 = n286 & n287;
  assign n289 = n286 | n287;
  assign n290 = ~n288 & n289;
  assign n291 = n506 & n290;
  assign n292 = n506 | n290;
  assign n293 = ~n291 & n292;
  assign n294 = x4 & x13;
  assign n295 = n293 & n294;
  assign n296 = n293 | n294;
  assign n297 = ~n295 & n296;
  assign n298 = n269 & n297;
  assign n299 = n269 | n297;
  assign n300 = ~n298 & n299;
  assign n301 = x3 & x14;
  assign n302 = n300 & n301;
  assign n303 = n300 | n301;
  assign n304 = ~n302 & n303;
  assign n305 = n504 & n304;
  assign n306 = n504 | n304;
  assign n307 = ~n305 & n306;
  assign n308 = x2 & x15;
  assign n309 = n307 & n308;
  assign n310 = n307 | n308;
  assign n311 = ~n309 & n310;
  assign n312 = n502 & n311;
  assign n313 = n502 | n311;
  assign n314 = ~n312 & n313;
  assign n523 = n309 | n502;
  assign n524 = (n309 & n311) | (n309 & n523) | (n311 & n523);
  assign n525 = n302 | n504;
  assign n526 = (n302 & n304) | (n302 & n525) | (n304 & n525);
  assign n527 = n295 | n297;
  assign n528 = (n269 & n295) | (n269 & n527) | (n295 & n527);
  assign n321 = x7 & x11;
  assign n743 = n321 & n738;
  assign n744 = n321 & n737;
  assign n745 = (n453 & n743) | (n453 & n744) | (n743 & n744);
  assign n534 = (n321 & n628) | (n321 & n745) | (n628 & n745);
  assign n746 = n321 | n738;
  assign n747 = n321 | n737;
  assign n748 = (n453 & n746) | (n453 & n747) | (n746 & n747);
  assign n536 = n628 | n748;
  assign n324 = ~n534 & n536;
  assign n538 = n281 & n324;
  assign n639 = (n283 & n324) | (n283 & n538) | (n324 & n538);
  assign n640 = (n507 & n538) | (n507 & n639) | (n538 & n639);
  assign n641 = (n233 & n538) | (n233 & n639) | (n538 & n639);
  assign n642 = (n493 & n640) | (n493 & n641) | (n640 & n641);
  assign n541 = n281 | n324;
  assign n643 = n283 | n541;
  assign n644 = (n507 & n541) | (n507 & n643) | (n541 & n643);
  assign n645 = (n233 & n541) | (n233 & n643) | (n541 & n643);
  assign n646 = (n493 & n644) | (n493 & n645) | (n644 & n645);
  assign n327 = ~n642 & n646;
  assign n328 = x6 & x12;
  assign n329 = n327 & n328;
  assign n330 = n327 | n328;
  assign n331 = ~n329 & n330;
  assign n529 = n288 | n290;
  assign n647 = n331 & n529;
  assign n648 = n288 & n331;
  assign n649 = (n506 & n647) | (n506 & n648) | (n647 & n648);
  assign n650 = n331 | n529;
  assign n651 = n288 | n331;
  assign n652 = (n506 & n650) | (n506 & n651) | (n650 & n651);
  assign n334 = ~n649 & n652;
  assign n335 = x5 & x13;
  assign n336 = n334 & n335;
  assign n337 = n334 | n335;
  assign n338 = ~n336 & n337;
  assign n339 = n528 & n338;
  assign n340 = n528 | n338;
  assign n341 = ~n339 & n340;
  assign n342 = x4 & x14;
  assign n343 = n341 & n342;
  assign n344 = n341 | n342;
  assign n345 = ~n343 & n344;
  assign n346 = n526 & n345;
  assign n347 = n526 | n345;
  assign n348 = ~n346 & n347;
  assign n349 = x3 & x15;
  assign n350 = n348 & n349;
  assign n351 = n348 | n349;
  assign n352 = ~n350 & n351;
  assign n353 = n524 & n352;
  assign n354 = n524 | n352;
  assign n355 = ~n353 & n354;
  assign n356 = n350 | n353;
  assign n361 = x7 & x12;
  assign n653 = n361 & n745;
  assign n654 = n321 & n361;
  assign n655 = (n628 & n653) | (n628 & n654) | (n653 & n654);
  assign n548 = (n361 & n642) | (n361 & n655) | (n642 & n655);
  assign n656 = n361 | n745;
  assign n657 = n321 | n361;
  assign n658 = (n628 & n656) | (n628 & n657) | (n656 & n657);
  assign n550 = n642 | n658;
  assign n364 = ~n548 & n550;
  assign n552 = n329 & n364;
  assign n659 = (n331 & n364) | (n331 & n552) | (n364 & n552);
  assign n660 = (n529 & n552) | (n529 & n659) | (n552 & n659);
  assign n661 = (n288 & n552) | (n288 & n659) | (n552 & n659);
  assign n662 = (n506 & n660) | (n506 & n661) | (n660 & n661);
  assign n555 = n329 | n364;
  assign n663 = n331 | n555;
  assign n664 = (n529 & n555) | (n529 & n663) | (n555 & n663);
  assign n665 = (n288 & n555) | (n288 & n663) | (n555 & n663);
  assign n666 = (n506 & n664) | (n506 & n665) | (n664 & n665);
  assign n367 = ~n662 & n666;
  assign n368 = x6 & x13;
  assign n369 = n367 & n368;
  assign n370 = n367 | n368;
  assign n371 = ~n369 & n370;
  assign n543 = n336 | n338;
  assign n667 = n371 & n543;
  assign n668 = n336 & n371;
  assign n669 = (n528 & n667) | (n528 & n668) | (n667 & n668);
  assign n670 = n371 | n543;
  assign n671 = n336 | n371;
  assign n672 = (n528 & n670) | (n528 & n671) | (n670 & n671);
  assign n374 = ~n669 & n672;
  assign n375 = x5 & x14;
  assign n376 = n374 & n375;
  assign n377 = n374 | n375;
  assign n378 = ~n376 & n377;
  assign n673 = n343 & n378;
  assign n674 = (n346 & n378) | (n346 & n673) | (n378 & n673);
  assign n675 = n343 | n378;
  assign n676 = n346 | n675;
  assign n381 = ~n674 & n676;
  assign n382 = x4 & x15;
  assign n383 = n381 & n382;
  assign n384 = n381 | n382;
  assign n385 = ~n383 & n384;
  assign n386 = n356 & n385;
  assign n387 = n356 | n385;
  assign n388 = ~n386 & n387;
  assign n677 = n383 | n385;
  assign n678 = (n356 & n383) | (n356 & n677) | (n383 & n677);
  assign n357 = n343 | n346;
  assign n393 = x7 & x13;
  assign n749 = n393 & n653;
  assign n750 = n393 & n654;
  assign n751 = (n628 & n749) | (n628 & n750) | (n749 & n750);
  assign n680 = n361 & n393;
  assign n681 = (n642 & n751) | (n642 & n680) | (n751 & n680);
  assign n562 = (n393 & n662) | (n393 & n681) | (n662 & n681);
  assign n752 = n393 | n653;
  assign n753 = n393 | n654;
  assign n754 = (n628 & n752) | (n628 & n753) | (n752 & n753);
  assign n683 = n361 | n393;
  assign n684 = (n642 & n754) | (n642 & n683) | (n754 & n683);
  assign n564 = n662 | n684;
  assign n396 = ~n562 & n564;
  assign n566 = n369 & n396;
  assign n685 = (n371 & n396) | (n371 & n566) | (n396 & n566);
  assign n686 = (n543 & n566) | (n543 & n685) | (n566 & n685);
  assign n687 = (n336 & n566) | (n336 & n685) | (n566 & n685);
  assign n688 = (n528 & n686) | (n528 & n687) | (n686 & n687);
  assign n569 = n369 | n396;
  assign n689 = n371 | n569;
  assign n690 = (n543 & n569) | (n543 & n689) | (n569 & n689);
  assign n691 = (n336 & n569) | (n336 & n689) | (n569 & n689);
  assign n692 = (n528 & n690) | (n528 & n691) | (n690 & n691);
  assign n399 = ~n688 & n692;
  assign n400 = x6 & x14;
  assign n401 = n399 & n400;
  assign n402 = n399 | n400;
  assign n403 = ~n401 & n402;
  assign n557 = n376 | n378;
  assign n693 = n403 & n557;
  assign n694 = n376 & n403;
  assign n695 = (n357 & n693) | (n357 & n694) | (n693 & n694);
  assign n696 = n403 | n557;
  assign n697 = n376 | n403;
  assign n698 = (n357 & n696) | (n357 & n697) | (n696 & n697);
  assign n406 = ~n695 & n698;
  assign n407 = x5 & x15;
  assign n408 = n406 & n407;
  assign n409 = n406 | n407;
  assign n410 = ~n408 & n409;
  assign n411 = n678 & n410;
  assign n412 = n678 | n410;
  assign n413 = ~n411 & n412;
  assign n571 = n408 | n410;
  assign n572 = (n678 & n408) | (n678 & n571) | (n408 & n571);
  assign n417 = x7 & x14;
  assign n755 = n417 & n751;
  assign n756 = n417 & n680;
  assign n757 = (n642 & n755) | (n642 & n756) | (n755 & n756);
  assign n700 = n393 & n417;
  assign n701 = (n662 & n757) | (n662 & n700) | (n757 & n700);
  assign n576 = (n417 & n688) | (n417 & n701) | (n688 & n701);
  assign n758 = n417 | n751;
  assign n759 = n417 | n680;
  assign n760 = (n642 & n758) | (n642 & n759) | (n758 & n759);
  assign n703 = n393 | n417;
  assign n704 = (n662 & n760) | (n662 & n703) | (n760 & n703);
  assign n578 = n688 | n704;
  assign n420 = ~n576 & n578;
  assign n580 = n401 & n420;
  assign n705 = (n403 & n420) | (n403 & n580) | (n420 & n580);
  assign n706 = (n557 & n580) | (n557 & n705) | (n580 & n705);
  assign n707 = (n376 & n580) | (n376 & n705) | (n580 & n705);
  assign n708 = (n357 & n706) | (n357 & n707) | (n706 & n707);
  assign n583 = n401 | n420;
  assign n709 = n403 | n583;
  assign n710 = (n557 & n583) | (n557 & n709) | (n583 & n709);
  assign n711 = (n376 & n583) | (n376 & n709) | (n583 & n709);
  assign n712 = (n357 & n710) | (n357 & n711) | (n710 & n711);
  assign n423 = ~n708 & n712;
  assign n424 = x6 & x15;
  assign n425 = n423 & n424;
  assign n426 = n423 | n424;
  assign n427 = ~n425 & n426;
  assign n428 = n572 & n427;
  assign n429 = n572 | n427;
  assign n430 = ~n428 & n429;
  assign n433 = x7 & x15;
  assign n761 = n433 & n757;
  assign n762 = n433 & n700;
  assign n763 = (n662 & n761) | (n662 & n762) | (n761 & n762);
  assign n714 = n417 & n433;
  assign n715 = (n688 & n763) | (n688 & n714) | (n763 & n714);
  assign n588 = (n433 & n708) | (n433 & n715) | (n708 & n715);
  assign n764 = n433 | n757;
  assign n765 = n433 | n700;
  assign n766 = (n662 & n764) | (n662 & n765) | (n764 & n765);
  assign n717 = n417 | n433;
  assign n718 = (n688 & n766) | (n688 & n717) | (n766 & n717);
  assign n590 = n708 | n718;
  assign n436 = ~n588 & n590;
  assign n592 = n425 & n436;
  assign n719 = (n427 & n436) | (n427 & n592) | (n436 & n592);
  assign n593 = (n572 & n719) | (n572 & n592) | (n719 & n592);
  assign n595 = n425 | n436;
  assign n720 = n427 | n595;
  assign n596 = (n572 & n720) | (n572 & n595) | (n720 & n595);
  assign n439 = ~n593 & n596;
  assign n721 = n588 | n719;
  assign n722 = n588 | n592;
  assign n723 = (n572 & n721) | (n572 & n722) | (n721 & n722);
  assign y0 = n17;
  assign y1 = n22;
  assign y2 = n34;
  assign y3 = n54;
  assign y4 = n82;
  assign y5 = n118;
  assign y6 = n162;
  assign y7 = n214;
  assign y8 = n266;
  assign y9 = n314;
  assign y10 = n355;
  assign y11 = n388;
  assign y12 = n413;
  assign y13 = n430;
  assign y14 = n439;
  assign y15 = n723;
endmodule

