module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085;
  assign n17 = x0 & x8;
  assign n18 = x0 | x8;
  assign n19 = ~n17 & n18;
  assign n20 = x1 & x9;
  assign n21 = x1 | x9;
  assign n22 = ~n20 & n21;
  assign n23 = n17 & n22;
  assign n24 = n17 | n22;
  assign n25 = ~n23 & n24;
  assign n69 = n17 | n20;
  assign n70 = (n20 & n22) | (n20 & n69) | (n22 & n69);
  assign n27 = x2 & x10;
  assign n28 = x2 | x10;
  assign n29 = ~n27 & n28;
  assign n30 = n70 & n29;
  assign n31 = n70 | n29;
  assign n32 = ~n30 & n31;
  assign n71 = n27 | n29;
  assign n72 = (n27 & n70) | (n27 & n71) | (n70 & n71);
  assign n34 = x3 & x11;
  assign n35 = x3 | x11;
  assign n36 = ~n34 & n35;
  assign n37 = n72 & n36;
  assign n38 = n72 | n36;
  assign n39 = ~n37 & n38;
  assign n41 = x4 & x12;
  assign n42 = x4 | x12;
  assign n43 = ~n41 & n42;
  assign n73 = n34 | n36;
  assign n75 = n43 & n73;
  assign n76 = n34 & n43;
  assign n77 = (n72 & n75) | (n72 & n76) | (n75 & n76);
  assign n78 = n43 | n73;
  assign n79 = n34 | n43;
  assign n80 = (n72 & n78) | (n72 & n79) | (n78 & n79);
  assign n46 = ~n77 & n80;
  assign n48 = x5 & x13;
  assign n49 = x5 | x13;
  assign n50 = ~n48 & n49;
  assign n81 = n41 & n50;
  assign n82 = (n50 & n77) | (n50 & n81) | (n77 & n81);
  assign n83 = n41 | n50;
  assign n84 = n77 | n83;
  assign n53 = ~n82 & n84;
  assign n55 = x6 & x14;
  assign n56 = x6 | x14;
  assign n57 = ~n55 & n56;
  assign n101 = n41 | n48;
  assign n102 = (n48 & n50) | (n48 & n101) | (n50 & n101);
  assign n88 = n57 & n102;
  assign n86 = n48 | n50;
  assign n89 = n57 & n86;
  assign n90 = (n77 & n88) | (n77 & n89) | (n88 & n89);
  assign n91 = n57 | n102;
  assign n92 = n57 | n86;
  assign n93 = (n77 & n91) | (n77 & n92) | (n91 & n92);
  assign n60 = ~n90 & n93;
  assign n62 = x7 & x15;
  assign n63 = x7 | x15;
  assign n64 = ~n62 & n63;
  assign n94 = n55 & n64;
  assign n103 = (n64 & n89) | (n64 & n94) | (n89 & n94);
  assign n104 = (n64 & n88) | (n64 & n94) | (n88 & n94);
  assign n105 = (n77 & n103) | (n77 & n104) | (n103 & n104);
  assign n96 = n55 | n64;
  assign n106 = n89 | n96;
  assign n107 = n88 | n96;
  assign n108 = (n77 & n106) | (n77 & n107) | (n106 & n107);
  assign n67 = ~n105 & n108;
  assign n99 = n62 | n64;
  assign n109 = n55 | n62;
  assign n110 = (n62 & n64) | (n62 & n109) | (n64 & n109);
  assign n111 = (n89 & n99) | (n89 & n110) | (n99 & n110);
  assign n112 = (n88 & n99) | (n88 & n110) | (n99 & n110);
  assign n113 = (n77 & n111) | (n77 & n112) | (n111 & n112);
  assign n146 = x16 & x32;
  assign n147 = x16 | x32;
  assign n148 = ~n146 & n147;
  assign n149 = x17 & x33;
  assign n150 = x17 | x33;
  assign n151 = ~n149 & n150;
  assign n152 = n146 & n151;
  assign n153 = n146 | n151;
  assign n154 = ~n152 & n153;
  assign n254 = n146 | n149;
  assign n255 = (n149 & n151) | (n149 & n254) | (n151 & n254);
  assign n156 = x18 & x34;
  assign n157 = x18 | x34;
  assign n158 = ~n156 & n157;
  assign n159 = n255 & n158;
  assign n160 = n255 | n158;
  assign n161 = ~n159 & n160;
  assign n256 = n156 | n158;
  assign n257 = (n156 & n255) | (n156 & n256) | (n255 & n256);
  assign n163 = x19 & x35;
  assign n164 = x19 | x35;
  assign n165 = ~n163 & n164;
  assign n166 = n257 & n165;
  assign n167 = n257 | n165;
  assign n168 = ~n166 & n167;
  assign n170 = x20 & x36;
  assign n171 = x20 | x36;
  assign n172 = ~n170 & n171;
  assign n258 = n163 | n165;
  assign n260 = n172 & n258;
  assign n261 = n163 & n172;
  assign n262 = (n257 & n260) | (n257 & n261) | (n260 & n261);
  assign n263 = n172 | n258;
  assign n264 = n163 | n172;
  assign n265 = (n257 & n263) | (n257 & n264) | (n263 & n264);
  assign n175 = ~n262 & n265;
  assign n177 = x21 & x37;
  assign n178 = x21 | x37;
  assign n179 = ~n177 & n178;
  assign n266 = n170 & n179;
  assign n267 = (n179 & n262) | (n179 & n266) | (n262 & n266);
  assign n268 = n170 | n179;
  assign n269 = n262 | n268;
  assign n182 = ~n267 & n269;
  assign n184 = x22 & x38;
  assign n185 = x22 | x38;
  assign n186 = ~n184 & n185;
  assign n341 = n170 | n177;
  assign n342 = (n177 & n179) | (n177 & n341) | (n179 & n341);
  assign n273 = n186 & n342;
  assign n271 = n177 | n179;
  assign n274 = n186 & n271;
  assign n275 = (n262 & n273) | (n262 & n274) | (n273 & n274);
  assign n276 = n186 | n342;
  assign n277 = n186 | n271;
  assign n278 = (n262 & n276) | (n262 & n277) | (n276 & n277);
  assign n189 = ~n275 & n278;
  assign n191 = x23 & x39;
  assign n192 = x23 | x39;
  assign n193 = ~n191 & n192;
  assign n279 = n184 & n193;
  assign n343 = (n193 & n274) | (n193 & n279) | (n274 & n279);
  assign n344 = (n193 & n273) | (n193 & n279) | (n273 & n279);
  assign n345 = (n262 & n343) | (n262 & n344) | (n343 & n344);
  assign n281 = n184 | n193;
  assign n346 = n274 | n281;
  assign n347 = n273 | n281;
  assign n348 = (n262 & n346) | (n262 & n347) | (n346 & n347);
  assign n196 = ~n345 & n348;
  assign n198 = x24 & x40;
  assign n199 = x24 | x40;
  assign n200 = ~n198 & n199;
  assign n349 = n184 | n191;
  assign n350 = (n191 & n193) | (n191 & n349) | (n193 & n349);
  assign n286 = n200 & n350;
  assign n284 = n191 | n193;
  assign n287 = n200 & n284;
  assign n351 = (n274 & n286) | (n274 & n287) | (n286 & n287);
  assign n352 = (n273 & n286) | (n273 & n287) | (n286 & n287);
  assign n353 = (n262 & n351) | (n262 & n352) | (n351 & n352);
  assign n289 = n200 | n350;
  assign n290 = n200 | n284;
  assign n354 = (n274 & n289) | (n274 & n290) | (n289 & n290);
  assign n355 = (n273 & n289) | (n273 & n290) | (n289 & n290);
  assign n356 = (n262 & n354) | (n262 & n355) | (n354 & n355);
  assign n203 = ~n353 & n356;
  assign n357 = n198 | n200;
  assign n358 = (n198 & n350) | (n198 & n357) | (n350 & n357);
  assign n359 = (n198 & n284) | (n198 & n357) | (n284 & n357);
  assign n360 = (n274 & n358) | (n274 & n359) | (n358 & n359);
  assign n361 = (n273 & n358) | (n273 & n359) | (n358 & n359);
  assign n362 = (n262 & n360) | (n262 & n361) | (n360 & n361);
  assign n205 = x25 & x41;
  assign n206 = x25 | x41;
  assign n207 = ~n205 & n206;
  assign n208 = n362 & n207;
  assign n209 = n362 | n207;
  assign n210 = ~n208 & n209;
  assign n212 = x26 & x42;
  assign n213 = x26 | x42;
  assign n214 = ~n212 & n213;
  assign n295 = n205 | n207;
  assign n297 = n214 & n295;
  assign n298 = n205 & n214;
  assign n299 = (n362 & n297) | (n362 & n298) | (n297 & n298);
  assign n300 = n214 | n295;
  assign n301 = n205 | n214;
  assign n302 = (n362 & n300) | (n362 & n301) | (n300 & n301);
  assign n217 = ~n299 & n302;
  assign n219 = x27 & x43;
  assign n220 = x27 | x43;
  assign n221 = ~n219 & n220;
  assign n363 = n212 | n214;
  assign n364 = (n212 & n295) | (n212 & n363) | (n295 & n363);
  assign n306 = n221 & n364;
  assign n365 = n205 | n212;
  assign n366 = (n212 & n214) | (n212 & n365) | (n214 & n365);
  assign n307 = n221 & n366;
  assign n308 = (n362 & n306) | (n362 & n307) | (n306 & n307);
  assign n309 = n221 | n364;
  assign n310 = n221 | n366;
  assign n311 = (n362 & n309) | (n362 & n310) | (n309 & n310);
  assign n224 = ~n308 & n311;
  assign n226 = x28 & x44;
  assign n227 = x28 | x44;
  assign n228 = ~n226 & n227;
  assign n367 = n219 | n221;
  assign n691 = n228 & n367;
  assign n692 = n219 & n228;
  assign n693 = (n364 & n691) | (n364 & n692) | (n691 & n692);
  assign n369 = (n219 & n366) | (n219 & n367) | (n366 & n367);
  assign n371 = n228 & n369;
  assign n372 = (n362 & n693) | (n362 & n371) | (n693 & n371);
  assign n694 = n228 | n367;
  assign n695 = n219 | n228;
  assign n696 = (n364 & n694) | (n364 & n695) | (n694 & n695);
  assign n374 = n228 | n369;
  assign n375 = (n362 & n696) | (n362 & n374) | (n696 & n374);
  assign n231 = ~n372 & n375;
  assign n233 = x29 & x45;
  assign n234 = x29 | x45;
  assign n235 = ~n233 & n234;
  assign n315 = n226 | n228;
  assign n317 = n235 & n315;
  assign n318 = n226 & n235;
  assign n368 = (n219 & n364) | (n219 & n367) | (n364 & n367);
  assign n376 = (n317 & n318) | (n317 & n368) | (n318 & n368);
  assign n377 = (n317 & n318) | (n317 & n369) | (n318 & n369);
  assign n378 = (n362 & n376) | (n362 & n377) | (n376 & n377);
  assign n320 = n235 | n315;
  assign n321 = n226 | n235;
  assign n379 = (n320 & n321) | (n320 & n368) | (n321 & n368);
  assign n380 = (n320 & n321) | (n320 & n369) | (n321 & n369);
  assign n381 = (n362 & n379) | (n362 & n380) | (n379 & n380);
  assign n238 = ~n378 & n381;
  assign n240 = x30 & x46;
  assign n241 = x30 | x46;
  assign n242 = ~n240 & n241;
  assign n382 = n233 | n235;
  assign n383 = (n233 & n315) | (n233 & n382) | (n315 & n382);
  assign n326 = n242 & n383;
  assign n384 = n226 | n233;
  assign n385 = (n233 & n235) | (n233 & n384) | (n235 & n384);
  assign n327 = n242 & n385;
  assign n386 = (n326 & n327) | (n326 & n368) | (n327 & n368);
  assign n387 = (n326 & n327) | (n326 & n369) | (n327 & n369);
  assign n388 = (n362 & n386) | (n362 & n387) | (n386 & n387);
  assign n329 = n242 | n383;
  assign n330 = n242 | n385;
  assign n389 = (n329 & n330) | (n329 & n368) | (n330 & n368);
  assign n390 = (n329 & n330) | (n329 & n369) | (n330 & n369);
  assign n391 = (n362 & n389) | (n362 & n390) | (n389 & n390);
  assign n245 = ~n388 & n391;
  assign n247 = x31 & x47;
  assign n248 = x31 | x47;
  assign n249 = ~n247 & n248;
  assign n392 = n240 | n242;
  assign n397 = (n240 & n385) | (n240 & n392) | (n385 & n392);
  assign n336 = n249 & n397;
  assign n394 = n249 & n392;
  assign n395 = n240 & n249;
  assign n396 = (n383 & n394) | (n383 & n395) | (n394 & n395);
  assign n398 = (n336 & n368) | (n336 & n396) | (n368 & n396);
  assign n399 = (n336 & n369) | (n336 & n396) | (n369 & n396);
  assign n400 = (n362 & n398) | (n362 & n399) | (n398 & n399);
  assign n339 = n249 | n397;
  assign n401 = n249 | n392;
  assign n402 = n240 | n249;
  assign n403 = (n383 & n401) | (n383 & n402) | (n401 & n402);
  assign n404 = (n339 & n368) | (n339 & n403) | (n368 & n403);
  assign n405 = (n339 & n369) | (n339 & n403) | (n369 & n403);
  assign n406 = (n362 & n404) | (n362 & n405) | (n404 & n405);
  assign n252 = ~n400 & n406;
  assign n253 = n247 | n400;
  assign n471 = x48 & x80;
  assign n472 = x48 | x80;
  assign n473 = ~n471 & n472;
  assign n474 = x49 & x81;
  assign n475 = x49 | x81;
  assign n476 = ~n474 & n475;
  assign n477 = n471 & n476;
  assign n478 = n471 | n476;
  assign n479 = ~n477 & n478;
  assign n697 = n471 | n474;
  assign n698 = (n474 & n476) | (n474 & n697) | (n476 & n697);
  assign n481 = x50 & x82;
  assign n482 = x50 | x82;
  assign n483 = ~n481 & n482;
  assign n484 = n698 & n483;
  assign n485 = n698 | n483;
  assign n486 = ~n484 & n485;
  assign n699 = n481 | n483;
  assign n700 = (n481 & n698) | (n481 & n699) | (n698 & n699);
  assign n488 = x51 & x83;
  assign n489 = x51 | x83;
  assign n490 = ~n488 & n489;
  assign n491 = n700 & n490;
  assign n492 = n700 | n490;
  assign n493 = ~n491 & n492;
  assign n495 = x52 & x84;
  assign n496 = x52 | x84;
  assign n497 = ~n495 & n496;
  assign n701 = n488 | n490;
  assign n703 = n497 & n701;
  assign n704 = n488 & n497;
  assign n705 = (n700 & n703) | (n700 & n704) | (n703 & n704);
  assign n706 = n497 | n701;
  assign n707 = n488 | n497;
  assign n708 = (n700 & n706) | (n700 & n707) | (n706 & n707);
  assign n500 = ~n705 & n708;
  assign n502 = x53 & x85;
  assign n503 = x53 | x85;
  assign n504 = ~n502 & n503;
  assign n709 = n495 & n504;
  assign n710 = (n504 & n705) | (n504 & n709) | (n705 & n709);
  assign n711 = n495 | n504;
  assign n712 = n705 | n711;
  assign n507 = ~n710 & n712;
  assign n509 = x54 & x86;
  assign n510 = x54 | x86;
  assign n511 = ~n509 & n510;
  assign n907 = n495 | n502;
  assign n908 = (n502 & n504) | (n502 & n907) | (n504 & n907);
  assign n716 = n511 & n908;
  assign n714 = n502 | n504;
  assign n717 = n511 & n714;
  assign n718 = (n705 & n716) | (n705 & n717) | (n716 & n717);
  assign n719 = n511 | n908;
  assign n720 = n511 | n714;
  assign n721 = (n705 & n719) | (n705 & n720) | (n719 & n720);
  assign n514 = ~n718 & n721;
  assign n516 = x55 & x87;
  assign n517 = x55 | x87;
  assign n518 = ~n516 & n517;
  assign n722 = n509 & n518;
  assign n909 = (n518 & n717) | (n518 & n722) | (n717 & n722);
  assign n910 = (n518 & n716) | (n518 & n722) | (n716 & n722);
  assign n911 = (n705 & n909) | (n705 & n910) | (n909 & n910);
  assign n724 = n509 | n518;
  assign n912 = n717 | n724;
  assign n913 = n716 | n724;
  assign n914 = (n705 & n912) | (n705 & n913) | (n912 & n913);
  assign n521 = ~n911 & n914;
  assign n523 = x56 & x88;
  assign n524 = x56 | x88;
  assign n525 = ~n523 & n524;
  assign n915 = n509 | n516;
  assign n916 = (n516 & n518) | (n516 & n915) | (n518 & n915);
  assign n729 = n525 & n916;
  assign n727 = n516 | n518;
  assign n730 = n525 & n727;
  assign n917 = (n717 & n729) | (n717 & n730) | (n729 & n730);
  assign n918 = (n716 & n729) | (n716 & n730) | (n729 & n730);
  assign n919 = (n705 & n917) | (n705 & n918) | (n917 & n918);
  assign n732 = n525 | n916;
  assign n733 = n525 | n727;
  assign n920 = (n717 & n732) | (n717 & n733) | (n732 & n733);
  assign n921 = (n716 & n732) | (n716 & n733) | (n732 & n733);
  assign n922 = (n705 & n920) | (n705 & n921) | (n920 & n921);
  assign n528 = ~n919 & n922;
  assign n923 = n523 | n525;
  assign n924 = (n523 & n916) | (n523 & n923) | (n916 & n923);
  assign n925 = (n523 & n727) | (n523 & n923) | (n727 & n923);
  assign n926 = (n717 & n924) | (n717 & n925) | (n924 & n925);
  assign n927 = (n716 & n924) | (n716 & n925) | (n924 & n925);
  assign n928 = (n705 & n926) | (n705 & n927) | (n926 & n927);
  assign n530 = x57 & x89;
  assign n531 = x57 | x89;
  assign n532 = ~n530 & n531;
  assign n533 = n928 & n532;
  assign n534 = n928 | n532;
  assign n535 = ~n533 & n534;
  assign n537 = x58 & x90;
  assign n538 = x58 | x90;
  assign n539 = ~n537 & n538;
  assign n738 = n530 | n532;
  assign n740 = n539 & n738;
  assign n741 = n530 & n539;
  assign n742 = (n928 & n740) | (n928 & n741) | (n740 & n741);
  assign n743 = n539 | n738;
  assign n744 = n530 | n539;
  assign n745 = (n928 & n743) | (n928 & n744) | (n743 & n744);
  assign n542 = ~n742 & n745;
  assign n544 = x59 & x91;
  assign n545 = x59 | x91;
  assign n546 = ~n544 & n545;
  assign n929 = n537 | n539;
  assign n930 = (n537 & n738) | (n537 & n929) | (n738 & n929);
  assign n749 = n546 & n930;
  assign n931 = n530 | n537;
  assign n932 = (n537 & n539) | (n537 & n931) | (n539 & n931);
  assign n750 = n546 & n932;
  assign n751 = (n928 & n749) | (n928 & n750) | (n749 & n750);
  assign n752 = n546 | n930;
  assign n753 = n546 | n932;
  assign n754 = (n928 & n752) | (n928 & n753) | (n752 & n753);
  assign n549 = ~n751 & n754;
  assign n551 = x60 & x92;
  assign n552 = x60 | x92;
  assign n553 = ~n551 & n552;
  assign n933 = n544 | n546;
  assign n934 = (n544 & n930) | (n544 & n933) | (n930 & n933);
  assign n936 = n553 & n934;
  assign n935 = (n544 & n932) | (n544 & n933) | (n932 & n933);
  assign n937 = n553 & n935;
  assign n938 = (n928 & n936) | (n928 & n937) | (n936 & n937);
  assign n939 = n553 | n934;
  assign n940 = n553 | n935;
  assign n941 = (n928 & n939) | (n928 & n940) | (n939 & n940);
  assign n556 = ~n938 & n941;
  assign n558 = x61 & x93;
  assign n559 = x61 | x93;
  assign n560 = ~n558 & n559;
  assign n758 = n551 | n553;
  assign n760 = n560 & n758;
  assign n761 = n551 & n560;
  assign n942 = (n760 & n761) | (n760 & n934) | (n761 & n934);
  assign n943 = (n760 & n761) | (n760 & n935) | (n761 & n935);
  assign n944 = (n928 & n942) | (n928 & n943) | (n942 & n943);
  assign n763 = n560 | n758;
  assign n764 = n551 | n560;
  assign n945 = (n763 & n764) | (n763 & n934) | (n764 & n934);
  assign n946 = (n763 & n764) | (n763 & n935) | (n764 & n935);
  assign n947 = (n928 & n945) | (n928 & n946) | (n945 & n946);
  assign n563 = ~n944 & n947;
  assign n565 = x62 & x94;
  assign n566 = x62 | x94;
  assign n567 = ~n565 & n566;
  assign n948 = n558 | n560;
  assign n949 = (n558 & n758) | (n558 & n948) | (n758 & n948);
  assign n769 = n567 & n949;
  assign n950 = n551 | n558;
  assign n951 = (n558 & n560) | (n558 & n950) | (n560 & n950);
  assign n770 = n567 & n951;
  assign n952 = (n769 & n770) | (n769 & n934) | (n770 & n934);
  assign n953 = (n769 & n770) | (n769 & n935) | (n770 & n935);
  assign n954 = (n928 & n952) | (n928 & n953) | (n952 & n953);
  assign n772 = n567 | n949;
  assign n773 = n567 | n951;
  assign n955 = (n772 & n773) | (n772 & n934) | (n773 & n934);
  assign n956 = (n772 & n773) | (n772 & n935) | (n773 & n935);
  assign n957 = (n928 & n955) | (n928 & n956) | (n955 & n956);
  assign n570 = ~n954 & n957;
  assign n572 = x63 & x95;
  assign n573 = x63 | x95;
  assign n574 = ~n572 & n573;
  assign n958 = n565 | n567;
  assign n963 = (n565 & n951) | (n565 & n958) | (n951 & n958);
  assign n779 = n574 & n963;
  assign n960 = n574 & n958;
  assign n961 = n565 & n574;
  assign n962 = (n949 & n960) | (n949 & n961) | (n960 & n961);
  assign n964 = (n779 & n934) | (n779 & n962) | (n934 & n962);
  assign n965 = (n779 & n935) | (n779 & n962) | (n935 & n962);
  assign n966 = (n928 & n964) | (n928 & n965) | (n964 & n965);
  assign n782 = n574 | n963;
  assign n967 = n574 | n958;
  assign n968 = n565 | n574;
  assign n969 = (n949 & n967) | (n949 & n968) | (n967 & n968);
  assign n970 = (n782 & n934) | (n782 & n969) | (n934 & n969);
  assign n971 = (n782 & n935) | (n782 & n969) | (n935 & n969);
  assign n972 = (n928 & n970) | (n928 & n971) | (n970 & n971);
  assign n577 = ~n966 & n972;
  assign n579 = x64 & x96;
  assign n580 = x64 | x96;
  assign n581 = ~n579 & n580;
  assign n784 = n572 & n581;
  assign n785 = (n581 & n966) | (n581 & n784) | (n966 & n784);
  assign n786 = n572 | n581;
  assign n787 = n966 | n786;
  assign n584 = ~n785 & n787;
  assign n586 = x65 & x97;
  assign n587 = x65 | x97;
  assign n588 = ~n586 & n587;
  assign n973 = n572 | n579;
  assign n974 = (n579 & n581) | (n579 & n973) | (n581 & n973);
  assign n791 = n588 & n974;
  assign n789 = n579 | n581;
  assign n792 = n588 & n789;
  assign n793 = (n966 & n791) | (n966 & n792) | (n791 & n792);
  assign n794 = n588 | n974;
  assign n795 = n588 | n789;
  assign n796 = (n966 & n794) | (n966 & n795) | (n794 & n795);
  assign n591 = ~n793 & n796;
  assign n593 = x66 & x98;
  assign n594 = x66 | x98;
  assign n595 = ~n593 & n594;
  assign n975 = n586 | n588;
  assign n976 = (n586 & n974) | (n586 & n975) | (n974 & n975);
  assign n800 = n595 & n976;
  assign n977 = (n586 & n789) | (n586 & n975) | (n789 & n975);
  assign n801 = n595 & n977;
  assign n802 = (n966 & n800) | (n966 & n801) | (n800 & n801);
  assign n803 = n595 | n976;
  assign n804 = n595 | n977;
  assign n805 = (n966 & n803) | (n966 & n804) | (n803 & n804);
  assign n598 = ~n802 & n805;
  assign n600 = x67 & x99;
  assign n601 = x67 | x99;
  assign n602 = ~n600 & n601;
  assign n978 = n593 | n595;
  assign n980 = n602 & n978;
  assign n981 = n593 & n602;
  assign n982 = (n976 & n980) | (n976 & n981) | (n980 & n981);
  assign n984 = (n977 & n980) | (n977 & n981) | (n980 & n981);
  assign n811 = (n966 & n982) | (n966 & n984) | (n982 & n984);
  assign n985 = n602 | n978;
  assign n986 = n593 | n602;
  assign n987 = (n976 & n985) | (n976 & n986) | (n985 & n986);
  assign n988 = (n977 & n985) | (n977 & n986) | (n985 & n986);
  assign n814 = (n966 & n987) | (n966 & n988) | (n987 & n988);
  assign n605 = ~n811 & n814;
  assign n607 = x68 & x100;
  assign n608 = x68 | x100;
  assign n609 = ~n607 & n608;
  assign n815 = n600 & n609;
  assign n989 = (n609 & n815) | (n609 & n984) | (n815 & n984);
  assign n990 = (n609 & n815) | (n609 & n982) | (n815 & n982);
  assign n991 = (n966 & n989) | (n966 & n990) | (n989 & n990);
  assign n817 = n600 | n609;
  assign n992 = n817 | n984;
  assign n993 = n817 | n982;
  assign n994 = (n966 & n992) | (n966 & n993) | (n992 & n993);
  assign n612 = ~n991 & n994;
  assign n614 = x69 & x101;
  assign n615 = x69 | x101;
  assign n616 = ~n614 & n615;
  assign n995 = n600 | n607;
  assign n996 = (n607 & n609) | (n607 & n995) | (n609 & n995);
  assign n822 = n616 & n996;
  assign n820 = n607 | n609;
  assign n823 = n616 & n820;
  assign n997 = (n822 & n823) | (n822 & n984) | (n823 & n984);
  assign n998 = (n822 & n823) | (n822 & n982) | (n823 & n982);
  assign n999 = (n966 & n997) | (n966 & n998) | (n997 & n998);
  assign n825 = n616 | n996;
  assign n826 = n616 | n820;
  assign n1000 = (n825 & n826) | (n825 & n984) | (n826 & n984);
  assign n1001 = (n825 & n826) | (n825 & n982) | (n826 & n982);
  assign n1002 = (n966 & n1000) | (n966 & n1001) | (n1000 & n1001);
  assign n619 = ~n999 & n1002;
  assign n621 = x70 & x102;
  assign n622 = x70 | x102;
  assign n623 = ~n621 & n622;
  assign n1003 = n614 | n616;
  assign n1004 = (n614 & n996) | (n614 & n1003) | (n996 & n1003);
  assign n831 = n623 & n1004;
  assign n1005 = (n614 & n820) | (n614 & n1003) | (n820 & n1003);
  assign n832 = n623 & n1005;
  assign n1006 = (n831 & n832) | (n831 & n984) | (n832 & n984);
  assign n1007 = (n831 & n832) | (n831 & n982) | (n832 & n982);
  assign n1008 = (n966 & n1006) | (n966 & n1007) | (n1006 & n1007);
  assign n834 = n623 | n1004;
  assign n835 = n623 | n1005;
  assign n1009 = (n834 & n835) | (n834 & n984) | (n835 & n984);
  assign n1010 = (n834 & n835) | (n834 & n982) | (n835 & n982);
  assign n1011 = (n966 & n1009) | (n966 & n1010) | (n1009 & n1010);
  assign n626 = ~n1008 & n1011;
  assign n628 = x71 & x103;
  assign n629 = x71 | x103;
  assign n630 = ~n628 & n629;
  assign n1012 = n621 | n623;
  assign n1014 = n630 & n1012;
  assign n1015 = n621 & n630;
  assign n1016 = (n1004 & n1014) | (n1004 & n1015) | (n1014 & n1015);
  assign n1018 = (n1005 & n1014) | (n1005 & n1015) | (n1014 & n1015);
  assign n1019 = (n984 & n1016) | (n984 & n1018) | (n1016 & n1018);
  assign n1020 = (n982 & n1016) | (n982 & n1018) | (n1016 & n1018);
  assign n1021 = (n966 & n1019) | (n966 & n1020) | (n1019 & n1020);
  assign n1022 = n630 | n1012;
  assign n1023 = n621 | n630;
  assign n1024 = (n1004 & n1022) | (n1004 & n1023) | (n1022 & n1023);
  assign n1025 = (n1005 & n1022) | (n1005 & n1023) | (n1022 & n1023);
  assign n1026 = (n984 & n1024) | (n984 & n1025) | (n1024 & n1025);
  assign n1027 = (n982 & n1024) | (n982 & n1025) | (n1024 & n1025);
  assign n1028 = (n966 & n1026) | (n966 & n1027) | (n1026 & n1027);
  assign n633 = ~n1021 & n1028;
  assign n846 = n628 | n1016;
  assign n847 = n628 | n1018;
  assign n1029 = (n846 & n847) | (n846 & n984) | (n847 & n984);
  assign n1030 = (n846 & n847) | (n846 & n982) | (n847 & n982);
  assign n1031 = (n966 & n1029) | (n966 & n1030) | (n1029 & n1030);
  assign n635 = x72 & x104;
  assign n636 = x72 | x104;
  assign n637 = ~n635 & n636;
  assign n638 = n1031 & n637;
  assign n639 = n1031 | n637;
  assign n640 = ~n638 & n639;
  assign n642 = x73 & x105;
  assign n643 = x73 | x105;
  assign n644 = ~n642 & n643;
  assign n849 = n635 | n637;
  assign n851 = n644 & n849;
  assign n852 = n635 & n644;
  assign n853 = (n1031 & n851) | (n1031 & n852) | (n851 & n852);
  assign n854 = n644 | n849;
  assign n855 = n635 | n644;
  assign n856 = (n1031 & n854) | (n1031 & n855) | (n854 & n855);
  assign n647 = ~n853 & n856;
  assign n649 = x74 & x106;
  assign n650 = x74 | x106;
  assign n651 = ~n649 & n650;
  assign n1032 = n642 | n644;
  assign n1033 = (n642 & n849) | (n642 & n1032) | (n849 & n1032);
  assign n860 = n651 & n1033;
  assign n1034 = n635 | n642;
  assign n1035 = (n642 & n644) | (n642 & n1034) | (n644 & n1034);
  assign n861 = n651 & n1035;
  assign n862 = (n1031 & n860) | (n1031 & n861) | (n860 & n861);
  assign n863 = n651 | n1033;
  assign n864 = n651 | n1035;
  assign n865 = (n1031 & n863) | (n1031 & n864) | (n863 & n864);
  assign n654 = ~n862 & n865;
  assign n656 = x75 & x107;
  assign n657 = x75 | x107;
  assign n658 = ~n656 & n657;
  assign n1036 = n649 | n651;
  assign n1038 = n658 & n1036;
  assign n1039 = n649 & n658;
  assign n1040 = (n1033 & n1038) | (n1033 & n1039) | (n1038 & n1039);
  assign n1041 = (n649 & n1035) | (n649 & n1036) | (n1035 & n1036);
  assign n870 = n658 & n1041;
  assign n871 = (n1031 & n1040) | (n1031 & n870) | (n1040 & n870);
  assign n1042 = n658 | n1036;
  assign n1043 = n649 | n658;
  assign n1044 = (n1033 & n1042) | (n1033 & n1043) | (n1042 & n1043);
  assign n873 = n658 | n1041;
  assign n874 = (n1031 & n1044) | (n1031 & n873) | (n1044 & n873);
  assign n661 = ~n871 & n874;
  assign n663 = x76 & x108;
  assign n664 = x76 | x108;
  assign n665 = ~n663 & n664;
  assign n1045 = n656 & n665;
  assign n1046 = (n665 & n1040) | (n665 & n1045) | (n1040 & n1045);
  assign n1047 = n656 | n658;
  assign n1049 = n665 & n1047;
  assign n1050 = (n1041 & n1045) | (n1041 & n1049) | (n1045 & n1049);
  assign n880 = (n1031 & n1046) | (n1031 & n1050) | (n1046 & n1050);
  assign n1051 = n656 | n665;
  assign n1052 = n1040 | n1051;
  assign n1053 = n665 | n1047;
  assign n1054 = (n1041 & n1051) | (n1041 & n1053) | (n1051 & n1053);
  assign n883 = (n1031 & n1052) | (n1031 & n1054) | (n1052 & n1054);
  assign n668 = ~n880 & n883;
  assign n670 = x77 & x109;
  assign n671 = x77 | x109;
  assign n672 = ~n670 & n671;
  assign n885 = n663 | n1050;
  assign n1058 = n672 & n885;
  assign n1055 = n663 | n1045;
  assign n1056 = n663 | n665;
  assign n1057 = (n1040 & n1055) | (n1040 & n1056) | (n1055 & n1056);
  assign n1059 = n672 & n1057;
  assign n1060 = (n1031 & n1058) | (n1031 & n1059) | (n1058 & n1059);
  assign n1061 = n672 | n885;
  assign n1062 = n672 | n1057;
  assign n1063 = (n1031 & n1061) | (n1031 & n1062) | (n1061 & n1062);
  assign n675 = ~n1060 & n1063;
  assign n677 = x78 & x110;
  assign n678 = x78 | x110;
  assign n679 = ~n677 & n678;
  assign n887 = n670 | n672;
  assign n889 = n679 & n887;
  assign n890 = n670 & n679;
  assign n1064 = (n885 & n889) | (n885 & n890) | (n889 & n890);
  assign n1065 = (n889 & n890) | (n889 & n1057) | (n890 & n1057);
  assign n1066 = (n1031 & n1064) | (n1031 & n1065) | (n1064 & n1065);
  assign n892 = n679 | n887;
  assign n893 = n670 | n679;
  assign n1067 = (n885 & n892) | (n885 & n893) | (n892 & n893);
  assign n1068 = (n892 & n893) | (n892 & n1057) | (n893 & n1057);
  assign n1069 = (n1031 & n1067) | (n1031 & n1068) | (n1067 & n1068);
  assign n682 = ~n1066 & n1069;
  assign n684 = x79 & x111;
  assign n685 = x79 | x111;
  assign n686 = ~n684 & n685;
  assign n1070 = n677 | n679;
  assign n1071 = (n677 & n887) | (n677 & n1070) | (n887 & n1070);
  assign n898 = n686 & n1071;
  assign n1072 = n670 | n677;
  assign n1073 = (n677 & n679) | (n677 & n1072) | (n679 & n1072);
  assign n899 = n686 & n1073;
  assign n1074 = (n885 & n898) | (n885 & n899) | (n898 & n899);
  assign n1075 = (n898 & n899) | (n898 & n1057) | (n899 & n1057);
  assign n1076 = (n1031 & n1074) | (n1031 & n1075) | (n1074 & n1075);
  assign n901 = n686 | n1071;
  assign n902 = n686 | n1073;
  assign n1077 = (n885 & n901) | (n885 & n902) | (n901 & n902);
  assign n1078 = (n901 & n902) | (n901 & n1057) | (n902 & n1057);
  assign n1079 = (n1031 & n1077) | (n1031 & n1078) | (n1077 & n1078);
  assign n689 = ~n1076 & n1079;
  assign n1080 = n684 | n686;
  assign n1081 = (n684 & n1071) | (n684 & n1080) | (n1071 & n1080);
  assign n1082 = (n684 & n1073) | (n684 & n1080) | (n1073 & n1080);
  assign n1083 = (n885 & n1081) | (n885 & n1082) | (n1081 & n1082);
  assign n1084 = (n1057 & n1081) | (n1057 & n1082) | (n1081 & n1082);
  assign n1085 = (n1031 & n1083) | (n1031 & n1084) | (n1083 & n1084);
  assign y0 = n19;
  assign y1 = n25;
  assign y2 = n32;
  assign y3 = n39;
  assign y4 = n46;
  assign y5 = n53;
  assign y6 = n60;
  assign y7 = n67;
  assign y8 = n113;
  assign y9 = n148;
  assign y10 = n154;
  assign y11 = n161;
  assign y12 = n168;
  assign y13 = n175;
  assign y14 = n182;
  assign y15 = n189;
  assign y16 = n196;
  assign y17 = n203;
  assign y18 = n210;
  assign y19 = n217;
  assign y20 = n224;
  assign y21 = n231;
  assign y22 = n238;
  assign y23 = n245;
  assign y24 = n252;
  assign y25 = n253;
  assign y26 = n473;
  assign y27 = n479;
  assign y28 = n486;
  assign y29 = n493;
  assign y30 = n500;
  assign y31 = n507;
  assign y32 = n514;
  assign y33 = n521;
  assign y34 = n528;
  assign y35 = n535;
  assign y36 = n542;
  assign y37 = n549;
  assign y38 = n556;
  assign y39 = n563;
  assign y40 = n570;
  assign y41 = n577;
  assign y42 = n584;
  assign y43 = n591;
  assign y44 = n598;
  assign y45 = n605;
  assign y46 = n612;
  assign y47 = n619;
  assign y48 = n626;
  assign y49 = n633;
  assign y50 = n640;
  assign y51 = n647;
  assign y52 = n654;
  assign y53 = n661;
  assign y54 = n668;
  assign y55 = n675;
  assign y56 = n682;
  assign y57 = n689;
  assign y58 = n1085;
endmodule

