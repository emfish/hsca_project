module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406;
  assign n17 = x0 & x8;
  assign n18 = x0 | x8;
  assign n19 = ~n17 & n18;
  assign n20 = x1 & x9;
  assign n21 = x1 | x9;
  assign n22 = ~n20 & n21;
  assign n23 = n17 & n22;
  assign n24 = n17 | n22;
  assign n25 = ~n23 & n24;
  assign n69 = n17 | n20;
  assign n70 = (n20 & n22) | (n20 & n69) | (n22 & n69);
  assign n27 = x2 & x10;
  assign n28 = x2 | x10;
  assign n29 = ~n27 & n28;
  assign n30 = n70 & n29;
  assign n31 = n70 | n29;
  assign n32 = ~n30 & n31;
  assign n71 = n27 | n29;
  assign n72 = (n27 & n70) | (n27 & n71) | (n70 & n71);
  assign n34 = x3 & x11;
  assign n35 = x3 | x11;
  assign n36 = ~n34 & n35;
  assign n37 = n72 & n36;
  assign n38 = n72 | n36;
  assign n39 = ~n37 & n38;
  assign n41 = x4 & x12;
  assign n42 = x4 | x12;
  assign n43 = ~n41 & n42;
  assign n73 = n34 | n36;
  assign n75 = n43 & n73;
  assign n76 = n34 & n43;
  assign n77 = (n72 & n75) | (n72 & n76) | (n75 & n76);
  assign n78 = n43 | n73;
  assign n79 = n34 | n43;
  assign n80 = (n72 & n78) | (n72 & n79) | (n78 & n79);
  assign n46 = ~n77 & n80;
  assign n48 = x5 & x13;
  assign n49 = x5 | x13;
  assign n50 = ~n48 & n49;
  assign n81 = n41 & n50;
  assign n82 = (n50 & n77) | (n50 & n81) | (n77 & n81);
  assign n83 = n41 | n50;
  assign n84 = n77 | n83;
  assign n53 = ~n82 & n84;
  assign n55 = x6 & x14;
  assign n56 = x6 | x14;
  assign n57 = ~n55 & n56;
  assign n101 = n41 | n48;
  assign n102 = (n48 & n50) | (n48 & n101) | (n50 & n101);
  assign n88 = n57 & n102;
  assign n86 = n48 | n50;
  assign n89 = n57 & n86;
  assign n90 = (n77 & n88) | (n77 & n89) | (n88 & n89);
  assign n91 = n57 | n102;
  assign n92 = n57 | n86;
  assign n93 = (n77 & n91) | (n77 & n92) | (n91 & n92);
  assign n60 = ~n90 & n93;
  assign n62 = x7 & x15;
  assign n63 = x7 | x15;
  assign n64 = ~n62 & n63;
  assign n94 = n55 & n64;
  assign n103 = (n64 & n89) | (n64 & n94) | (n89 & n94);
  assign n104 = (n64 & n88) | (n64 & n94) | (n88 & n94);
  assign n105 = (n77 & n103) | (n77 & n104) | (n103 & n104);
  assign n96 = n55 | n64;
  assign n106 = n89 | n96;
  assign n107 = n88 | n96;
  assign n108 = (n77 & n106) | (n77 & n107) | (n106 & n107);
  assign n67 = ~n105 & n108;
  assign n99 = n62 | n64;
  assign n109 = n55 | n62;
  assign n110 = (n62 & n64) | (n62 & n109) | (n64 & n109);
  assign n111 = (n89 & n99) | (n89 & n110) | (n99 & n110);
  assign n112 = (n88 & n99) | (n88 & n110) | (n99 & n110);
  assign n113 = (n77 & n111) | (n77 & n112) | (n111 & n112);
  assign n146 = x16 & x32;
  assign n147 = x16 | x32;
  assign n148 = ~n146 & n147;
  assign n149 = x17 & x33;
  assign n150 = x17 | x33;
  assign n151 = ~n149 & n150;
  assign n152 = n146 & n151;
  assign n153 = n146 | n151;
  assign n154 = ~n152 & n153;
  assign n254 = n146 | n149;
  assign n255 = (n149 & n151) | (n149 & n254) | (n151 & n254);
  assign n156 = x18 & x34;
  assign n157 = x18 | x34;
  assign n158 = ~n156 & n157;
  assign n159 = n255 & n158;
  assign n160 = n255 | n158;
  assign n161 = ~n159 & n160;
  assign n256 = n156 | n158;
  assign n257 = (n156 & n255) | (n156 & n256) | (n255 & n256);
  assign n163 = x19 & x35;
  assign n164 = x19 | x35;
  assign n165 = ~n163 & n164;
  assign n166 = n257 & n165;
  assign n167 = n257 | n165;
  assign n168 = ~n166 & n167;
  assign n170 = x20 & x36;
  assign n171 = x20 | x36;
  assign n172 = ~n170 & n171;
  assign n258 = n163 | n165;
  assign n260 = n172 & n258;
  assign n261 = n163 & n172;
  assign n262 = (n257 & n260) | (n257 & n261) | (n260 & n261);
  assign n263 = n172 | n258;
  assign n264 = n163 | n172;
  assign n265 = (n257 & n263) | (n257 & n264) | (n263 & n264);
  assign n175 = ~n262 & n265;
  assign n177 = x21 & x37;
  assign n178 = x21 | x37;
  assign n179 = ~n177 & n178;
  assign n266 = n170 & n179;
  assign n267 = (n179 & n262) | (n179 & n266) | (n262 & n266);
  assign n268 = n170 | n179;
  assign n269 = n262 | n268;
  assign n182 = ~n267 & n269;
  assign n184 = x22 & x38;
  assign n185 = x22 | x38;
  assign n186 = ~n184 & n185;
  assign n341 = n170 | n177;
  assign n342 = (n177 & n179) | (n177 & n341) | (n179 & n341);
  assign n273 = n186 & n342;
  assign n271 = n177 | n179;
  assign n274 = n186 & n271;
  assign n275 = (n262 & n273) | (n262 & n274) | (n273 & n274);
  assign n276 = n186 | n342;
  assign n277 = n186 | n271;
  assign n278 = (n262 & n276) | (n262 & n277) | (n276 & n277);
  assign n189 = ~n275 & n278;
  assign n191 = x23 & x39;
  assign n192 = x23 | x39;
  assign n193 = ~n191 & n192;
  assign n279 = n184 & n193;
  assign n343 = (n193 & n274) | (n193 & n279) | (n274 & n279);
  assign n344 = (n193 & n273) | (n193 & n279) | (n273 & n279);
  assign n345 = (n262 & n343) | (n262 & n344) | (n343 & n344);
  assign n281 = n184 | n193;
  assign n346 = n274 | n281;
  assign n347 = n273 | n281;
  assign n348 = (n262 & n346) | (n262 & n347) | (n346 & n347);
  assign n196 = ~n345 & n348;
  assign n198 = x24 & x40;
  assign n199 = x24 | x40;
  assign n200 = ~n198 & n199;
  assign n349 = n184 | n191;
  assign n350 = (n191 & n193) | (n191 & n349) | (n193 & n349);
  assign n286 = n200 & n350;
  assign n284 = n191 | n193;
  assign n287 = n200 & n284;
  assign n351 = (n274 & n286) | (n274 & n287) | (n286 & n287);
  assign n352 = (n273 & n286) | (n273 & n287) | (n286 & n287);
  assign n353 = (n262 & n351) | (n262 & n352) | (n351 & n352);
  assign n289 = n200 | n350;
  assign n290 = n200 | n284;
  assign n354 = (n274 & n289) | (n274 & n290) | (n289 & n290);
  assign n355 = (n273 & n289) | (n273 & n290) | (n289 & n290);
  assign n356 = (n262 & n354) | (n262 & n355) | (n354 & n355);
  assign n203 = ~n353 & n356;
  assign n357 = n198 | n200;
  assign n358 = (n198 & n350) | (n198 & n357) | (n350 & n357);
  assign n359 = (n198 & n284) | (n198 & n357) | (n284 & n357);
  assign n360 = (n274 & n358) | (n274 & n359) | (n358 & n359);
  assign n361 = (n273 & n358) | (n273 & n359) | (n358 & n359);
  assign n362 = (n262 & n360) | (n262 & n361) | (n360 & n361);
  assign n205 = x25 & x41;
  assign n206 = x25 | x41;
  assign n207 = ~n205 & n206;
  assign n208 = n362 & n207;
  assign n209 = n362 | n207;
  assign n210 = ~n208 & n209;
  assign n212 = x26 & x42;
  assign n213 = x26 | x42;
  assign n214 = ~n212 & n213;
  assign n295 = n205 | n207;
  assign n297 = n214 & n295;
  assign n298 = n205 & n214;
  assign n299 = (n362 & n297) | (n362 & n298) | (n297 & n298);
  assign n300 = n214 | n295;
  assign n301 = n205 | n214;
  assign n302 = (n362 & n300) | (n362 & n301) | (n300 & n301);
  assign n217 = ~n299 & n302;
  assign n219 = x27 & x43;
  assign n220 = x27 | x43;
  assign n221 = ~n219 & n220;
  assign n363 = n212 | n214;
  assign n364 = (n212 & n295) | (n212 & n363) | (n295 & n363);
  assign n306 = n221 & n364;
  assign n365 = n205 | n212;
  assign n366 = (n212 & n214) | (n212 & n365) | (n214 & n365);
  assign n307 = n221 & n366;
  assign n308 = (n362 & n306) | (n362 & n307) | (n306 & n307);
  assign n309 = n221 | n364;
  assign n310 = n221 | n366;
  assign n311 = (n362 & n309) | (n362 & n310) | (n309 & n310);
  assign n224 = ~n308 & n311;
  assign n226 = x28 & x44;
  assign n227 = x28 | x44;
  assign n228 = ~n226 & n227;
  assign n367 = n219 | n221;
  assign n368 = (n219 & n364) | (n219 & n367) | (n364 & n367);
  assign n370 = n228 & n368;
  assign n369 = (n219 & n366) | (n219 & n367) | (n366 & n367);
  assign n371 = n228 & n369;
  assign n372 = (n362 & n370) | (n362 & n371) | (n370 & n371);
  assign n373 = n228 | n368;
  assign n374 = n228 | n369;
  assign n375 = (n362 & n373) | (n362 & n374) | (n373 & n374);
  assign n231 = ~n372 & n375;
  assign n233 = x29 & x45;
  assign n234 = x29 | x45;
  assign n235 = ~n233 & n234;
  assign n315 = n226 | n228;
  assign n317 = n235 & n315;
  assign n318 = n226 & n235;
  assign n376 = (n317 & n318) | (n317 & n368) | (n318 & n368);
  assign n377 = (n317 & n318) | (n317 & n369) | (n318 & n369);
  assign n378 = (n362 & n376) | (n362 & n377) | (n376 & n377);
  assign n320 = n235 | n315;
  assign n321 = n226 | n235;
  assign n379 = (n320 & n321) | (n320 & n368) | (n321 & n368);
  assign n380 = (n320 & n321) | (n320 & n369) | (n321 & n369);
  assign n381 = (n362 & n379) | (n362 & n380) | (n379 & n380);
  assign n238 = ~n378 & n381;
  assign n240 = x30 & x46;
  assign n241 = x30 | x46;
  assign n242 = ~n240 & n241;
  assign n382 = n233 | n235;
  assign n383 = (n233 & n315) | (n233 & n382) | (n315 & n382);
  assign n326 = n242 & n383;
  assign n384 = n226 | n233;
  assign n385 = (n233 & n235) | (n233 & n384) | (n235 & n384);
  assign n327 = n242 & n385;
  assign n386 = (n326 & n327) | (n326 & n368) | (n327 & n368);
  assign n387 = (n326 & n327) | (n326 & n369) | (n327 & n369);
  assign n388 = (n362 & n386) | (n362 & n387) | (n386 & n387);
  assign n329 = n242 | n383;
  assign n330 = n242 | n385;
  assign n389 = (n329 & n330) | (n329 & n368) | (n330 & n368);
  assign n390 = (n329 & n330) | (n329 & n369) | (n330 & n369);
  assign n391 = (n362 & n389) | (n362 & n390) | (n389 & n390);
  assign n245 = ~n388 & n391;
  assign n247 = x31 & x47;
  assign n248 = x31 | x47;
  assign n249 = ~n247 & n248;
  assign n392 = n240 | n242;
  assign n397 = (n240 & n385) | (n240 & n392) | (n385 & n392);
  assign n336 = n249 & n397;
  assign n394 = n249 & n392;
  assign n395 = n240 & n249;
  assign n396 = (n383 & n394) | (n383 & n395) | (n394 & n395);
  assign n398 = (n336 & n368) | (n336 & n396) | (n368 & n396);
  assign n399 = (n336 & n369) | (n336 & n396) | (n369 & n396);
  assign n400 = (n362 & n398) | (n362 & n399) | (n398 & n399);
  assign n339 = n249 | n397;
  assign n401 = n249 | n392;
  assign n402 = n240 | n249;
  assign n403 = (n383 & n401) | (n383 & n402) | (n401 & n402);
  assign n404 = (n339 & n368) | (n339 & n403) | (n368 & n403);
  assign n405 = (n339 & n369) | (n339 & n403) | (n369 & n403);
  assign n406 = (n362 & n404) | (n362 & n405) | (n404 & n405);
  assign n252 = ~n400 & n406;
  assign n253 = n247 | n400;
  assign y0 = n19;
  assign y1 = n25;
  assign y2 = n32;
  assign y3 = n39;
  assign y4 = n46;
  assign y5 = n53;
  assign y6 = n60;
  assign y7 = n67;
  assign y8 = n113;
  assign y9 = n148;
  assign y10 = n154;
  assign y11 = n161;
  assign y12 = n168;
  assign y13 = n175;
  assign y14 = n182;
  assign y15 = n189;
  assign y16 = n196;
  assign y17 = n203;
  assign y18 = n210;
  assign y19 = n217;
  assign y20 = n224;
  assign y21 = n231;
  assign y22 = n238;
  assign y23 = n245;
  assign y24 = n252;
  assign y25 = n253;
endmodule

