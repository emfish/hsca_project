module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, y0, y1, y2, y3, y4, y5, y6, y7, y8);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113;
  assign n17 = x0 & x8;
  assign n18 = x0 | x8;
  assign n19 = ~n17 & n18;
  assign n20 = x1 & x9;
  assign n21 = x1 | x9;
  assign n22 = ~n20 & n21;
  assign n23 = n17 & n22;
  assign n24 = n17 | n22;
  assign n25 = ~n23 & n24;
  assign n69 = n17 | n20;
  assign n70 = (n20 & n22) | (n20 & n69) | (n22 & n69);
  assign n27 = x2 & x10;
  assign n28 = x2 | x10;
  assign n29 = ~n27 & n28;
  assign n30 = n70 & n29;
  assign n31 = n70 | n29;
  assign n32 = ~n30 & n31;
  assign n71 = n27 | n29;
  assign n72 = (n27 & n70) | (n27 & n71) | (n70 & n71);
  assign n34 = x3 & x11;
  assign n35 = x3 | x11;
  assign n36 = ~n34 & n35;
  assign n37 = n72 & n36;
  assign n38 = n72 | n36;
  assign n39 = ~n37 & n38;
  assign n41 = x4 & x12;
  assign n42 = x4 | x12;
  assign n43 = ~n41 & n42;
  assign n73 = n34 | n36;
  assign n75 = n43 & n73;
  assign n76 = n34 & n43;
  assign n77 = (n72 & n75) | (n72 & n76) | (n75 & n76);
  assign n78 = n43 | n73;
  assign n79 = n34 | n43;
  assign n80 = (n72 & n78) | (n72 & n79) | (n78 & n79);
  assign n46 = ~n77 & n80;
  assign n48 = x5 & x13;
  assign n49 = x5 | x13;
  assign n50 = ~n48 & n49;
  assign n81 = n41 & n50;
  assign n82 = (n50 & n77) | (n50 & n81) | (n77 & n81);
  assign n83 = n41 | n50;
  assign n84 = n77 | n83;
  assign n53 = ~n82 & n84;
  assign n55 = x6 & x14;
  assign n56 = x6 | x14;
  assign n57 = ~n55 & n56;
  assign n101 = n41 | n48;
  assign n102 = (n48 & n50) | (n48 & n101) | (n50 & n101);
  assign n88 = n57 & n102;
  assign n86 = n48 | n50;
  assign n89 = n57 & n86;
  assign n90 = (n77 & n88) | (n77 & n89) | (n88 & n89);
  assign n91 = n57 | n102;
  assign n92 = n57 | n86;
  assign n93 = (n77 & n91) | (n77 & n92) | (n91 & n92);
  assign n60 = ~n90 & n93;
  assign n62 = x7 & x15;
  assign n63 = x7 | x15;
  assign n64 = ~n62 & n63;
  assign n94 = n55 & n64;
  assign n103 = (n64 & n89) | (n64 & n94) | (n89 & n94);
  assign n104 = (n64 & n88) | (n64 & n94) | (n88 & n94);
  assign n105 = (n77 & n103) | (n77 & n104) | (n103 & n104);
  assign n96 = n55 | n64;
  assign n106 = n89 | n96;
  assign n107 = n88 | n96;
  assign n108 = (n77 & n106) | (n77 & n107) | (n106 & n107);
  assign n67 = ~n105 & n108;
  assign n99 = n62 | n64;
  assign n109 = n55 | n62;
  assign n110 = (n62 & n64) | (n62 & n109) | (n64 & n109);
  assign n111 = (n89 & n99) | (n89 & n110) | (n99 & n110);
  assign n112 = (n88 & n99) | (n88 & n110) | (n99 & n110);
  assign n113 = (n77 & n111) | (n77 & n112) | (n111 & n112);
  assign y0 = n19;
  assign y1 = n25;
  assign y2 = n32;
  assign y3 = n39;
  assign y4 = n46;
  assign y5 = n53;
  assign y6 = n60;
  assign y7 = n67;
  assign y8 = n113;
endmodule

