module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792;
  assign n17 = x0 & x8;
  assign n18 = x0 | x8;
  assign n19 = ~n17 & n18;
  assign n20 = x1 & x9;
  assign n21 = x1 | x9;
  assign n22 = ~n20 & n21;
  assign n23 = n17 & n22;
  assign n24 = n17 | n22;
  assign n25 = ~n23 & n24;
  assign n69 = n17 | n20;
  assign n70 = (n20 & n22) | (n20 & n69) | (n22 & n69);
  assign n27 = x2 & x10;
  assign n28 = x2 | x10;
  assign n29 = ~n27 & n28;
  assign n30 = n70 & n29;
  assign n31 = n70 | n29;
  assign n32 = ~n30 & n31;
  assign n71 = n27 | n29;
  assign n72 = (n27 & n70) | (n27 & n71) | (n70 & n71);
  assign n34 = x3 & x11;
  assign n35 = x3 | x11;
  assign n36 = ~n34 & n35;
  assign n37 = n72 & n36;
  assign n38 = n72 | n36;
  assign n39 = ~n37 & n38;
  assign n41 = x4 & x12;
  assign n42 = x4 | x12;
  assign n43 = ~n41 & n42;
  assign n73 = n34 | n36;
  assign n75 = n43 & n73;
  assign n76 = n34 & n43;
  assign n77 = (n72 & n75) | (n72 & n76) | (n75 & n76);
  assign n78 = n43 | n73;
  assign n79 = n34 | n43;
  assign n80 = (n72 & n78) | (n72 & n79) | (n78 & n79);
  assign n46 = ~n77 & n80;
  assign n48 = x5 & x13;
  assign n49 = x5 | x13;
  assign n50 = ~n48 & n49;
  assign n81 = n41 & n50;
  assign n82 = (n50 & n77) | (n50 & n81) | (n77 & n81);
  assign n83 = n41 | n50;
  assign n84 = n77 | n83;
  assign n53 = ~n82 & n84;
  assign n55 = x6 & x14;
  assign n56 = x6 | x14;
  assign n57 = ~n55 & n56;
  assign n101 = n41 | n48;
  assign n102 = (n48 & n50) | (n48 & n101) | (n50 & n101);
  assign n88 = n57 & n102;
  assign n86 = n48 | n50;
  assign n89 = n57 & n86;
  assign n90 = (n77 & n88) | (n77 & n89) | (n88 & n89);
  assign n91 = n57 | n102;
  assign n92 = n57 | n86;
  assign n93 = (n77 & n91) | (n77 & n92) | (n91 & n92);
  assign n60 = ~n90 & n93;
  assign n62 = x7 & x15;
  assign n63 = x7 | x15;
  assign n64 = ~n62 & n63;
  assign n94 = n55 & n64;
  assign n103 = (n64 & n89) | (n64 & n94) | (n89 & n94);
  assign n104 = (n64 & n88) | (n64 & n94) | (n88 & n94);
  assign n105 = (n77 & n103) | (n77 & n104) | (n103 & n104);
  assign n96 = n55 | n64;
  assign n106 = n89 | n96;
  assign n107 = n88 | n96;
  assign n108 = (n77 & n106) | (n77 & n107) | (n106 & n107);
  assign n67 = ~n105 & n108;
  assign n99 = n62 | n64;
  assign n109 = n55 | n62;
  assign n110 = (n62 & n64) | (n62 & n109) | (n64 & n109);
  assign n111 = (n89 & n99) | (n89 & n110) | (n99 & n110);
  assign n112 = (n88 & n99) | (n88 & n110) | (n99 & n110);
  assign n113 = (n77 & n111) | (n77 & n112) | (n111 & n112);
  assign n146 = x16 & x32;
  assign n147 = x16 | x32;
  assign n148 = ~n146 & n147;
  assign n149 = x17 & x33;
  assign n150 = x17 | x33;
  assign n151 = ~n149 & n150;
  assign n152 = n146 & n151;
  assign n153 = n146 | n151;
  assign n154 = ~n152 & n153;
  assign n254 = n146 | n149;
  assign n255 = (n149 & n151) | (n149 & n254) | (n151 & n254);
  assign n156 = x18 & x34;
  assign n157 = x18 | x34;
  assign n158 = ~n156 & n157;
  assign n159 = n255 & n158;
  assign n160 = n255 | n158;
  assign n161 = ~n159 & n160;
  assign n256 = n156 | n158;
  assign n257 = (n156 & n255) | (n156 & n256) | (n255 & n256);
  assign n163 = x19 & x35;
  assign n164 = x19 | x35;
  assign n165 = ~n163 & n164;
  assign n166 = n257 & n165;
  assign n167 = n257 | n165;
  assign n168 = ~n166 & n167;
  assign n170 = x20 & x36;
  assign n171 = x20 | x36;
  assign n172 = ~n170 & n171;
  assign n258 = n163 | n165;
  assign n260 = n172 & n258;
  assign n261 = n163 & n172;
  assign n262 = (n257 & n260) | (n257 & n261) | (n260 & n261);
  assign n263 = n172 | n258;
  assign n264 = n163 | n172;
  assign n265 = (n257 & n263) | (n257 & n264) | (n263 & n264);
  assign n175 = ~n262 & n265;
  assign n177 = x21 & x37;
  assign n178 = x21 | x37;
  assign n179 = ~n177 & n178;
  assign n266 = n170 & n179;
  assign n267 = (n179 & n262) | (n179 & n266) | (n262 & n266);
  assign n268 = n170 | n179;
  assign n269 = n262 | n268;
  assign n182 = ~n267 & n269;
  assign n184 = x22 & x38;
  assign n185 = x22 | x38;
  assign n186 = ~n184 & n185;
  assign n341 = n170 | n177;
  assign n342 = (n177 & n179) | (n177 & n341) | (n179 & n341);
  assign n273 = n186 & n342;
  assign n271 = n177 | n179;
  assign n274 = n186 & n271;
  assign n275 = (n262 & n273) | (n262 & n274) | (n273 & n274);
  assign n276 = n186 | n342;
  assign n277 = n186 | n271;
  assign n278 = (n262 & n276) | (n262 & n277) | (n276 & n277);
  assign n189 = ~n275 & n278;
  assign n191 = x23 & x39;
  assign n192 = x23 | x39;
  assign n193 = ~n191 & n192;
  assign n279 = n184 & n193;
  assign n343 = (n193 & n274) | (n193 & n279) | (n274 & n279);
  assign n344 = (n193 & n273) | (n193 & n279) | (n273 & n279);
  assign n345 = (n262 & n343) | (n262 & n344) | (n343 & n344);
  assign n281 = n184 | n193;
  assign n346 = n274 | n281;
  assign n347 = n273 | n281;
  assign n348 = (n262 & n346) | (n262 & n347) | (n346 & n347);
  assign n196 = ~n345 & n348;
  assign n198 = x24 & x40;
  assign n199 = x24 | x40;
  assign n200 = ~n198 & n199;
  assign n349 = n184 | n191;
  assign n350 = (n191 & n193) | (n191 & n349) | (n193 & n349);
  assign n286 = n200 & n350;
  assign n284 = n191 | n193;
  assign n287 = n200 & n284;
  assign n351 = (n274 & n286) | (n274 & n287) | (n286 & n287);
  assign n352 = (n273 & n286) | (n273 & n287) | (n286 & n287);
  assign n353 = (n262 & n351) | (n262 & n352) | (n351 & n352);
  assign n289 = n200 | n350;
  assign n290 = n200 | n284;
  assign n354 = (n274 & n289) | (n274 & n290) | (n289 & n290);
  assign n355 = (n273 & n289) | (n273 & n290) | (n289 & n290);
  assign n356 = (n262 & n354) | (n262 & n355) | (n354 & n355);
  assign n203 = ~n353 & n356;
  assign n357 = n198 | n200;
  assign n358 = (n198 & n350) | (n198 & n357) | (n350 & n357);
  assign n359 = (n198 & n284) | (n198 & n357) | (n284 & n357);
  assign n360 = (n274 & n358) | (n274 & n359) | (n358 & n359);
  assign n361 = (n273 & n358) | (n273 & n359) | (n358 & n359);
  assign n362 = (n262 & n360) | (n262 & n361) | (n360 & n361);
  assign n205 = x25 & x41;
  assign n206 = x25 | x41;
  assign n207 = ~n205 & n206;
  assign n208 = n362 & n207;
  assign n209 = n362 | n207;
  assign n210 = ~n208 & n209;
  assign n212 = x26 & x42;
  assign n213 = x26 | x42;
  assign n214 = ~n212 & n213;
  assign n295 = n205 | n207;
  assign n297 = n214 & n295;
  assign n298 = n205 & n214;
  assign n299 = (n362 & n297) | (n362 & n298) | (n297 & n298);
  assign n300 = n214 | n295;
  assign n301 = n205 | n214;
  assign n302 = (n362 & n300) | (n362 & n301) | (n300 & n301);
  assign n217 = ~n299 & n302;
  assign n219 = x27 & x43;
  assign n220 = x27 | x43;
  assign n221 = ~n219 & n220;
  assign n363 = n212 | n214;
  assign n364 = (n212 & n295) | (n212 & n363) | (n295 & n363);
  assign n306 = n221 & n364;
  assign n365 = n205 | n212;
  assign n366 = (n212 & n214) | (n212 & n365) | (n214 & n365);
  assign n307 = n221 & n366;
  assign n308 = (n362 & n306) | (n362 & n307) | (n306 & n307);
  assign n309 = n221 | n364;
  assign n310 = n221 | n366;
  assign n311 = (n362 & n309) | (n362 & n310) | (n309 & n310);
  assign n224 = ~n308 & n311;
  assign n226 = x28 & x44;
  assign n227 = x28 | x44;
  assign n228 = ~n226 & n227;
  assign n367 = n219 | n221;
  assign n691 = n228 & n367;
  assign n692 = n219 & n228;
  assign n693 = (n364 & n691) | (n364 & n692) | (n691 & n692);
  assign n369 = (n219 & n366) | (n219 & n367) | (n366 & n367);
  assign n371 = n228 & n369;
  assign n372 = (n362 & n693) | (n362 & n371) | (n693 & n371);
  assign n694 = n228 | n367;
  assign n695 = n219 | n228;
  assign n696 = (n364 & n694) | (n364 & n695) | (n694 & n695);
  assign n374 = n228 | n369;
  assign n375 = (n362 & n696) | (n362 & n374) | (n696 & n374);
  assign n231 = ~n372 & n375;
  assign n233 = x29 & x45;
  assign n234 = x29 | x45;
  assign n235 = ~n233 & n234;
  assign n315 = n226 | n228;
  assign n317 = n235 & n315;
  assign n318 = n226 & n235;
  assign n368 = (n219 & n364) | (n219 & n367) | (n364 & n367);
  assign n376 = (n317 & n318) | (n317 & n368) | (n318 & n368);
  assign n377 = (n317 & n318) | (n317 & n369) | (n318 & n369);
  assign n378 = (n362 & n376) | (n362 & n377) | (n376 & n377);
  assign n320 = n235 | n315;
  assign n321 = n226 | n235;
  assign n379 = (n320 & n321) | (n320 & n368) | (n321 & n368);
  assign n380 = (n320 & n321) | (n320 & n369) | (n321 & n369);
  assign n381 = (n362 & n379) | (n362 & n380) | (n379 & n380);
  assign n238 = ~n378 & n381;
  assign n240 = x30 & x46;
  assign n241 = x30 | x46;
  assign n242 = ~n240 & n241;
  assign n382 = n233 | n235;
  assign n383 = (n233 & n315) | (n233 & n382) | (n315 & n382);
  assign n326 = n242 & n383;
  assign n384 = n226 | n233;
  assign n385 = (n233 & n235) | (n233 & n384) | (n235 & n384);
  assign n327 = n242 & n385;
  assign n386 = (n326 & n327) | (n326 & n368) | (n327 & n368);
  assign n387 = (n326 & n327) | (n326 & n369) | (n327 & n369);
  assign n388 = (n362 & n386) | (n362 & n387) | (n386 & n387);
  assign n329 = n242 | n383;
  assign n330 = n242 | n385;
  assign n389 = (n329 & n330) | (n329 & n368) | (n330 & n368);
  assign n390 = (n329 & n330) | (n329 & n369) | (n330 & n369);
  assign n391 = (n362 & n389) | (n362 & n390) | (n389 & n390);
  assign n245 = ~n388 & n391;
  assign n247 = x31 & x47;
  assign n248 = x31 | x47;
  assign n249 = ~n247 & n248;
  assign n392 = n240 | n242;
  assign n397 = (n240 & n385) | (n240 & n392) | (n385 & n392);
  assign n336 = n249 & n397;
  assign n394 = n249 & n392;
  assign n395 = n240 & n249;
  assign n396 = (n383 & n394) | (n383 & n395) | (n394 & n395);
  assign n398 = (n336 & n368) | (n336 & n396) | (n368 & n396);
  assign n399 = (n336 & n369) | (n336 & n396) | (n369 & n396);
  assign n400 = (n362 & n398) | (n362 & n399) | (n398 & n399);
  assign n339 = n249 | n397;
  assign n401 = n249 | n392;
  assign n402 = n240 | n249;
  assign n403 = (n383 & n401) | (n383 & n402) | (n401 & n402);
  assign n404 = (n339 & n368) | (n339 & n403) | (n368 & n403);
  assign n405 = (n339 & n369) | (n339 & n403) | (n369 & n403);
  assign n406 = (n362 & n404) | (n362 & n405) | (n404 & n405);
  assign n252 = ~n400 & n406;
  assign n253 = n247 | n400;
  assign n471 = x48 & x80;
  assign n472 = x48 | x80;
  assign n473 = ~n471 & n472;
  assign n474 = x49 & x81;
  assign n475 = x49 | x81;
  assign n476 = ~n474 & n475;
  assign n477 = n471 & n476;
  assign n478 = n471 | n476;
  assign n479 = ~n477 & n478;
  assign n697 = n471 | n474;
  assign n698 = (n474 & n476) | (n474 & n697) | (n476 & n697);
  assign n481 = x50 & x82;
  assign n482 = x50 | x82;
  assign n483 = ~n481 & n482;
  assign n484 = n698 & n483;
  assign n485 = n698 | n483;
  assign n486 = ~n484 & n485;
  assign n699 = n481 | n483;
  assign n700 = (n481 & n698) | (n481 & n699) | (n698 & n699);
  assign n488 = x51 & x83;
  assign n489 = x51 | x83;
  assign n490 = ~n488 & n489;
  assign n491 = n700 & n490;
  assign n492 = n700 | n490;
  assign n493 = ~n491 & n492;
  assign n495 = x52 & x84;
  assign n496 = x52 | x84;
  assign n497 = ~n495 & n496;
  assign n701 = n488 | n490;
  assign n703 = n497 & n701;
  assign n704 = n488 & n497;
  assign n705 = (n700 & n703) | (n700 & n704) | (n703 & n704);
  assign n706 = n497 | n701;
  assign n707 = n488 | n497;
  assign n708 = (n700 & n706) | (n700 & n707) | (n706 & n707);
  assign n500 = ~n705 & n708;
  assign n502 = x53 & x85;
  assign n503 = x53 | x85;
  assign n504 = ~n502 & n503;
  assign n709 = n495 & n504;
  assign n710 = (n504 & n705) | (n504 & n709) | (n705 & n709);
  assign n711 = n495 | n504;
  assign n712 = n705 | n711;
  assign n507 = ~n710 & n712;
  assign n509 = x54 & x86;
  assign n510 = x54 | x86;
  assign n511 = ~n509 & n510;
  assign n907 = n495 | n502;
  assign n908 = (n502 & n504) | (n502 & n907) | (n504 & n907);
  assign n716 = n511 & n908;
  assign n714 = n502 | n504;
  assign n717 = n511 & n714;
  assign n718 = (n705 & n716) | (n705 & n717) | (n716 & n717);
  assign n719 = n511 | n908;
  assign n720 = n511 | n714;
  assign n721 = (n705 & n719) | (n705 & n720) | (n719 & n720);
  assign n514 = ~n718 & n721;
  assign n516 = x55 & x87;
  assign n517 = x55 | x87;
  assign n518 = ~n516 & n517;
  assign n722 = n509 & n518;
  assign n909 = (n518 & n717) | (n518 & n722) | (n717 & n722);
  assign n910 = (n518 & n716) | (n518 & n722) | (n716 & n722);
  assign n911 = (n705 & n909) | (n705 & n910) | (n909 & n910);
  assign n724 = n509 | n518;
  assign n912 = n717 | n724;
  assign n913 = n716 | n724;
  assign n914 = (n705 & n912) | (n705 & n913) | (n912 & n913);
  assign n521 = ~n911 & n914;
  assign n523 = x56 & x88;
  assign n524 = x56 | x88;
  assign n525 = ~n523 & n524;
  assign n915 = n509 | n516;
  assign n916 = (n516 & n518) | (n516 & n915) | (n518 & n915);
  assign n729 = n525 & n916;
  assign n727 = n516 | n518;
  assign n730 = n525 & n727;
  assign n917 = (n717 & n729) | (n717 & n730) | (n729 & n730);
  assign n918 = (n716 & n729) | (n716 & n730) | (n729 & n730);
  assign n919 = (n705 & n917) | (n705 & n918) | (n917 & n918);
  assign n732 = n525 | n916;
  assign n733 = n525 | n727;
  assign n920 = (n717 & n732) | (n717 & n733) | (n732 & n733);
  assign n921 = (n716 & n732) | (n716 & n733) | (n732 & n733);
  assign n922 = (n705 & n920) | (n705 & n921) | (n920 & n921);
  assign n528 = ~n919 & n922;
  assign n923 = n523 | n525;
  assign n924 = (n523 & n916) | (n523 & n923) | (n916 & n923);
  assign n925 = (n523 & n727) | (n523 & n923) | (n727 & n923);
  assign n926 = (n717 & n924) | (n717 & n925) | (n924 & n925);
  assign n927 = (n716 & n924) | (n716 & n925) | (n924 & n925);
  assign n928 = (n705 & n926) | (n705 & n927) | (n926 & n927);
  assign n530 = x57 & x89;
  assign n531 = x57 | x89;
  assign n532 = ~n530 & n531;
  assign n533 = n928 & n532;
  assign n534 = n928 | n532;
  assign n535 = ~n533 & n534;
  assign n537 = x58 & x90;
  assign n538 = x58 | x90;
  assign n539 = ~n537 & n538;
  assign n738 = n530 | n532;
  assign n740 = n539 & n738;
  assign n741 = n530 & n539;
  assign n742 = (n928 & n740) | (n928 & n741) | (n740 & n741);
  assign n743 = n539 | n738;
  assign n744 = n530 | n539;
  assign n745 = (n928 & n743) | (n928 & n744) | (n743 & n744);
  assign n542 = ~n742 & n745;
  assign n544 = x59 & x91;
  assign n545 = x59 | x91;
  assign n546 = ~n544 & n545;
  assign n929 = n537 | n539;
  assign n930 = (n537 & n738) | (n537 & n929) | (n738 & n929);
  assign n749 = n546 & n930;
  assign n931 = n530 | n537;
  assign n932 = (n537 & n539) | (n537 & n931) | (n539 & n931);
  assign n750 = n546 & n932;
  assign n751 = (n928 & n749) | (n928 & n750) | (n749 & n750);
  assign n752 = n546 | n930;
  assign n753 = n546 | n932;
  assign n754 = (n928 & n752) | (n928 & n753) | (n752 & n753);
  assign n549 = ~n751 & n754;
  assign n551 = x60 & x92;
  assign n552 = x60 | x92;
  assign n553 = ~n551 & n552;
  assign n933 = n544 | n546;
  assign n1658 = n553 & n933;
  assign n1659 = n544 & n553;
  assign n1660 = (n930 & n1658) | (n930 & n1659) | (n1658 & n1659);
  assign n935 = (n544 & n932) | (n544 & n933) | (n932 & n933);
  assign n937 = n553 & n935;
  assign n938 = (n928 & n1660) | (n928 & n937) | (n1660 & n937);
  assign n1661 = n553 | n933;
  assign n1662 = n544 | n553;
  assign n1663 = (n930 & n1661) | (n930 & n1662) | (n1661 & n1662);
  assign n940 = n553 | n935;
  assign n941 = (n928 & n1663) | (n928 & n940) | (n1663 & n940);
  assign n556 = ~n938 & n941;
  assign n558 = x61 & x93;
  assign n559 = x61 | x93;
  assign n560 = ~n558 & n559;
  assign n758 = n551 | n553;
  assign n760 = n560 & n758;
  assign n761 = n551 & n560;
  assign n934 = (n544 & n930) | (n544 & n933) | (n930 & n933);
  assign n942 = (n760 & n761) | (n760 & n934) | (n761 & n934);
  assign n943 = (n760 & n761) | (n760 & n935) | (n761 & n935);
  assign n944 = (n928 & n942) | (n928 & n943) | (n942 & n943);
  assign n763 = n560 | n758;
  assign n764 = n551 | n560;
  assign n945 = (n763 & n764) | (n763 & n934) | (n764 & n934);
  assign n946 = (n763 & n764) | (n763 & n935) | (n764 & n935);
  assign n947 = (n928 & n945) | (n928 & n946) | (n945 & n946);
  assign n563 = ~n944 & n947;
  assign n565 = x62 & x94;
  assign n566 = x62 | x94;
  assign n567 = ~n565 & n566;
  assign n948 = n558 | n560;
  assign n949 = (n558 & n758) | (n558 & n948) | (n758 & n948);
  assign n769 = n567 & n949;
  assign n950 = n551 | n558;
  assign n951 = (n558 & n560) | (n558 & n950) | (n560 & n950);
  assign n770 = n567 & n951;
  assign n952 = (n769 & n770) | (n769 & n934) | (n770 & n934);
  assign n953 = (n769 & n770) | (n769 & n935) | (n770 & n935);
  assign n954 = (n928 & n952) | (n928 & n953) | (n952 & n953);
  assign n772 = n567 | n949;
  assign n773 = n567 | n951;
  assign n955 = (n772 & n773) | (n772 & n934) | (n773 & n934);
  assign n956 = (n772 & n773) | (n772 & n935) | (n773 & n935);
  assign n957 = (n928 & n955) | (n928 & n956) | (n955 & n956);
  assign n570 = ~n954 & n957;
  assign n572 = x63 & x95;
  assign n573 = x63 | x95;
  assign n574 = ~n572 & n573;
  assign n958 = n565 | n567;
  assign n963 = (n565 & n951) | (n565 & n958) | (n951 & n958);
  assign n779 = n574 & n963;
  assign n960 = n574 & n958;
  assign n961 = n565 & n574;
  assign n962 = (n949 & n960) | (n949 & n961) | (n960 & n961);
  assign n964 = (n779 & n934) | (n779 & n962) | (n934 & n962);
  assign n965 = (n779 & n935) | (n779 & n962) | (n935 & n962);
  assign n966 = (n928 & n964) | (n928 & n965) | (n964 & n965);
  assign n782 = n574 | n963;
  assign n967 = n574 | n958;
  assign n968 = n565 | n574;
  assign n969 = (n949 & n967) | (n949 & n968) | (n967 & n968);
  assign n970 = (n782 & n934) | (n782 & n969) | (n934 & n969);
  assign n971 = (n782 & n935) | (n782 & n969) | (n935 & n969);
  assign n972 = (n928 & n970) | (n928 & n971) | (n970 & n971);
  assign n577 = ~n966 & n972;
  assign n579 = x64 & x96;
  assign n580 = x64 | x96;
  assign n581 = ~n579 & n580;
  assign n784 = n572 & n581;
  assign n785 = (n581 & n966) | (n581 & n784) | (n966 & n784);
  assign n786 = n572 | n581;
  assign n787 = n966 | n786;
  assign n584 = ~n785 & n787;
  assign n586 = x65 & x97;
  assign n587 = x65 | x97;
  assign n588 = ~n586 & n587;
  assign n973 = n572 | n579;
  assign n974 = (n579 & n581) | (n579 & n973) | (n581 & n973);
  assign n791 = n588 & n974;
  assign n789 = n579 | n581;
  assign n792 = n588 & n789;
  assign n793 = (n966 & n791) | (n966 & n792) | (n791 & n792);
  assign n794 = n588 | n974;
  assign n795 = n588 | n789;
  assign n796 = (n966 & n794) | (n966 & n795) | (n794 & n795);
  assign n591 = ~n793 & n796;
  assign n593 = x66 & x98;
  assign n594 = x66 | x98;
  assign n595 = ~n593 & n594;
  assign n975 = n586 | n588;
  assign n976 = (n586 & n974) | (n586 & n975) | (n974 & n975);
  assign n800 = n595 & n976;
  assign n977 = (n586 & n789) | (n586 & n975) | (n789 & n975);
  assign n801 = n595 & n977;
  assign n802 = (n966 & n800) | (n966 & n801) | (n800 & n801);
  assign n803 = n595 | n976;
  assign n804 = n595 | n977;
  assign n805 = (n966 & n803) | (n966 & n804) | (n803 & n804);
  assign n598 = ~n802 & n805;
  assign n600 = x67 & x99;
  assign n601 = x67 | x99;
  assign n602 = ~n600 & n601;
  assign n978 = n593 | n595;
  assign n980 = n602 & n978;
  assign n981 = n593 & n602;
  assign n982 = (n976 & n980) | (n976 & n981) | (n980 & n981);
  assign n984 = (n977 & n980) | (n977 & n981) | (n980 & n981);
  assign n811 = (n966 & n982) | (n966 & n984) | (n982 & n984);
  assign n985 = n602 | n978;
  assign n986 = n593 | n602;
  assign n987 = (n976 & n985) | (n976 & n986) | (n985 & n986);
  assign n988 = (n977 & n985) | (n977 & n986) | (n985 & n986);
  assign n814 = (n966 & n987) | (n966 & n988) | (n987 & n988);
  assign n605 = ~n811 & n814;
  assign n607 = x68 & x100;
  assign n608 = x68 | x100;
  assign n609 = ~n607 & n608;
  assign n815 = n600 & n609;
  assign n989 = (n609 & n815) | (n609 & n984) | (n815 & n984);
  assign n990 = (n609 & n815) | (n609 & n982) | (n815 & n982);
  assign n991 = (n966 & n989) | (n966 & n990) | (n989 & n990);
  assign n817 = n600 | n609;
  assign n992 = n817 | n984;
  assign n993 = n817 | n982;
  assign n994 = (n966 & n992) | (n966 & n993) | (n992 & n993);
  assign n612 = ~n991 & n994;
  assign n614 = x69 & x101;
  assign n615 = x69 | x101;
  assign n616 = ~n614 & n615;
  assign n995 = n600 | n607;
  assign n996 = (n607 & n609) | (n607 & n995) | (n609 & n995);
  assign n822 = n616 & n996;
  assign n820 = n607 | n609;
  assign n823 = n616 & n820;
  assign n997 = (n822 & n823) | (n822 & n984) | (n823 & n984);
  assign n998 = (n822 & n823) | (n822 & n982) | (n823 & n982);
  assign n999 = (n966 & n997) | (n966 & n998) | (n997 & n998);
  assign n825 = n616 | n996;
  assign n826 = n616 | n820;
  assign n1000 = (n825 & n826) | (n825 & n984) | (n826 & n984);
  assign n1001 = (n825 & n826) | (n825 & n982) | (n826 & n982);
  assign n1002 = (n966 & n1000) | (n966 & n1001) | (n1000 & n1001);
  assign n619 = ~n999 & n1002;
  assign n621 = x70 & x102;
  assign n622 = x70 | x102;
  assign n623 = ~n621 & n622;
  assign n1003 = n614 | n616;
  assign n1004 = (n614 & n996) | (n614 & n1003) | (n996 & n1003);
  assign n831 = n623 & n1004;
  assign n1005 = (n614 & n820) | (n614 & n1003) | (n820 & n1003);
  assign n832 = n623 & n1005;
  assign n1006 = (n831 & n832) | (n831 & n984) | (n832 & n984);
  assign n1007 = (n831 & n832) | (n831 & n982) | (n832 & n982);
  assign n1008 = (n966 & n1006) | (n966 & n1007) | (n1006 & n1007);
  assign n834 = n623 | n1004;
  assign n835 = n623 | n1005;
  assign n1009 = (n834 & n835) | (n834 & n984) | (n835 & n984);
  assign n1010 = (n834 & n835) | (n834 & n982) | (n835 & n982);
  assign n1011 = (n966 & n1009) | (n966 & n1010) | (n1009 & n1010);
  assign n626 = ~n1008 & n1011;
  assign n628 = x71 & x103;
  assign n629 = x71 | x103;
  assign n630 = ~n628 & n629;
  assign n1012 = n621 | n623;
  assign n1014 = n630 & n1012;
  assign n1015 = n621 & n630;
  assign n1016 = (n1004 & n1014) | (n1004 & n1015) | (n1014 & n1015);
  assign n1018 = (n1005 & n1014) | (n1005 & n1015) | (n1014 & n1015);
  assign n1019 = (n984 & n1016) | (n984 & n1018) | (n1016 & n1018);
  assign n1020 = (n982 & n1016) | (n982 & n1018) | (n1016 & n1018);
  assign n1021 = (n966 & n1019) | (n966 & n1020) | (n1019 & n1020);
  assign n1022 = n630 | n1012;
  assign n1023 = n621 | n630;
  assign n1024 = (n1004 & n1022) | (n1004 & n1023) | (n1022 & n1023);
  assign n1025 = (n1005 & n1022) | (n1005 & n1023) | (n1022 & n1023);
  assign n1026 = (n984 & n1024) | (n984 & n1025) | (n1024 & n1025);
  assign n1027 = (n982 & n1024) | (n982 & n1025) | (n1024 & n1025);
  assign n1028 = (n966 & n1026) | (n966 & n1027) | (n1026 & n1027);
  assign n633 = ~n1021 & n1028;
  assign n846 = n628 | n1016;
  assign n847 = n628 | n1018;
  assign n1029 = (n846 & n847) | (n846 & n984) | (n847 & n984);
  assign n1030 = (n846 & n847) | (n846 & n982) | (n847 & n982);
  assign n1031 = (n966 & n1029) | (n966 & n1030) | (n1029 & n1030);
  assign n635 = x72 & x104;
  assign n636 = x72 | x104;
  assign n637 = ~n635 & n636;
  assign n638 = n1031 & n637;
  assign n639 = n1031 | n637;
  assign n640 = ~n638 & n639;
  assign n642 = x73 & x105;
  assign n643 = x73 | x105;
  assign n644 = ~n642 & n643;
  assign n849 = n635 | n637;
  assign n851 = n644 & n849;
  assign n852 = n635 & n644;
  assign n853 = (n1031 & n851) | (n1031 & n852) | (n851 & n852);
  assign n854 = n644 | n849;
  assign n855 = n635 | n644;
  assign n856 = (n1031 & n854) | (n1031 & n855) | (n854 & n855);
  assign n647 = ~n853 & n856;
  assign n649 = x74 & x106;
  assign n650 = x74 | x106;
  assign n651 = ~n649 & n650;
  assign n1032 = n642 | n644;
  assign n1033 = (n642 & n849) | (n642 & n1032) | (n849 & n1032);
  assign n860 = n651 & n1033;
  assign n1034 = n635 | n642;
  assign n1035 = (n642 & n644) | (n642 & n1034) | (n644 & n1034);
  assign n861 = n651 & n1035;
  assign n862 = (n1031 & n860) | (n1031 & n861) | (n860 & n861);
  assign n863 = n651 | n1033;
  assign n864 = n651 | n1035;
  assign n865 = (n1031 & n863) | (n1031 & n864) | (n863 & n864);
  assign n654 = ~n862 & n865;
  assign n656 = x75 & x107;
  assign n657 = x75 | x107;
  assign n658 = ~n656 & n657;
  assign n1036 = n649 | n651;
  assign n1038 = n658 & n1036;
  assign n1039 = n649 & n658;
  assign n1040 = (n1033 & n1038) | (n1033 & n1039) | (n1038 & n1039);
  assign n1041 = (n649 & n1035) | (n649 & n1036) | (n1035 & n1036);
  assign n870 = n658 & n1041;
  assign n871 = (n1031 & n1040) | (n1031 & n870) | (n1040 & n870);
  assign n1042 = n658 | n1036;
  assign n1043 = n649 | n658;
  assign n1044 = (n1033 & n1042) | (n1033 & n1043) | (n1042 & n1043);
  assign n873 = n658 | n1041;
  assign n874 = (n1031 & n1044) | (n1031 & n873) | (n1044 & n873);
  assign n661 = ~n871 & n874;
  assign n663 = x76 & x108;
  assign n664 = x76 | x108;
  assign n665 = ~n663 & n664;
  assign n1045 = n656 & n665;
  assign n1046 = (n665 & n1040) | (n665 & n1045) | (n1040 & n1045);
  assign n1047 = n656 | n658;
  assign n1049 = n665 & n1047;
  assign n1050 = (n1041 & n1045) | (n1041 & n1049) | (n1045 & n1049);
  assign n880 = (n1031 & n1046) | (n1031 & n1050) | (n1046 & n1050);
  assign n1051 = n656 | n665;
  assign n1052 = n1040 | n1051;
  assign n1053 = n665 | n1047;
  assign n1054 = (n1041 & n1051) | (n1041 & n1053) | (n1051 & n1053);
  assign n883 = (n1031 & n1052) | (n1031 & n1054) | (n1052 & n1054);
  assign n668 = ~n880 & n883;
  assign n670 = x77 & x109;
  assign n671 = x77 | x109;
  assign n672 = ~n670 & n671;
  assign n1664 = n663 & n672;
  assign n1665 = (n672 & n1050) | (n672 & n1664) | (n1050 & n1664);
  assign n1056 = n663 | n665;
  assign n1668 = n672 & n1056;
  assign n1666 = n656 | n663;
  assign n1667 = (n663 & n665) | (n663 & n1666) | (n665 & n1666);
  assign n1669 = n672 & n1667;
  assign n1670 = (n1040 & n1668) | (n1040 & n1669) | (n1668 & n1669);
  assign n1060 = (n1031 & n1665) | (n1031 & n1670) | (n1665 & n1670);
  assign n1671 = n663 | n672;
  assign n1672 = n1050 | n1671;
  assign n1673 = n672 | n1056;
  assign n1674 = n672 | n1667;
  assign n1675 = (n1040 & n1673) | (n1040 & n1674) | (n1673 & n1674);
  assign n1063 = (n1031 & n1672) | (n1031 & n1675) | (n1672 & n1675);
  assign n675 = ~n1060 & n1063;
  assign n677 = x78 & x110;
  assign n678 = x78 | x110;
  assign n679 = ~n677 & n678;
  assign n887 = n670 | n672;
  assign n889 = n679 & n887;
  assign n890 = n670 & n679;
  assign n1676 = (n663 & n889) | (n663 & n890) | (n889 & n890);
  assign n1677 = n889 | n890;
  assign n1678 = (n1050 & n1676) | (n1050 & n1677) | (n1676 & n1677);
  assign n1679 = (n889 & n890) | (n889 & n1056) | (n890 & n1056);
  assign n1680 = (n889 & n890) | (n889 & n1667) | (n890 & n1667);
  assign n1681 = (n1040 & n1679) | (n1040 & n1680) | (n1679 & n1680);
  assign n1066 = (n1031 & n1678) | (n1031 & n1681) | (n1678 & n1681);
  assign n892 = n679 | n887;
  assign n893 = n670 | n679;
  assign n1682 = (n663 & n892) | (n663 & n893) | (n892 & n893);
  assign n1683 = n892 | n893;
  assign n1684 = (n1050 & n1682) | (n1050 & n1683) | (n1682 & n1683);
  assign n1685 = (n892 & n893) | (n892 & n1056) | (n893 & n1056);
  assign n1686 = (n892 & n893) | (n892 & n1667) | (n893 & n1667);
  assign n1687 = (n1040 & n1685) | (n1040 & n1686) | (n1685 & n1686);
  assign n1069 = (n1031 & n1684) | (n1031 & n1687) | (n1684 & n1687);
  assign n682 = ~n1066 & n1069;
  assign n885 = n663 | n1050;
  assign n684 = x79 & x111;
  assign n685 = x79 | x111;
  assign n686 = ~n684 & n685;
  assign n1070 = n677 | n679;
  assign n1071 = (n677 & n887) | (n677 & n1070) | (n887 & n1070);
  assign n898 = n686 & n1071;
  assign n1072 = n670 | n677;
  assign n1073 = (n677 & n679) | (n677 & n1072) | (n679 & n1072);
  assign n899 = n686 & n1073;
  assign n1074 = (n885 & n898) | (n885 & n899) | (n898 & n899);
  assign n1057 = (n1040 & n1667) | (n1040 & n1056) | (n1667 & n1056);
  assign n1075 = (n898 & n899) | (n898 & n1057) | (n899 & n1057);
  assign n1076 = (n1031 & n1074) | (n1031 & n1075) | (n1074 & n1075);
  assign n901 = n686 | n1071;
  assign n902 = n686 | n1073;
  assign n1077 = (n885 & n901) | (n885 & n902) | (n901 & n902);
  assign n1078 = (n901 & n902) | (n901 & n1057) | (n902 & n1057);
  assign n1079 = (n1031 & n1077) | (n1031 & n1078) | (n1077 & n1078);
  assign n689 = ~n1076 & n1079;
  assign n1080 = n684 | n686;
  assign n1081 = (n684 & n1071) | (n684 & n1080) | (n1071 & n1080);
  assign n1082 = (n684 & n1073) | (n684 & n1080) | (n1073 & n1080);
  assign n1083 = (n885 & n1081) | (n885 & n1082) | (n1081 & n1082);
  assign n1084 = (n1057 & n1081) | (n1057 & n1082) | (n1081 & n1082);
  assign n1085 = (n1031 & n1083) | (n1031 & n1084) | (n1083 & n1084);
  assign n1214 = x112 & x176;
  assign n1215 = x112 | x176;
  assign n1216 = ~n1214 & n1215;
  assign n1217 = x113 & x177;
  assign n1218 = x113 | x177;
  assign n1219 = ~n1217 & n1218;
  assign n1220 = n1214 & n1219;
  assign n1221 = n1214 | n1219;
  assign n1222 = ~n1220 & n1221;
  assign n1688 = n1214 | n1217;
  assign n1689 = (n1217 & n1219) | (n1217 & n1688) | (n1219 & n1688);
  assign n1224 = x114 & x178;
  assign n1225 = x114 | x178;
  assign n1226 = ~n1224 & n1225;
  assign n1227 = n1689 & n1226;
  assign n1228 = n1689 | n1226;
  assign n1229 = ~n1227 & n1228;
  assign n1690 = n1224 | n1226;
  assign n1691 = (n1224 & n1689) | (n1224 & n1690) | (n1689 & n1690);
  assign n1231 = x115 & x179;
  assign n1232 = x115 | x179;
  assign n1233 = ~n1231 & n1232;
  assign n1234 = n1691 & n1233;
  assign n1235 = n1691 | n1233;
  assign n1236 = ~n1234 & n1235;
  assign n1238 = x116 & x180;
  assign n1239 = x116 | x180;
  assign n1240 = ~n1238 & n1239;
  assign n1692 = n1231 | n1233;
  assign n1694 = n1240 & n1692;
  assign n1695 = n1231 & n1240;
  assign n1696 = (n1691 & n1694) | (n1691 & n1695) | (n1694 & n1695);
  assign n1697 = n1240 | n1692;
  assign n1698 = n1231 | n1240;
  assign n1699 = (n1691 & n1697) | (n1691 & n1698) | (n1697 & n1698);
  assign n1243 = ~n1696 & n1699;
  assign n1245 = x117 & x181;
  assign n1246 = x117 | x181;
  assign n1247 = ~n1245 & n1246;
  assign n1700 = n1238 & n1247;
  assign n1701 = (n1247 & n1696) | (n1247 & n1700) | (n1696 & n1700);
  assign n1702 = n1238 | n1247;
  assign n1703 = n1696 | n1702;
  assign n1250 = ~n1701 & n1703;
  assign n1252 = x118 & x182;
  assign n1253 = x118 | x182;
  assign n1254 = ~n1252 & n1253;
  assign n2157 = n1238 | n1245;
  assign n2158 = (n1245 & n1247) | (n1245 & n2157) | (n1247 & n2157);
  assign n1707 = n1254 & n2158;
  assign n1705 = n1245 | n1247;
  assign n1708 = n1254 & n1705;
  assign n1709 = (n1696 & n1707) | (n1696 & n1708) | (n1707 & n1708);
  assign n1710 = n1254 | n2158;
  assign n1711 = n1254 | n1705;
  assign n1712 = (n1696 & n1710) | (n1696 & n1711) | (n1710 & n1711);
  assign n1257 = ~n1709 & n1712;
  assign n1259 = x119 & x183;
  assign n1260 = x119 | x183;
  assign n1261 = ~n1259 & n1260;
  assign n1713 = n1252 & n1261;
  assign n2159 = (n1261 & n1708) | (n1261 & n1713) | (n1708 & n1713);
  assign n2160 = (n1261 & n1707) | (n1261 & n1713) | (n1707 & n1713);
  assign n2161 = (n1696 & n2159) | (n1696 & n2160) | (n2159 & n2160);
  assign n1715 = n1252 | n1261;
  assign n2162 = n1708 | n1715;
  assign n2163 = n1707 | n1715;
  assign n2164 = (n1696 & n2162) | (n1696 & n2163) | (n2162 & n2163);
  assign n1264 = ~n2161 & n2164;
  assign n1266 = x120 & x184;
  assign n1267 = x120 | x184;
  assign n1268 = ~n1266 & n1267;
  assign n2165 = n1252 | n1259;
  assign n2166 = (n1259 & n1261) | (n1259 & n2165) | (n1261 & n2165);
  assign n1720 = n1268 & n2166;
  assign n1718 = n1259 | n1261;
  assign n1721 = n1268 & n1718;
  assign n2167 = (n1708 & n1720) | (n1708 & n1721) | (n1720 & n1721);
  assign n2168 = (n1707 & n1720) | (n1707 & n1721) | (n1720 & n1721);
  assign n2169 = (n1696 & n2167) | (n1696 & n2168) | (n2167 & n2168);
  assign n1723 = n1268 | n2166;
  assign n1724 = n1268 | n1718;
  assign n2170 = (n1708 & n1723) | (n1708 & n1724) | (n1723 & n1724);
  assign n2171 = (n1707 & n1723) | (n1707 & n1724) | (n1723 & n1724);
  assign n2172 = (n1696 & n2170) | (n1696 & n2171) | (n2170 & n2171);
  assign n1271 = ~n2169 & n2172;
  assign n2173 = n1266 | n1268;
  assign n2174 = (n1266 & n2166) | (n1266 & n2173) | (n2166 & n2173);
  assign n2175 = (n1266 & n1718) | (n1266 & n2173) | (n1718 & n2173);
  assign n2176 = (n1708 & n2174) | (n1708 & n2175) | (n2174 & n2175);
  assign n2177 = (n1707 & n2174) | (n1707 & n2175) | (n2174 & n2175);
  assign n2178 = (n1696 & n2176) | (n1696 & n2177) | (n2176 & n2177);
  assign n1273 = x121 & x185;
  assign n1274 = x121 | x185;
  assign n1275 = ~n1273 & n1274;
  assign n1276 = n2178 & n1275;
  assign n1277 = n2178 | n1275;
  assign n1278 = ~n1276 & n1277;
  assign n1280 = x122 & x186;
  assign n1281 = x122 | x186;
  assign n1282 = ~n1280 & n1281;
  assign n1729 = n1273 | n1275;
  assign n1731 = n1282 & n1729;
  assign n1732 = n1273 & n1282;
  assign n1733 = (n2178 & n1731) | (n2178 & n1732) | (n1731 & n1732);
  assign n1734 = n1282 | n1729;
  assign n1735 = n1273 | n1282;
  assign n1736 = (n2178 & n1734) | (n2178 & n1735) | (n1734 & n1735);
  assign n1285 = ~n1733 & n1736;
  assign n1287 = x123 & x187;
  assign n1288 = x123 | x187;
  assign n1289 = ~n1287 & n1288;
  assign n2179 = n1280 | n1282;
  assign n2180 = (n1280 & n1729) | (n1280 & n2179) | (n1729 & n2179);
  assign n1740 = n1289 & n2180;
  assign n2181 = n1273 | n1280;
  assign n2182 = (n1280 & n1282) | (n1280 & n2181) | (n1282 & n2181);
  assign n1741 = n1289 & n2182;
  assign n1742 = (n2178 & n1740) | (n2178 & n1741) | (n1740 & n1741);
  assign n1743 = n1289 | n2180;
  assign n1744 = n1289 | n2182;
  assign n1745 = (n2178 & n1743) | (n2178 & n1744) | (n1743 & n1744);
  assign n1292 = ~n1742 & n1745;
  assign n1294 = x124 & x188;
  assign n1295 = x124 | x188;
  assign n1296 = ~n1294 & n1295;
  assign n2183 = n1287 | n1289;
  assign n2696 = n1296 & n2183;
  assign n2697 = n1287 & n1296;
  assign n2698 = (n2180 & n2696) | (n2180 & n2697) | (n2696 & n2697);
  assign n2185 = (n1287 & n2182) | (n1287 & n2183) | (n2182 & n2183);
  assign n2187 = n1296 & n2185;
  assign n2188 = (n2178 & n2698) | (n2178 & n2187) | (n2698 & n2187);
  assign n2699 = n1296 | n2183;
  assign n2700 = n1287 | n1296;
  assign n2701 = (n2180 & n2699) | (n2180 & n2700) | (n2699 & n2700);
  assign n2190 = n1296 | n2185;
  assign n2191 = (n2178 & n2701) | (n2178 & n2190) | (n2701 & n2190);
  assign n1299 = ~n2188 & n2191;
  assign n1301 = x125 & x189;
  assign n1302 = x125 | x189;
  assign n1303 = ~n1301 & n1302;
  assign n1749 = n1294 | n1296;
  assign n1751 = n1303 & n1749;
  assign n1752 = n1294 & n1303;
  assign n2184 = (n1287 & n2180) | (n1287 & n2183) | (n2180 & n2183);
  assign n2192 = (n1751 & n1752) | (n1751 & n2184) | (n1752 & n2184);
  assign n2193 = (n1751 & n1752) | (n1751 & n2185) | (n1752 & n2185);
  assign n2194 = (n2178 & n2192) | (n2178 & n2193) | (n2192 & n2193);
  assign n1754 = n1303 | n1749;
  assign n1755 = n1294 | n1303;
  assign n2195 = (n1754 & n1755) | (n1754 & n2184) | (n1755 & n2184);
  assign n2196 = (n1754 & n1755) | (n1754 & n2185) | (n1755 & n2185);
  assign n2197 = (n2178 & n2195) | (n2178 & n2196) | (n2195 & n2196);
  assign n1306 = ~n2194 & n2197;
  assign n1308 = x126 & x190;
  assign n1309 = x126 | x190;
  assign n1310 = ~n1308 & n1309;
  assign n2198 = n1301 | n1303;
  assign n2199 = (n1301 & n1749) | (n1301 & n2198) | (n1749 & n2198);
  assign n1760 = n1310 & n2199;
  assign n2200 = n1294 | n1301;
  assign n2201 = (n1301 & n1303) | (n1301 & n2200) | (n1303 & n2200);
  assign n1761 = n1310 & n2201;
  assign n2202 = (n1760 & n1761) | (n1760 & n2184) | (n1761 & n2184);
  assign n2203 = (n1760 & n1761) | (n1760 & n2185) | (n1761 & n2185);
  assign n2204 = (n2178 & n2202) | (n2178 & n2203) | (n2202 & n2203);
  assign n1763 = n1310 | n2199;
  assign n1764 = n1310 | n2201;
  assign n2205 = (n1763 & n1764) | (n1763 & n2184) | (n1764 & n2184);
  assign n2206 = (n1763 & n1764) | (n1763 & n2185) | (n1764 & n2185);
  assign n2207 = (n2178 & n2205) | (n2178 & n2206) | (n2205 & n2206);
  assign n1313 = ~n2204 & n2207;
  assign n1315 = x127 & x191;
  assign n1316 = x127 | x191;
  assign n1317 = ~n1315 & n1316;
  assign n2208 = n1308 | n1310;
  assign n2213 = (n1308 & n2201) | (n1308 & n2208) | (n2201 & n2208);
  assign n1770 = n1317 & n2213;
  assign n2210 = n1317 & n2208;
  assign n2211 = n1308 & n1317;
  assign n2212 = (n2199 & n2210) | (n2199 & n2211) | (n2210 & n2211);
  assign n2214 = (n1770 & n2184) | (n1770 & n2212) | (n2184 & n2212);
  assign n2215 = (n1770 & n2185) | (n1770 & n2212) | (n2185 & n2212);
  assign n2216 = (n2178 & n2214) | (n2178 & n2215) | (n2214 & n2215);
  assign n1773 = n1317 | n2213;
  assign n2217 = n1317 | n2208;
  assign n2218 = n1308 | n1317;
  assign n2219 = (n2199 & n2217) | (n2199 & n2218) | (n2217 & n2218);
  assign n2220 = (n1773 & n2184) | (n1773 & n2219) | (n2184 & n2219);
  assign n2221 = (n1773 & n2185) | (n1773 & n2219) | (n2185 & n2219);
  assign n2222 = (n2178 & n2220) | (n2178 & n2221) | (n2220 & n2221);
  assign n1320 = ~n2216 & n2222;
  assign n1322 = x128 & x192;
  assign n1323 = x128 | x192;
  assign n1324 = ~n1322 & n1323;
  assign n1775 = n1315 & n1324;
  assign n1776 = (n1324 & n2216) | (n1324 & n1775) | (n2216 & n1775);
  assign n1777 = n1315 | n1324;
  assign n1778 = n2216 | n1777;
  assign n1327 = ~n1776 & n1778;
  assign n1329 = x129 & x193;
  assign n1330 = x129 | x193;
  assign n1331 = ~n1329 & n1330;
  assign n2223 = n1315 | n1322;
  assign n2224 = (n1322 & n1324) | (n1322 & n2223) | (n1324 & n2223);
  assign n1782 = n1331 & n2224;
  assign n1780 = n1322 | n1324;
  assign n1783 = n1331 & n1780;
  assign n1784 = (n2216 & n1782) | (n2216 & n1783) | (n1782 & n1783);
  assign n1785 = n1331 | n2224;
  assign n1786 = n1331 | n1780;
  assign n1787 = (n2216 & n1785) | (n2216 & n1786) | (n1785 & n1786);
  assign n1334 = ~n1784 & n1787;
  assign n1336 = x130 & x194;
  assign n1337 = x130 | x194;
  assign n1338 = ~n1336 & n1337;
  assign n2225 = n1329 | n1331;
  assign n2226 = (n1329 & n2224) | (n1329 & n2225) | (n2224 & n2225);
  assign n1791 = n1338 & n2226;
  assign n2227 = (n1329 & n1780) | (n1329 & n2225) | (n1780 & n2225);
  assign n1792 = n1338 & n2227;
  assign n1793 = (n2216 & n1791) | (n2216 & n1792) | (n1791 & n1792);
  assign n1794 = n1338 | n2226;
  assign n1795 = n1338 | n2227;
  assign n1796 = (n2216 & n1794) | (n2216 & n1795) | (n1794 & n1795);
  assign n1341 = ~n1793 & n1796;
  assign n1343 = x131 & x195;
  assign n1344 = x131 | x195;
  assign n1345 = ~n1343 & n1344;
  assign n2228 = n1336 | n1338;
  assign n2230 = n1345 & n2228;
  assign n2231 = n1336 & n1345;
  assign n2232 = (n2226 & n2230) | (n2226 & n2231) | (n2230 & n2231);
  assign n2234 = (n2227 & n2230) | (n2227 & n2231) | (n2230 & n2231);
  assign n1802 = (n2216 & n2232) | (n2216 & n2234) | (n2232 & n2234);
  assign n2235 = n1345 | n2228;
  assign n2236 = n1336 | n1345;
  assign n2237 = (n2226 & n2235) | (n2226 & n2236) | (n2235 & n2236);
  assign n2238 = (n2227 & n2235) | (n2227 & n2236) | (n2235 & n2236);
  assign n1805 = (n2216 & n2237) | (n2216 & n2238) | (n2237 & n2238);
  assign n1348 = ~n1802 & n1805;
  assign n1350 = x132 & x196;
  assign n1351 = x132 | x196;
  assign n1352 = ~n1350 & n1351;
  assign n1806 = n1343 & n1352;
  assign n2239 = (n1352 & n1806) | (n1352 & n2234) | (n1806 & n2234);
  assign n2240 = (n1352 & n1806) | (n1352 & n2232) | (n1806 & n2232);
  assign n2241 = (n2216 & n2239) | (n2216 & n2240) | (n2239 & n2240);
  assign n1808 = n1343 | n1352;
  assign n2242 = n1808 | n2234;
  assign n2243 = n1808 | n2232;
  assign n2244 = (n2216 & n2242) | (n2216 & n2243) | (n2242 & n2243);
  assign n1355 = ~n2241 & n2244;
  assign n1357 = x133 & x197;
  assign n1358 = x133 | x197;
  assign n1359 = ~n1357 & n1358;
  assign n2245 = n1343 | n1350;
  assign n2246 = (n1350 & n1352) | (n1350 & n2245) | (n1352 & n2245);
  assign n1813 = n1359 & n2246;
  assign n1811 = n1350 | n1352;
  assign n1814 = n1359 & n1811;
  assign n2247 = (n1813 & n1814) | (n1813 & n2234) | (n1814 & n2234);
  assign n2248 = (n1813 & n1814) | (n1813 & n2232) | (n1814 & n2232);
  assign n2249 = (n2216 & n2247) | (n2216 & n2248) | (n2247 & n2248);
  assign n1816 = n1359 | n2246;
  assign n1817 = n1359 | n1811;
  assign n2250 = (n1816 & n1817) | (n1816 & n2234) | (n1817 & n2234);
  assign n2251 = (n1816 & n1817) | (n1816 & n2232) | (n1817 & n2232);
  assign n2252 = (n2216 & n2250) | (n2216 & n2251) | (n2250 & n2251);
  assign n1362 = ~n2249 & n2252;
  assign n1364 = x134 & x198;
  assign n1365 = x134 | x198;
  assign n1366 = ~n1364 & n1365;
  assign n2253 = n1357 | n1359;
  assign n2254 = (n1357 & n2246) | (n1357 & n2253) | (n2246 & n2253);
  assign n1822 = n1366 & n2254;
  assign n2255 = (n1357 & n1811) | (n1357 & n2253) | (n1811 & n2253);
  assign n1823 = n1366 & n2255;
  assign n2256 = (n1822 & n1823) | (n1822 & n2234) | (n1823 & n2234);
  assign n2257 = (n1822 & n1823) | (n1822 & n2232) | (n1823 & n2232);
  assign n2258 = (n2216 & n2256) | (n2216 & n2257) | (n2256 & n2257);
  assign n1825 = n1366 | n2254;
  assign n1826 = n1366 | n2255;
  assign n2259 = (n1825 & n1826) | (n1825 & n2234) | (n1826 & n2234);
  assign n2260 = (n1825 & n1826) | (n1825 & n2232) | (n1826 & n2232);
  assign n2261 = (n2216 & n2259) | (n2216 & n2260) | (n2259 & n2260);
  assign n1369 = ~n2258 & n2261;
  assign n1371 = x135 & x199;
  assign n1372 = x135 | x199;
  assign n1373 = ~n1371 & n1372;
  assign n2262 = n1364 | n1366;
  assign n2264 = n1373 & n2262;
  assign n2265 = n1364 & n1373;
  assign n2266 = (n2254 & n2264) | (n2254 & n2265) | (n2264 & n2265);
  assign n2268 = (n2255 & n2264) | (n2255 & n2265) | (n2264 & n2265);
  assign n2269 = (n2234 & n2266) | (n2234 & n2268) | (n2266 & n2268);
  assign n2270 = (n2232 & n2266) | (n2232 & n2268) | (n2266 & n2268);
  assign n2271 = (n2216 & n2269) | (n2216 & n2270) | (n2269 & n2270);
  assign n2272 = n1373 | n2262;
  assign n2273 = n1364 | n1373;
  assign n2274 = (n2254 & n2272) | (n2254 & n2273) | (n2272 & n2273);
  assign n2275 = (n2255 & n2272) | (n2255 & n2273) | (n2272 & n2273);
  assign n2276 = (n2234 & n2274) | (n2234 & n2275) | (n2274 & n2275);
  assign n2277 = (n2232 & n2274) | (n2232 & n2275) | (n2274 & n2275);
  assign n2278 = (n2216 & n2276) | (n2216 & n2277) | (n2276 & n2277);
  assign n1376 = ~n2271 & n2278;
  assign n1837 = n1371 | n2266;
  assign n1838 = n1371 | n2268;
  assign n2279 = (n1837 & n1838) | (n1837 & n2234) | (n1838 & n2234);
  assign n2280 = (n1837 & n1838) | (n1837 & n2232) | (n1838 & n2232);
  assign n2281 = (n2216 & n2279) | (n2216 & n2280) | (n2279 & n2280);
  assign n1378 = x136 & x200;
  assign n1379 = x136 | x200;
  assign n1380 = ~n1378 & n1379;
  assign n1381 = n2281 & n1380;
  assign n1382 = n2281 | n1380;
  assign n1383 = ~n1381 & n1382;
  assign n1385 = x137 & x201;
  assign n1386 = x137 | x201;
  assign n1387 = ~n1385 & n1386;
  assign n1840 = n1378 | n1380;
  assign n1842 = n1387 & n1840;
  assign n1843 = n1378 & n1387;
  assign n1844 = (n2281 & n1842) | (n2281 & n1843) | (n1842 & n1843);
  assign n1845 = n1387 | n1840;
  assign n1846 = n1378 | n1387;
  assign n1847 = (n2281 & n1845) | (n2281 & n1846) | (n1845 & n1846);
  assign n1390 = ~n1844 & n1847;
  assign n1392 = x138 & x202;
  assign n1393 = x138 | x202;
  assign n1394 = ~n1392 & n1393;
  assign n2282 = n1385 | n1387;
  assign n2283 = (n1385 & n1840) | (n1385 & n2282) | (n1840 & n2282);
  assign n1851 = n1394 & n2283;
  assign n2284 = n1378 | n1385;
  assign n2285 = (n1385 & n1387) | (n1385 & n2284) | (n1387 & n2284);
  assign n1852 = n1394 & n2285;
  assign n1853 = (n2281 & n1851) | (n2281 & n1852) | (n1851 & n1852);
  assign n1854 = n1394 | n2283;
  assign n1855 = n1394 | n2285;
  assign n1856 = (n2281 & n1854) | (n2281 & n1855) | (n1854 & n1855);
  assign n1397 = ~n1853 & n1856;
  assign n1399 = x139 & x203;
  assign n1400 = x139 | x203;
  assign n1401 = ~n1399 & n1400;
  assign n2286 = n1392 | n1394;
  assign n2288 = n1401 & n2286;
  assign n2289 = n1392 & n1401;
  assign n2290 = (n2283 & n2288) | (n2283 & n2289) | (n2288 & n2289);
  assign n2291 = (n1392 & n2285) | (n1392 & n2286) | (n2285 & n2286);
  assign n1861 = n1401 & n2291;
  assign n1862 = (n2281 & n2290) | (n2281 & n1861) | (n2290 & n1861);
  assign n2292 = n1401 | n2286;
  assign n2293 = n1392 | n1401;
  assign n2294 = (n2283 & n2292) | (n2283 & n2293) | (n2292 & n2293);
  assign n1864 = n1401 | n2291;
  assign n1865 = (n2281 & n2294) | (n2281 & n1864) | (n2294 & n1864);
  assign n1404 = ~n1862 & n1865;
  assign n1406 = x140 & x204;
  assign n1407 = x140 | x204;
  assign n1408 = ~n1406 & n1407;
  assign n2295 = n1399 & n1408;
  assign n2296 = (n1408 & n2290) | (n1408 & n2295) | (n2290 & n2295);
  assign n2297 = n1399 | n1401;
  assign n2299 = n1408 & n2297;
  assign n2300 = (n2291 & n2295) | (n2291 & n2299) | (n2295 & n2299);
  assign n1871 = (n2281 & n2296) | (n2281 & n2300) | (n2296 & n2300);
  assign n2301 = n1399 | n1408;
  assign n2302 = n2290 | n2301;
  assign n2303 = n1408 | n2297;
  assign n2304 = (n2291 & n2301) | (n2291 & n2303) | (n2301 & n2303);
  assign n1874 = (n2281 & n2302) | (n2281 & n2304) | (n2302 & n2304);
  assign n1411 = ~n1871 & n1874;
  assign n1413 = x141 & x205;
  assign n1414 = x141 | x205;
  assign n1415 = ~n1413 & n1414;
  assign n2702 = n1406 & n1415;
  assign n2703 = (n1415 & n2300) | (n1415 & n2702) | (n2300 & n2702);
  assign n2306 = n1406 | n1408;
  assign n2706 = n1415 & n2306;
  assign n2704 = n1399 | n1406;
  assign n2705 = (n1406 & n1408) | (n1406 & n2704) | (n1408 & n2704);
  assign n2707 = n1415 & n2705;
  assign n2708 = (n2290 & n2706) | (n2290 & n2707) | (n2706 & n2707);
  assign n2310 = (n2281 & n2703) | (n2281 & n2708) | (n2703 & n2708);
  assign n2709 = n1406 | n1415;
  assign n2710 = n2300 | n2709;
  assign n2711 = n1415 | n2306;
  assign n2712 = n1415 | n2705;
  assign n2713 = (n2290 & n2711) | (n2290 & n2712) | (n2711 & n2712);
  assign n2313 = (n2281 & n2710) | (n2281 & n2713) | (n2710 & n2713);
  assign n1418 = ~n2310 & n2313;
  assign n1420 = x142 & x206;
  assign n1421 = x142 | x206;
  assign n1422 = ~n1420 & n1421;
  assign n1878 = n1413 | n1415;
  assign n1880 = n1422 & n1878;
  assign n1881 = n1413 & n1422;
  assign n2714 = (n1406 & n1880) | (n1406 & n1881) | (n1880 & n1881);
  assign n2715 = n1880 | n1881;
  assign n2716 = (n2300 & n2714) | (n2300 & n2715) | (n2714 & n2715);
  assign n2717 = (n1880 & n1881) | (n1880 & n2306) | (n1881 & n2306);
  assign n2718 = (n1880 & n1881) | (n1880 & n2705) | (n1881 & n2705);
  assign n2719 = (n2290 & n2717) | (n2290 & n2718) | (n2717 & n2718);
  assign n2316 = (n2281 & n2716) | (n2281 & n2719) | (n2716 & n2719);
  assign n1883 = n1422 | n1878;
  assign n1884 = n1413 | n1422;
  assign n2720 = (n1406 & n1883) | (n1406 & n1884) | (n1883 & n1884);
  assign n2721 = n1883 | n1884;
  assign n2722 = (n2300 & n2720) | (n2300 & n2721) | (n2720 & n2721);
  assign n2723 = (n1883 & n1884) | (n1883 & n2306) | (n1884 & n2306);
  assign n2724 = (n1883 & n1884) | (n1883 & n2705) | (n1884 & n2705);
  assign n2725 = (n2290 & n2723) | (n2290 & n2724) | (n2723 & n2724);
  assign n2319 = (n2281 & n2722) | (n2281 & n2725) | (n2722 & n2725);
  assign n1425 = ~n2316 & n2319;
  assign n1876 = n1406 | n2300;
  assign n1427 = x143 & x207;
  assign n1428 = x143 | x207;
  assign n1429 = ~n1427 & n1428;
  assign n2320 = n1420 | n1422;
  assign n2321 = (n1420 & n1878) | (n1420 & n2320) | (n1878 & n2320);
  assign n1889 = n1429 & n2321;
  assign n2322 = n1413 | n1420;
  assign n2323 = (n1420 & n1422) | (n1420 & n2322) | (n1422 & n2322);
  assign n1890 = n1429 & n2323;
  assign n2324 = (n1876 & n1889) | (n1876 & n1890) | (n1889 & n1890);
  assign n2307 = (n2290 & n2705) | (n2290 & n2306) | (n2705 & n2306);
  assign n2325 = (n1889 & n1890) | (n1889 & n2307) | (n1890 & n2307);
  assign n2326 = (n2281 & n2324) | (n2281 & n2325) | (n2324 & n2325);
  assign n1892 = n1429 | n2321;
  assign n1893 = n1429 | n2323;
  assign n2327 = (n1876 & n1892) | (n1876 & n1893) | (n1892 & n1893);
  assign n2328 = (n1892 & n1893) | (n1892 & n2307) | (n1893 & n2307);
  assign n2329 = (n2281 & n2327) | (n2281 & n2328) | (n2327 & n2328);
  assign n1432 = ~n2326 & n2329;
  assign n1434 = x144 & x208;
  assign n1435 = x144 | x208;
  assign n1436 = ~n1434 & n1435;
  assign n2330 = n1427 | n1429;
  assign n2335 = (n1427 & n2323) | (n1427 & n2330) | (n2323 & n2330);
  assign n1899 = n1436 & n2335;
  assign n2332 = n1436 & n2330;
  assign n2333 = n1427 & n1436;
  assign n2334 = (n2321 & n2332) | (n2321 & n2333) | (n2332 & n2333);
  assign n2336 = (n1876 & n1899) | (n1876 & n2334) | (n1899 & n2334);
  assign n2337 = (n1899 & n2307) | (n1899 & n2334) | (n2307 & n2334);
  assign n2338 = (n2281 & n2336) | (n2281 & n2337) | (n2336 & n2337);
  assign n1902 = n1436 | n2335;
  assign n2339 = n1436 | n2330;
  assign n2340 = n1427 | n1436;
  assign n2341 = (n2321 & n2339) | (n2321 & n2340) | (n2339 & n2340);
  assign n2342 = (n1876 & n1902) | (n1876 & n2341) | (n1902 & n2341);
  assign n2343 = (n1902 & n2307) | (n1902 & n2341) | (n2307 & n2341);
  assign n2344 = (n2281 & n2342) | (n2281 & n2343) | (n2342 & n2343);
  assign n1439 = ~n2338 & n2344;
  assign n1441 = x145 & x209;
  assign n1442 = x145 | x209;
  assign n1443 = ~n1441 & n1442;
  assign n2345 = n1434 & n1443;
  assign n2346 = (n1443 & n2334) | (n1443 & n2345) | (n2334 & n2345);
  assign n2347 = n1434 | n1436;
  assign n2349 = n1443 & n2347;
  assign n2350 = (n2335 & n2345) | (n2335 & n2349) | (n2345 & n2349);
  assign n2351 = (n1876 & n2346) | (n1876 & n2350) | (n2346 & n2350);
  assign n2352 = (n2307 & n2346) | (n2307 & n2350) | (n2346 & n2350);
  assign n2353 = (n2281 & n2351) | (n2281 & n2352) | (n2351 & n2352);
  assign n2354 = n1434 | n1443;
  assign n2355 = n2334 | n2354;
  assign n2356 = n1443 | n2347;
  assign n2357 = (n2335 & n2354) | (n2335 & n2356) | (n2354 & n2356);
  assign n2358 = (n1876 & n2355) | (n1876 & n2357) | (n2355 & n2357);
  assign n2359 = (n2307 & n2355) | (n2307 & n2357) | (n2355 & n2357);
  assign n2360 = (n2281 & n2358) | (n2281 & n2359) | (n2358 & n2359);
  assign n1446 = ~n2353 & n2360;
  assign n1448 = x146 & x210;
  assign n1449 = x146 | x210;
  assign n1450 = ~n1448 & n1449;
  assign n2726 = n1434 | n1441;
  assign n2727 = (n1441 & n1443) | (n1441 & n2726) | (n1443 & n2726);
  assign n2364 = n1450 & n2727;
  assign n2362 = n1441 | n1443;
  assign n2365 = n1450 & n2362;
  assign n2366 = (n2334 & n2364) | (n2334 & n2365) | (n2364 & n2365);
  assign n2367 = n1441 & n1450;
  assign n2368 = (n1450 & n2350) | (n1450 & n2367) | (n2350 & n2367);
  assign n2369 = (n1876 & n2366) | (n1876 & n2368) | (n2366 & n2368);
  assign n2370 = (n2307 & n2366) | (n2307 & n2368) | (n2366 & n2368);
  assign n2371 = (n2281 & n2369) | (n2281 & n2370) | (n2369 & n2370);
  assign n2372 = n1450 | n2727;
  assign n2373 = n1450 | n2362;
  assign n2374 = (n2334 & n2372) | (n2334 & n2373) | (n2372 & n2373);
  assign n2375 = n1441 | n1450;
  assign n2376 = n2350 | n2375;
  assign n2377 = (n1876 & n2374) | (n1876 & n2376) | (n2374 & n2376);
  assign n2378 = (n2307 & n2374) | (n2307 & n2376) | (n2374 & n2376);
  assign n2379 = (n2281 & n2377) | (n2281 & n2378) | (n2377 & n2378);
  assign n1453 = ~n2371 & n2379;
  assign n1455 = x147 & x211;
  assign n1456 = x147 | x211;
  assign n1457 = ~n1455 & n1456;
  assign n1922 = n1448 & n1457;
  assign n2380 = (n1457 & n1922) | (n1457 & n2370) | (n1922 & n2370);
  assign n2381 = (n1457 & n1922) | (n1457 & n2369) | (n1922 & n2369);
  assign n2382 = (n2281 & n2380) | (n2281 & n2381) | (n2380 & n2381);
  assign n1924 = n1448 | n1457;
  assign n2383 = n1924 | n2370;
  assign n2384 = n1924 | n2369;
  assign n2385 = (n2281 & n2383) | (n2281 & n2384) | (n2383 & n2384);
  assign n1460 = ~n2382 & n2385;
  assign n1462 = x148 & x212;
  assign n1463 = x148 | x212;
  assign n1464 = ~n1462 & n1463;
  assign n2386 = n1448 | n1455;
  assign n2387 = (n1455 & n1457) | (n1455 & n2386) | (n1457 & n2386);
  assign n1929 = n1464 & n2387;
  assign n1927 = n1455 | n1457;
  assign n1930 = n1464 & n1927;
  assign n2388 = (n1929 & n1930) | (n1929 & n2370) | (n1930 & n2370);
  assign n2389 = (n1929 & n1930) | (n1929 & n2369) | (n1930 & n2369);
  assign n2390 = (n2281 & n2388) | (n2281 & n2389) | (n2388 & n2389);
  assign n1932 = n1464 | n2387;
  assign n1933 = n1464 | n1927;
  assign n2391 = (n1932 & n1933) | (n1932 & n2370) | (n1933 & n2370);
  assign n2392 = (n1932 & n1933) | (n1932 & n2369) | (n1933 & n2369);
  assign n2393 = (n2281 & n2391) | (n2281 & n2392) | (n2391 & n2392);
  assign n1467 = ~n2390 & n2393;
  assign n1469 = x149 & x213;
  assign n1470 = x149 | x213;
  assign n1471 = ~n1469 & n1470;
  assign n2394 = n1462 | n1464;
  assign n2395 = (n1462 & n2387) | (n1462 & n2394) | (n2387 & n2394);
  assign n1938 = n1471 & n2395;
  assign n2396 = (n1462 & n1927) | (n1462 & n2394) | (n1927 & n2394);
  assign n1939 = n1471 & n2396;
  assign n2397 = (n1938 & n1939) | (n1938 & n2370) | (n1939 & n2370);
  assign n2398 = (n1938 & n1939) | (n1938 & n2369) | (n1939 & n2369);
  assign n2399 = (n2281 & n2397) | (n2281 & n2398) | (n2397 & n2398);
  assign n1941 = n1471 | n2395;
  assign n1942 = n1471 | n2396;
  assign n2400 = (n1941 & n1942) | (n1941 & n2370) | (n1942 & n2370);
  assign n2401 = (n1941 & n1942) | (n1941 & n2369) | (n1942 & n2369);
  assign n2402 = (n2281 & n2400) | (n2281 & n2401) | (n2400 & n2401);
  assign n1474 = ~n2399 & n2402;
  assign n1476 = x150 & x214;
  assign n1477 = x150 | x214;
  assign n1478 = ~n1476 & n1477;
  assign n2403 = n1469 | n1471;
  assign n2405 = n1478 & n2403;
  assign n2406 = n1469 & n1478;
  assign n2407 = (n2395 & n2405) | (n2395 & n2406) | (n2405 & n2406);
  assign n2409 = (n2396 & n2405) | (n2396 & n2406) | (n2405 & n2406);
  assign n2410 = (n2370 & n2407) | (n2370 & n2409) | (n2407 & n2409);
  assign n2411 = (n2369 & n2407) | (n2369 & n2409) | (n2407 & n2409);
  assign n2412 = (n2281 & n2410) | (n2281 & n2411) | (n2410 & n2411);
  assign n2413 = n1478 | n2403;
  assign n2414 = n1469 | n1478;
  assign n2415 = (n2395 & n2413) | (n2395 & n2414) | (n2413 & n2414);
  assign n2416 = (n2396 & n2413) | (n2396 & n2414) | (n2413 & n2414);
  assign n2417 = (n2370 & n2415) | (n2370 & n2416) | (n2415 & n2416);
  assign n2418 = (n2369 & n2415) | (n2369 & n2416) | (n2415 & n2416);
  assign n2419 = (n2281 & n2417) | (n2281 & n2418) | (n2417 & n2418);
  assign n1481 = ~n2412 & n2419;
  assign n1483 = x151 & x215;
  assign n1484 = x151 | x215;
  assign n1485 = ~n1483 & n1484;
  assign n2420 = n1476 & n1485;
  assign n2421 = (n1485 & n2407) | (n1485 & n2420) | (n2407 & n2420);
  assign n2422 = (n1485 & n2409) | (n1485 & n2420) | (n2409 & n2420);
  assign n2423 = (n2370 & n2421) | (n2370 & n2422) | (n2421 & n2422);
  assign n2424 = (n2369 & n2421) | (n2369 & n2422) | (n2421 & n2422);
  assign n2425 = (n2281 & n2423) | (n2281 & n2424) | (n2423 & n2424);
  assign n2426 = n1476 | n1485;
  assign n2427 = n2407 | n2426;
  assign n2428 = n2409 | n2426;
  assign n2429 = (n2370 & n2427) | (n2370 & n2428) | (n2427 & n2428);
  assign n2430 = (n2369 & n2427) | (n2369 & n2428) | (n2427 & n2428);
  assign n2431 = (n2281 & n2429) | (n2281 & n2430) | (n2429 & n2430);
  assign n1488 = ~n2425 & n2431;
  assign n1490 = x152 & x216;
  assign n1491 = x152 | x216;
  assign n1492 = ~n1490 & n1491;
  assign n2728 = n1476 | n1483;
  assign n2729 = (n1483 & n1485) | (n1483 & n2728) | (n1485 & n2728);
  assign n2435 = n1492 & n2729;
  assign n2433 = n1483 | n1485;
  assign n2436 = n1492 & n2433;
  assign n2437 = (n2407 & n2435) | (n2407 & n2436) | (n2435 & n2436);
  assign n2439 = (n2409 & n2435) | (n2409 & n2436) | (n2435 & n2436);
  assign n2440 = (n2370 & n2437) | (n2370 & n2439) | (n2437 & n2439);
  assign n2441 = (n2369 & n2437) | (n2369 & n2439) | (n2437 & n2439);
  assign n2442 = (n2281 & n2440) | (n2281 & n2441) | (n2440 & n2441);
  assign n2443 = n1492 | n2729;
  assign n2444 = n1492 | n2433;
  assign n2445 = (n2407 & n2443) | (n2407 & n2444) | (n2443 & n2444);
  assign n2446 = (n2409 & n2443) | (n2409 & n2444) | (n2443 & n2444);
  assign n2447 = (n2370 & n2445) | (n2370 & n2446) | (n2445 & n2446);
  assign n2448 = (n2369 & n2445) | (n2369 & n2446) | (n2445 & n2446);
  assign n2449 = (n2281 & n2447) | (n2281 & n2448) | (n2447 & n2448);
  assign n1495 = ~n2442 & n2449;
  assign n1497 = x153 & x217;
  assign n1498 = x153 | x217;
  assign n1499 = ~n1497 & n1498;
  assign n1971 = n1490 & n1499;
  assign n1972 = (n1499 & n2442) | (n1499 & n1971) | (n2442 & n1971);
  assign n1973 = n1490 | n1499;
  assign n1974 = n2442 | n1973;
  assign n1502 = ~n1972 & n1974;
  assign n1504 = x154 & x218;
  assign n1505 = x154 | x218;
  assign n1506 = ~n1504 & n1505;
  assign n2450 = n1490 | n1497;
  assign n2451 = (n1497 & n1499) | (n1497 & n2450) | (n1499 & n2450);
  assign n1978 = n1506 & n2451;
  assign n1976 = n1497 | n1499;
  assign n1979 = n1506 & n1976;
  assign n1980 = (n2442 & n1978) | (n2442 & n1979) | (n1978 & n1979);
  assign n1981 = n1506 | n2451;
  assign n1982 = n1506 | n1976;
  assign n1983 = (n2442 & n1981) | (n2442 & n1982) | (n1981 & n1982);
  assign n1509 = ~n1980 & n1983;
  assign n1511 = x155 & x219;
  assign n1512 = x155 | x219;
  assign n1513 = ~n1511 & n1512;
  assign n2452 = n1504 | n1506;
  assign n2453 = (n1504 & n2451) | (n1504 & n2452) | (n2451 & n2452);
  assign n1987 = n1513 & n2453;
  assign n2454 = (n1504 & n1976) | (n1504 & n2452) | (n1976 & n2452);
  assign n1988 = n1513 & n2454;
  assign n1989 = (n2442 & n1987) | (n2442 & n1988) | (n1987 & n1988);
  assign n1990 = n1513 | n2453;
  assign n1991 = n1513 | n2454;
  assign n1992 = (n2442 & n1990) | (n2442 & n1991) | (n1990 & n1991);
  assign n1516 = ~n1989 & n1992;
  assign n1518 = x156 & x220;
  assign n1519 = x156 | x220;
  assign n1520 = ~n1518 & n1519;
  assign n2455 = n1511 | n1513;
  assign n2457 = n1520 & n2455;
  assign n2458 = n1511 & n1520;
  assign n2459 = (n2453 & n2457) | (n2453 & n2458) | (n2457 & n2458);
  assign n2461 = (n2454 & n2457) | (n2454 & n2458) | (n2457 & n2458);
  assign n1998 = (n2442 & n2459) | (n2442 & n2461) | (n2459 & n2461);
  assign n2462 = n1520 | n2455;
  assign n2463 = n1511 | n1520;
  assign n2464 = (n2453 & n2462) | (n2453 & n2463) | (n2462 & n2463);
  assign n2465 = (n2454 & n2462) | (n2454 & n2463) | (n2462 & n2463);
  assign n2001 = (n2442 & n2464) | (n2442 & n2465) | (n2464 & n2465);
  assign n1523 = ~n1998 & n2001;
  assign n1525 = x157 & x221;
  assign n1526 = x157 | x221;
  assign n1527 = ~n1525 & n1526;
  assign n2466 = n1518 & n1527;
  assign n2467 = (n1527 & n2459) | (n1527 & n2466) | (n2459 & n2466);
  assign n2468 = (n1527 & n2461) | (n1527 & n2466) | (n2461 & n2466);
  assign n2007 = (n2442 & n2467) | (n2442 & n2468) | (n2467 & n2468);
  assign n2469 = n1518 | n1527;
  assign n2470 = n2459 | n2469;
  assign n2471 = n2461 | n2469;
  assign n2010 = (n2442 & n2470) | (n2442 & n2471) | (n2470 & n2471);
  assign n1530 = ~n2007 & n2010;
  assign n1532 = x158 & x222;
  assign n1533 = x158 | x222;
  assign n1534 = ~n1532 & n1533;
  assign n2730 = n1518 | n1525;
  assign n2731 = (n1525 & n1527) | (n1525 & n2730) | (n1527 & n2730);
  assign n2475 = n1534 & n2731;
  assign n2473 = n1525 | n1527;
  assign n2476 = n1534 & n2473;
  assign n2477 = (n2459 & n2475) | (n2459 & n2476) | (n2475 & n2476);
  assign n2479 = (n2461 & n2475) | (n2461 & n2476) | (n2475 & n2476);
  assign n2016 = (n2442 & n2477) | (n2442 & n2479) | (n2477 & n2479);
  assign n2480 = n1534 | n2731;
  assign n2481 = n1534 | n2473;
  assign n2482 = (n2459 & n2480) | (n2459 & n2481) | (n2480 & n2481);
  assign n2483 = (n2461 & n2480) | (n2461 & n2481) | (n2480 & n2481);
  assign n2019 = (n2442 & n2482) | (n2442 & n2483) | (n2482 & n2483);
  assign n1537 = ~n2016 & n2019;
  assign n1539 = x159 & x223;
  assign n1540 = x159 | x223;
  assign n1541 = ~n1539 & n1540;
  assign n2732 = n1532 | n2476;
  assign n2733 = n1532 | n2475;
  assign n2734 = (n2461 & n2732) | (n2461 & n2733) | (n2732 & n2733);
  assign n2484 = n1541 & n2734;
  assign n2735 = (n2459 & n2732) | (n2459 & n2733) | (n2732 & n2733);
  assign n2485 = n1541 & n2735;
  assign n2486 = (n2442 & n2484) | (n2442 & n2485) | (n2484 & n2485);
  assign n2487 = n1541 | n2734;
  assign n2488 = n1541 | n2735;
  assign n2489 = (n2442 & n2487) | (n2442 & n2488) | (n2487 & n2488);
  assign n1544 = ~n2486 & n2489;
  assign n1546 = x160 & x224;
  assign n1547 = x160 | x224;
  assign n1548 = ~n1546 & n1547;
  assign n2023 = n1539 | n1541;
  assign n2025 = n1548 & n2023;
  assign n2026 = n1539 & n1548;
  assign n2490 = (n2734 & n2025) | (n2734 & n2026) | (n2025 & n2026);
  assign n2491 = (n2735 & n2025) | (n2735 & n2026) | (n2025 & n2026);
  assign n2492 = (n2442 & n2490) | (n2442 & n2491) | (n2490 & n2491);
  assign n2028 = n1548 | n2023;
  assign n2029 = n1539 | n1548;
  assign n2493 = (n2734 & n2028) | (n2734 & n2029) | (n2028 & n2029);
  assign n2494 = (n2735 & n2028) | (n2735 & n2029) | (n2028 & n2029);
  assign n2495 = (n2442 & n2493) | (n2442 & n2494) | (n2493 & n2494);
  assign n1551 = ~n2492 & n2495;
  assign n1553 = x161 & x225;
  assign n1554 = x161 | x225;
  assign n1555 = ~n1553 & n1554;
  assign n2496 = n1546 | n1548;
  assign n2497 = (n1546 & n2023) | (n1546 & n2496) | (n2023 & n2496);
  assign n2034 = n1555 & n2497;
  assign n2498 = n1539 | n1546;
  assign n2499 = (n1546 & n1548) | (n1546 & n2498) | (n1548 & n2498);
  assign n2035 = n1555 & n2499;
  assign n2500 = (n2734 & n2034) | (n2734 & n2035) | (n2034 & n2035);
  assign n2501 = (n2735 & n2034) | (n2735 & n2035) | (n2034 & n2035);
  assign n2502 = (n2442 & n2500) | (n2442 & n2501) | (n2500 & n2501);
  assign n2037 = n1555 | n2497;
  assign n2038 = n1555 | n2499;
  assign n2503 = (n2734 & n2037) | (n2734 & n2038) | (n2037 & n2038);
  assign n2504 = (n2735 & n2037) | (n2735 & n2038) | (n2037 & n2038);
  assign n2505 = (n2442 & n2503) | (n2442 & n2504) | (n2503 & n2504);
  assign n1558 = ~n2502 & n2505;
  assign n1560 = x162 & x226;
  assign n1561 = x162 | x226;
  assign n1562 = ~n1560 & n1561;
  assign n2506 = n1553 | n1555;
  assign n2511 = (n1553 & n2499) | (n1553 & n2506) | (n2499 & n2506);
  assign n2044 = n1562 & n2511;
  assign n2508 = n1562 & n2506;
  assign n2509 = n1553 & n1562;
  assign n2510 = (n2497 & n2508) | (n2497 & n2509) | (n2508 & n2509);
  assign n2512 = (n2734 & n2044) | (n2734 & n2510) | (n2044 & n2510);
  assign n2513 = (n2735 & n2044) | (n2735 & n2510) | (n2044 & n2510);
  assign n2514 = (n2442 & n2512) | (n2442 & n2513) | (n2512 & n2513);
  assign n2047 = n1562 | n2511;
  assign n2515 = n1562 | n2506;
  assign n2516 = n1553 | n1562;
  assign n2517 = (n2497 & n2515) | (n2497 & n2516) | (n2515 & n2516);
  assign n2518 = (n2734 & n2047) | (n2734 & n2517) | (n2047 & n2517);
  assign n2519 = (n2735 & n2047) | (n2735 & n2517) | (n2047 & n2517);
  assign n2520 = (n2442 & n2518) | (n2442 & n2519) | (n2518 & n2519);
  assign n1565 = ~n2514 & n2520;
  assign n1567 = x163 & x227;
  assign n1568 = x163 | x227;
  assign n1569 = ~n1567 & n1568;
  assign n2521 = n1560 & n1569;
  assign n2522 = (n1569 & n2510) | (n1569 & n2521) | (n2510 & n2521);
  assign n2523 = n1560 | n1562;
  assign n2525 = n1569 & n2523;
  assign n2526 = (n2511 & n2521) | (n2511 & n2525) | (n2521 & n2525);
  assign n2527 = (n2734 & n2522) | (n2734 & n2526) | (n2522 & n2526);
  assign n2528 = (n2735 & n2522) | (n2735 & n2526) | (n2522 & n2526);
  assign n2529 = (n2442 & n2527) | (n2442 & n2528) | (n2527 & n2528);
  assign n2530 = n1560 | n1569;
  assign n2531 = n2510 | n2530;
  assign n2532 = n1569 | n2523;
  assign n2533 = (n2511 & n2530) | (n2511 & n2532) | (n2530 & n2532);
  assign n2534 = (n2734 & n2531) | (n2734 & n2533) | (n2531 & n2533);
  assign n2535 = (n2735 & n2531) | (n2735 & n2533) | (n2531 & n2533);
  assign n2536 = (n2442 & n2534) | (n2442 & n2535) | (n2534 & n2535);
  assign n1572 = ~n2529 & n2536;
  assign n1574 = x164 & x228;
  assign n1575 = x164 | x228;
  assign n1576 = ~n1574 & n1575;
  assign n2736 = n1560 | n1567;
  assign n2737 = (n1567 & n1569) | (n1567 & n2736) | (n1569 & n2736);
  assign n2540 = n1576 & n2737;
  assign n2538 = n1567 | n1569;
  assign n2541 = n1576 & n2538;
  assign n2542 = (n2510 & n2540) | (n2510 & n2541) | (n2540 & n2541);
  assign n2543 = n1567 & n1576;
  assign n2544 = (n1576 & n2526) | (n1576 & n2543) | (n2526 & n2543);
  assign n2545 = (n2734 & n2542) | (n2734 & n2544) | (n2542 & n2544);
  assign n2546 = (n2735 & n2542) | (n2735 & n2544) | (n2542 & n2544);
  assign n2547 = (n2442 & n2545) | (n2442 & n2546) | (n2545 & n2546);
  assign n2548 = n1576 | n2737;
  assign n2549 = n1576 | n2538;
  assign n2550 = (n2510 & n2548) | (n2510 & n2549) | (n2548 & n2549);
  assign n2551 = n1567 | n1576;
  assign n2552 = n2526 | n2551;
  assign n2553 = (n2734 & n2550) | (n2734 & n2552) | (n2550 & n2552);
  assign n2554 = (n2735 & n2550) | (n2735 & n2552) | (n2550 & n2552);
  assign n2555 = (n2442 & n2553) | (n2442 & n2554) | (n2553 & n2554);
  assign n1579 = ~n2547 & n2555;
  assign n1581 = x165 & x229;
  assign n1582 = x165 | x229;
  assign n1583 = ~n1581 & n1582;
  assign n2556 = n1574 & n1583;
  assign n2738 = (n1583 & n2541) | (n1583 & n2556) | (n2541 & n2556);
  assign n2739 = (n1583 & n2540) | (n1583 & n2556) | (n2540 & n2556);
  assign n2740 = (n2510 & n2738) | (n2510 & n2739) | (n2738 & n2739);
  assign n2741 = n1567 | n1574;
  assign n2742 = (n1574 & n1576) | (n1574 & n2741) | (n1576 & n2741);
  assign n2561 = n1583 & n2742;
  assign n2559 = n1574 | n1576;
  assign n2562 = n1583 & n2559;
  assign n2563 = (n2526 & n2561) | (n2526 & n2562) | (n2561 & n2562);
  assign n2564 = (n2734 & n2740) | (n2734 & n2563) | (n2740 & n2563);
  assign n2565 = (n2735 & n2740) | (n2735 & n2563) | (n2740 & n2563);
  assign n2566 = (n2442 & n2564) | (n2442 & n2565) | (n2564 & n2565);
  assign n2567 = n1574 | n1583;
  assign n2743 = n2541 | n2567;
  assign n2744 = n2540 | n2567;
  assign n2745 = (n2510 & n2743) | (n2510 & n2744) | (n2743 & n2744);
  assign n2569 = n1583 | n2742;
  assign n2570 = n1583 | n2559;
  assign n2571 = (n2526 & n2569) | (n2526 & n2570) | (n2569 & n2570);
  assign n2572 = (n2734 & n2745) | (n2734 & n2571) | (n2745 & n2571);
  assign n2573 = (n2735 & n2745) | (n2735 & n2571) | (n2745 & n2571);
  assign n2574 = (n2442 & n2572) | (n2442 & n2573) | (n2572 & n2573);
  assign n1586 = ~n2566 & n2574;
  assign n1588 = x166 & x230;
  assign n1589 = x166 | x230;
  assign n1590 = ~n1588 & n1589;
  assign n2746 = n1581 | n2562;
  assign n2747 = n1581 | n2561;
  assign n2748 = (n2526 & n2746) | (n2526 & n2747) | (n2746 & n2747);
  assign n2576 = n1581 | n1583;
  assign n2749 = n1574 | n1581;
  assign n2750 = (n1581 & n1583) | (n1581 & n2749) | (n1583 & n2749);
  assign n2751 = (n2541 & n2576) | (n2541 & n2750) | (n2576 & n2750);
  assign n2752 = (n2540 & n2576) | (n2540 & n2750) | (n2576 & n2750);
  assign n2753 = (n2510 & n2751) | (n2510 & n2752) | (n2751 & n2752);
  assign n2579 = (n2735 & n2748) | (n2735 & n2753) | (n2748 & n2753);
  assign n2581 = n1590 & n2579;
  assign n2578 = (n2734 & n2748) | (n2734 & n2753) | (n2748 & n2753);
  assign n2582 = n1590 & n2578;
  assign n2583 = (n2442 & n2581) | (n2442 & n2582) | (n2581 & n2582);
  assign n2584 = n1590 | n2579;
  assign n2585 = n1590 | n2578;
  assign n2586 = (n2442 & n2584) | (n2442 & n2585) | (n2584 & n2585);
  assign n1593 = ~n2583 & n2586;
  assign n1595 = x167 & x231;
  assign n1596 = x167 | x231;
  assign n1597 = ~n1595 & n1596;
  assign n2079 = n1588 | n1590;
  assign n2081 = n1597 & n2079;
  assign n2082 = n1588 & n1597;
  assign n2587 = (n2081 & n2082) | (n2081 & n2579) | (n2082 & n2579);
  assign n2588 = (n2081 & n2082) | (n2081 & n2578) | (n2082 & n2578);
  assign n2589 = (n2442 & n2587) | (n2442 & n2588) | (n2587 & n2588);
  assign n2084 = n1597 | n2079;
  assign n2085 = n1588 | n1597;
  assign n2590 = (n2084 & n2085) | (n2084 & n2579) | (n2085 & n2579);
  assign n2591 = (n2084 & n2085) | (n2084 & n2578) | (n2085 & n2578);
  assign n2592 = (n2442 & n2590) | (n2442 & n2591) | (n2590 & n2591);
  assign n1600 = ~n2589 & n2592;
  assign n1602 = x168 & x232;
  assign n1603 = x168 | x232;
  assign n1604 = ~n1602 & n1603;
  assign n2593 = n1595 | n1597;
  assign n2594 = (n1595 & n2079) | (n1595 & n2593) | (n2079 & n2593);
  assign n2090 = n1604 & n2594;
  assign n2595 = n1588 | n1595;
  assign n2596 = (n1595 & n1597) | (n1595 & n2595) | (n1597 & n2595);
  assign n2091 = n1604 & n2596;
  assign n2597 = (n2090 & n2091) | (n2090 & n2579) | (n2091 & n2579);
  assign n2598 = (n2090 & n2091) | (n2090 & n2578) | (n2091 & n2578);
  assign n2599 = (n2442 & n2597) | (n2442 & n2598) | (n2597 & n2598);
  assign n2093 = n1604 | n2594;
  assign n2094 = n1604 | n2596;
  assign n2600 = (n2093 & n2094) | (n2093 & n2579) | (n2094 & n2579);
  assign n2601 = (n2093 & n2094) | (n2093 & n2578) | (n2094 & n2578);
  assign n2602 = (n2442 & n2600) | (n2442 & n2601) | (n2600 & n2601);
  assign n1607 = ~n2599 & n2602;
  assign n1609 = x169 & x233;
  assign n1610 = x169 | x233;
  assign n1611 = ~n1609 & n1610;
  assign n2603 = n1602 | n1604;
  assign n2608 = (n1602 & n2596) | (n1602 & n2603) | (n2596 & n2603);
  assign n2100 = n1611 & n2608;
  assign n2605 = n1611 & n2603;
  assign n2606 = n1602 & n1611;
  assign n2607 = (n2594 & n2605) | (n2594 & n2606) | (n2605 & n2606);
  assign n2609 = (n2100 & n2579) | (n2100 & n2607) | (n2579 & n2607);
  assign n2610 = (n2100 & n2578) | (n2100 & n2607) | (n2578 & n2607);
  assign n2611 = (n2442 & n2609) | (n2442 & n2610) | (n2609 & n2610);
  assign n2103 = n1611 | n2608;
  assign n2612 = n1611 | n2603;
  assign n2613 = n1602 | n1611;
  assign n2614 = (n2594 & n2612) | (n2594 & n2613) | (n2612 & n2613);
  assign n2615 = (n2103 & n2579) | (n2103 & n2614) | (n2579 & n2614);
  assign n2616 = (n2103 & n2578) | (n2103 & n2614) | (n2578 & n2614);
  assign n2617 = (n2442 & n2615) | (n2442 & n2616) | (n2615 & n2616);
  assign n1614 = ~n2611 & n2617;
  assign n1616 = x170 & x234;
  assign n1617 = x170 | x234;
  assign n1618 = ~n1616 & n1617;
  assign n2618 = n1609 & n1618;
  assign n2619 = (n1618 & n2607) | (n1618 & n2618) | (n2607 & n2618);
  assign n2620 = n1609 | n1611;
  assign n2622 = n1618 & n2620;
  assign n2623 = (n2608 & n2618) | (n2608 & n2622) | (n2618 & n2622);
  assign n2624 = (n2579 & n2619) | (n2579 & n2623) | (n2619 & n2623);
  assign n2625 = (n2578 & n2619) | (n2578 & n2623) | (n2619 & n2623);
  assign n2626 = (n2442 & n2624) | (n2442 & n2625) | (n2624 & n2625);
  assign n2627 = n1609 | n1618;
  assign n2628 = n2607 | n2627;
  assign n2629 = n1618 | n2620;
  assign n2630 = (n2608 & n2627) | (n2608 & n2629) | (n2627 & n2629);
  assign n2631 = (n2579 & n2628) | (n2579 & n2630) | (n2628 & n2630);
  assign n2632 = (n2578 & n2628) | (n2578 & n2630) | (n2628 & n2630);
  assign n2633 = (n2442 & n2631) | (n2442 & n2632) | (n2631 & n2632);
  assign n1621 = ~n2626 & n2633;
  assign n1623 = x171 & x235;
  assign n1624 = x171 | x235;
  assign n1625 = ~n1623 & n1624;
  assign n2754 = n1609 | n1616;
  assign n2755 = (n1616 & n1618) | (n1616 & n2754) | (n1618 & n2754);
  assign n2637 = n1625 & n2755;
  assign n2635 = n1616 | n1618;
  assign n2638 = n1625 & n2635;
  assign n2639 = (n2607 & n2637) | (n2607 & n2638) | (n2637 & n2638);
  assign n2640 = n1616 & n1625;
  assign n2641 = (n1625 & n2623) | (n1625 & n2640) | (n2623 & n2640);
  assign n2642 = (n2579 & n2639) | (n2579 & n2641) | (n2639 & n2641);
  assign n2643 = (n2578 & n2639) | (n2578 & n2641) | (n2639 & n2641);
  assign n2644 = (n2442 & n2642) | (n2442 & n2643) | (n2642 & n2643);
  assign n2645 = n1625 | n2755;
  assign n2646 = n1625 | n2635;
  assign n2647 = (n2607 & n2645) | (n2607 & n2646) | (n2645 & n2646);
  assign n2648 = n1616 | n1625;
  assign n2649 = n2623 | n2648;
  assign n2650 = (n2579 & n2647) | (n2579 & n2649) | (n2647 & n2649);
  assign n2651 = (n2578 & n2647) | (n2578 & n2649) | (n2647 & n2649);
  assign n2652 = (n2442 & n2650) | (n2442 & n2651) | (n2650 & n2651);
  assign n1628 = ~n2644 & n2652;
  assign n1630 = x172 & x236;
  assign n1631 = x172 | x236;
  assign n1632 = ~n1630 & n1631;
  assign n2653 = n1623 & n1632;
  assign n2756 = (n1632 & n2638) | (n1632 & n2653) | (n2638 & n2653);
  assign n2757 = (n1632 & n2637) | (n1632 & n2653) | (n2637 & n2653);
  assign n2758 = (n2607 & n2756) | (n2607 & n2757) | (n2756 & n2757);
  assign n2759 = n1616 | n1623;
  assign n2760 = (n1623 & n1625) | (n1623 & n2759) | (n1625 & n2759);
  assign n2658 = n1632 & n2760;
  assign n2656 = n1623 | n1625;
  assign n2659 = n1632 & n2656;
  assign n2660 = (n2623 & n2658) | (n2623 & n2659) | (n2658 & n2659);
  assign n2661 = (n2579 & n2758) | (n2579 & n2660) | (n2758 & n2660);
  assign n2662 = (n2578 & n2758) | (n2578 & n2660) | (n2758 & n2660);
  assign n2663 = (n2442 & n2661) | (n2442 & n2662) | (n2661 & n2662);
  assign n2664 = n1623 | n1632;
  assign n2761 = n2638 | n2664;
  assign n2762 = n2637 | n2664;
  assign n2763 = (n2607 & n2761) | (n2607 & n2762) | (n2761 & n2762);
  assign n2666 = n1632 | n2760;
  assign n2667 = n1632 | n2656;
  assign n2668 = (n2623 & n2666) | (n2623 & n2667) | (n2666 & n2667);
  assign n2669 = (n2579 & n2763) | (n2579 & n2668) | (n2763 & n2668);
  assign n2670 = (n2578 & n2763) | (n2578 & n2668) | (n2763 & n2668);
  assign n2671 = (n2442 & n2669) | (n2442 & n2670) | (n2669 & n2670);
  assign n1635 = ~n2663 & n2671;
  assign n1637 = x173 & x237;
  assign n1638 = x173 | x237;
  assign n1639 = ~n1637 & n1638;
  assign n2764 = n1623 | n1630;
  assign n2765 = (n1630 & n1632) | (n1630 & n2764) | (n1632 & n2764);
  assign n2675 = n1639 & n2765;
  assign n2673 = n1630 | n1632;
  assign n2676 = n1639 & n2673;
  assign n2766 = (n2638 & n2675) | (n2638 & n2676) | (n2675 & n2676);
  assign n2767 = (n2637 & n2675) | (n2637 & n2676) | (n2675 & n2676);
  assign n2768 = (n2607 & n2766) | (n2607 & n2767) | (n2766 & n2767);
  assign n2678 = n1630 & n1639;
  assign n2769 = (n1639 & n2659) | (n1639 & n2678) | (n2659 & n2678);
  assign n2770 = (n1639 & n2658) | (n1639 & n2678) | (n2658 & n2678);
  assign n2771 = (n2623 & n2769) | (n2623 & n2770) | (n2769 & n2770);
  assign n2680 = (n2579 & n2768) | (n2579 & n2771) | (n2768 & n2771);
  assign n2681 = (n2578 & n2768) | (n2578 & n2771) | (n2768 & n2771);
  assign n2682 = (n2442 & n2680) | (n2442 & n2681) | (n2680 & n2681);
  assign n2683 = n1639 | n2765;
  assign n2684 = n1639 | n2673;
  assign n2772 = (n2638 & n2683) | (n2638 & n2684) | (n2683 & n2684);
  assign n2773 = (n2637 & n2683) | (n2637 & n2684) | (n2683 & n2684);
  assign n2774 = (n2607 & n2772) | (n2607 & n2773) | (n2772 & n2773);
  assign n2686 = n1630 | n1639;
  assign n2775 = n2659 | n2686;
  assign n2776 = n2658 | n2686;
  assign n2777 = (n2623 & n2775) | (n2623 & n2776) | (n2775 & n2776);
  assign n2688 = (n2579 & n2774) | (n2579 & n2777) | (n2774 & n2777);
  assign n2689 = (n2578 & n2774) | (n2578 & n2777) | (n2774 & n2777);
  assign n2690 = (n2442 & n2688) | (n2442 & n2689) | (n2688 & n2689);
  assign n1642 = ~n2682 & n2690;
  assign n1644 = x174 & x238;
  assign n1645 = x174 | x238;
  assign n1646 = ~n1644 & n1645;
  assign n2141 = n1637 & n1646;
  assign n2778 = (n1646 & n2141) | (n1646 & n2681) | (n2141 & n2681);
  assign n2779 = (n1646 & n2141) | (n1646 & n2680) | (n2141 & n2680);
  assign n2780 = (n2442 & n2778) | (n2442 & n2779) | (n2778 & n2779);
  assign n2143 = n1637 | n1646;
  assign n2781 = n2143 | n2681;
  assign n2782 = n2143 | n2680;
  assign n2783 = (n2442 & n2781) | (n2442 & n2782) | (n2781 & n2782);
  assign n1649 = ~n2780 & n2783;
  assign n1651 = x175 & x239;
  assign n1652 = x175 | x239;
  assign n1653 = ~n1651 & n1652;
  assign n2691 = n1637 | n1644;
  assign n2692 = (n1644 & n1646) | (n1644 & n2691) | (n1646 & n2691);
  assign n2148 = n1653 & n2692;
  assign n2146 = n1644 | n1646;
  assign n2149 = n1653 & n2146;
  assign n2784 = (n2148 & n2149) | (n2148 & n2681) | (n2149 & n2681);
  assign n2785 = (n2148 & n2149) | (n2148 & n2680) | (n2149 & n2680);
  assign n2786 = (n2442 & n2784) | (n2442 & n2785) | (n2784 & n2785);
  assign n2151 = n1653 | n2692;
  assign n2152 = n1653 | n2146;
  assign n2787 = (n2151 & n2152) | (n2151 & n2681) | (n2152 & n2681);
  assign n2788 = (n2151 & n2152) | (n2151 & n2680) | (n2152 & n2680);
  assign n2789 = (n2442 & n2787) | (n2442 & n2788) | (n2787 & n2788);
  assign n1656 = ~n2786 & n2789;
  assign n2693 = n1651 | n1653;
  assign n2694 = (n1651 & n2692) | (n1651 & n2693) | (n2692 & n2693);
  assign n2695 = (n1651 & n2146) | (n1651 & n2693) | (n2146 & n2693);
  assign n2790 = (n2681 & n2694) | (n2681 & n2695) | (n2694 & n2695);
  assign n2791 = (n2680 & n2694) | (n2680 & n2695) | (n2694 & n2695);
  assign n2792 = (n2442 & n2790) | (n2442 & n2791) | (n2790 & n2791);
  assign y0 = n19;
  assign y1 = n25;
  assign y2 = n32;
  assign y3 = n39;
  assign y4 = n46;
  assign y5 = n53;
  assign y6 = n60;
  assign y7 = n67;
  assign y8 = n113;
  assign y9 = n148;
  assign y10 = n154;
  assign y11 = n161;
  assign y12 = n168;
  assign y13 = n175;
  assign y14 = n182;
  assign y15 = n189;
  assign y16 = n196;
  assign y17 = n203;
  assign y18 = n210;
  assign y19 = n217;
  assign y20 = n224;
  assign y21 = n231;
  assign y22 = n238;
  assign y23 = n245;
  assign y24 = n252;
  assign y25 = n253;
  assign y26 = n473;
  assign y27 = n479;
  assign y28 = n486;
  assign y29 = n493;
  assign y30 = n500;
  assign y31 = n507;
  assign y32 = n514;
  assign y33 = n521;
  assign y34 = n528;
  assign y35 = n535;
  assign y36 = n542;
  assign y37 = n549;
  assign y38 = n556;
  assign y39 = n563;
  assign y40 = n570;
  assign y41 = n577;
  assign y42 = n584;
  assign y43 = n591;
  assign y44 = n598;
  assign y45 = n605;
  assign y46 = n612;
  assign y47 = n619;
  assign y48 = n626;
  assign y49 = n633;
  assign y50 = n640;
  assign y51 = n647;
  assign y52 = n654;
  assign y53 = n661;
  assign y54 = n668;
  assign y55 = n675;
  assign y56 = n682;
  assign y57 = n689;
  assign y58 = n1085;
  assign y59 = n1216;
  assign y60 = n1222;
  assign y61 = n1229;
  assign y62 = n1236;
  assign y63 = n1243;
  assign y64 = n1250;
  assign y65 = n1257;
  assign y66 = n1264;
  assign y67 = n1271;
  assign y68 = n1278;
  assign y69 = n1285;
  assign y70 = n1292;
  assign y71 = n1299;
  assign y72 = n1306;
  assign y73 = n1313;
  assign y74 = n1320;
  assign y75 = n1327;
  assign y76 = n1334;
  assign y77 = n1341;
  assign y78 = n1348;
  assign y79 = n1355;
  assign y80 = n1362;
  assign y81 = n1369;
  assign y82 = n1376;
  assign y83 = n1383;
  assign y84 = n1390;
  assign y85 = n1397;
  assign y86 = n1404;
  assign y87 = n1411;
  assign y88 = n1418;
  assign y89 = n1425;
  assign y90 = n1432;
  assign y91 = n1439;
  assign y92 = n1446;
  assign y93 = n1453;
  assign y94 = n1460;
  assign y95 = n1467;
  assign y96 = n1474;
  assign y97 = n1481;
  assign y98 = n1488;
  assign y99 = n1495;
  assign y100 = n1502;
  assign y101 = n1509;
  assign y102 = n1516;
  assign y103 = n1523;
  assign y104 = n1530;
  assign y105 = n1537;
  assign y106 = n1544;
  assign y107 = n1551;
  assign y108 = n1558;
  assign y109 = n1565;
  assign y110 = n1572;
  assign y111 = n1579;
  assign y112 = n1586;
  assign y113 = n1593;
  assign y114 = n1600;
  assign y115 = n1607;
  assign y116 = n1614;
  assign y117 = n1621;
  assign y118 = n1628;
  assign y119 = n1635;
  assign y120 = n1642;
  assign y121 = n1649;
  assign y122 = n1656;
  assign y123 = n2792;
endmodule

