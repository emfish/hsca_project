module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930;
  assign n17 = x0 & x8;
  assign n18 = x1 & x8;
  assign n19 = x0 & x9;
  assign n20 = n18 & n19;
  assign n21 = n18 | n19;
  assign n22 = ~n20 & n21;
  assign n23 = x2 & x8;
  assign n24 = x1 & x9;
  assign n25 = n23 & n24;
  assign n26 = n23 | n24;
  assign n27 = ~n25 & n26;
  assign n28 = n20 & n27;
  assign n29 = n20 | n27;
  assign n30 = ~n28 & n29;
  assign n31 = x0 & x10;
  assign n32 = n30 & n31;
  assign n33 = n30 | n31;
  assign n34 = ~n32 & n33;
  assign n441 = n20 | n25;
  assign n442 = (n25 & n27) | (n25 & n441) | (n27 & n441);
  assign n36 = x3 & x8;
  assign n37 = x2 & x9;
  assign n38 = n36 & n37;
  assign n39 = n36 | n37;
  assign n40 = ~n38 & n39;
  assign n41 = n442 & n40;
  assign n42 = n442 | n40;
  assign n43 = ~n41 & n42;
  assign n44 = x1 & x10;
  assign n45 = n43 & n44;
  assign n46 = n43 | n44;
  assign n47 = ~n45 & n46;
  assign n48 = n32 & n47;
  assign n49 = n32 | n47;
  assign n50 = ~n48 & n49;
  assign n51 = x0 & x11;
  assign n52 = n50 & n51;
  assign n53 = n50 | n51;
  assign n54 = ~n52 & n53;
  assign n443 = n32 | n45;
  assign n444 = (n45 & n47) | (n45 & n443) | (n47 & n443);
  assign n445 = n38 | n40;
  assign n446 = (n38 & n442) | (n38 & n445) | (n442 & n445);
  assign n57 = x4 & x8;
  assign n58 = x3 & x9;
  assign n59 = n57 & n58;
  assign n60 = n57 | n58;
  assign n61 = ~n59 & n60;
  assign n62 = n446 & n61;
  assign n63 = n446 | n61;
  assign n64 = ~n62 & n63;
  assign n65 = x2 & x10;
  assign n66 = n64 & n65;
  assign n67 = n64 | n65;
  assign n68 = ~n66 & n67;
  assign n69 = n444 & n68;
  assign n70 = n444 | n68;
  assign n71 = ~n69 & n70;
  assign n72 = x1 & x11;
  assign n73 = n71 & n72;
  assign n74 = n71 | n72;
  assign n75 = ~n73 & n74;
  assign n76 = n52 & n75;
  assign n77 = n52 | n75;
  assign n78 = ~n76 & n77;
  assign n79 = x0 & x12;
  assign n80 = n78 & n79;
  assign n81 = n78 | n79;
  assign n82 = ~n80 & n81;
  assign n447 = n52 | n73;
  assign n448 = (n73 & n75) | (n73 & n447) | (n75 & n447);
  assign n86 = x5 & x8;
  assign n87 = x4 & x9;
  assign n88 = n86 & n87;
  assign n89 = n86 | n87;
  assign n90 = ~n88 & n89;
  assign n449 = n59 | n61;
  assign n451 = n90 & n449;
  assign n452 = n59 & n90;
  assign n453 = (n446 & n451) | (n446 & n452) | (n451 & n452);
  assign n454 = n90 | n449;
  assign n455 = n59 | n90;
  assign n456 = (n446 & n454) | (n446 & n455) | (n454 & n455);
  assign n93 = ~n453 & n456;
  assign n94 = x3 & x10;
  assign n95 = n93 & n94;
  assign n96 = n93 | n94;
  assign n97 = ~n95 & n96;
  assign n457 = n66 & n97;
  assign n458 = (n69 & n97) | (n69 & n457) | (n97 & n457);
  assign n459 = n66 | n97;
  assign n460 = n69 | n459;
  assign n100 = ~n458 & n460;
  assign n101 = x2 & x11;
  assign n102 = n100 & n101;
  assign n103 = n100 | n101;
  assign n104 = ~n102 & n103;
  assign n105 = n448 & n104;
  assign n106 = n448 | n104;
  assign n107 = ~n105 & n106;
  assign n108 = x1 & x12;
  assign n109 = n107 & n108;
  assign n110 = n107 | n108;
  assign n111 = ~n109 & n110;
  assign n112 = n80 & n111;
  assign n113 = n80 | n111;
  assign n114 = ~n112 & n113;
  assign n115 = x0 & x13;
  assign n116 = n114 & n115;
  assign n117 = n114 | n115;
  assign n118 = ~n116 & n117;
  assign n461 = n80 | n109;
  assign n462 = (n109 & n111) | (n109 & n461) | (n111 & n461);
  assign n120 = n102 | n105;
  assign n123 = x6 & x8;
  assign n124 = x5 & x9;
  assign n125 = n123 & n124;
  assign n126 = n123 | n124;
  assign n127 = ~n125 & n126;
  assign n463 = n88 & n127;
  assign n464 = (n127 & n453) | (n127 & n463) | (n453 & n463);
  assign n465 = n88 | n127;
  assign n466 = n453 | n465;
  assign n130 = ~n464 & n466;
  assign n131 = x4 & x10;
  assign n132 = n130 & n131;
  assign n133 = n130 | n131;
  assign n134 = ~n132 & n133;
  assign n467 = n95 & n134;
  assign n468 = (n134 & n458) | (n134 & n467) | (n458 & n467);
  assign n469 = n95 | n134;
  assign n470 = n458 | n469;
  assign n137 = ~n468 & n470;
  assign n138 = x3 & x11;
  assign n139 = n137 & n138;
  assign n140 = n137 | n138;
  assign n141 = ~n139 & n140;
  assign n142 = n120 & n141;
  assign n143 = n120 | n141;
  assign n144 = ~n142 & n143;
  assign n145 = x2 & x12;
  assign n146 = n144 & n145;
  assign n147 = n144 | n145;
  assign n148 = ~n146 & n147;
  assign n149 = n462 & n148;
  assign n150 = n462 | n148;
  assign n151 = ~n149 & n150;
  assign n152 = x1 & x13;
  assign n153 = n151 & n152;
  assign n154 = n151 | n152;
  assign n155 = ~n153 & n154;
  assign n156 = n116 & n155;
  assign n157 = n116 | n155;
  assign n158 = ~n156 & n157;
  assign n159 = x0 & x14;
  assign n160 = n158 & n159;
  assign n161 = n158 | n159;
  assign n162 = ~n160 & n161;
  assign n724 = n115 | n152;
  assign n725 = (n114 & n152) | (n114 & n724) | (n152 & n724);
  assign n598 = (n116 & n151) | (n116 & n725) | (n151 & n725);
  assign n472 = (n153 & n155) | (n153 & n598) | (n155 & n598);
  assign n473 = n146 | n462;
  assign n474 = (n146 & n148) | (n146 & n473) | (n148 & n473);
  assign n475 = n139 | n141;
  assign n476 = (n120 & n139) | (n120 & n475) | (n139 & n475);
  assign n168 = x7 & x8;
  assign n169 = x6 & x9;
  assign n170 = n168 & n169;
  assign n171 = n168 | n169;
  assign n172 = ~n170 & n171;
  assign n599 = n88 | n125;
  assign n600 = (n125 & n127) | (n125 & n599) | (n127 & n599);
  assign n480 = n172 & n600;
  assign n478 = n125 | n127;
  assign n481 = n172 & n478;
  assign n482 = (n453 & n480) | (n453 & n481) | (n480 & n481);
  assign n483 = n172 | n600;
  assign n484 = n172 | n478;
  assign n485 = (n453 & n483) | (n453 & n484) | (n483 & n484);
  assign n175 = ~n482 & n485;
  assign n176 = x5 & x10;
  assign n177 = n175 & n176;
  assign n178 = n175 | n176;
  assign n179 = ~n177 & n178;
  assign n486 = n132 & n179;
  assign n487 = (n179 & n468) | (n179 & n486) | (n468 & n486);
  assign n488 = n132 | n179;
  assign n489 = n468 | n488;
  assign n182 = ~n487 & n489;
  assign n183 = x4 & x11;
  assign n184 = n182 & n183;
  assign n185 = n182 | n183;
  assign n186 = ~n184 & n185;
  assign n187 = n476 & n186;
  assign n188 = n476 | n186;
  assign n189 = ~n187 & n188;
  assign n190 = x3 & x12;
  assign n191 = n189 & n190;
  assign n192 = n189 | n190;
  assign n193 = ~n191 & n192;
  assign n194 = n474 & n193;
  assign n195 = n474 | n193;
  assign n196 = ~n194 & n195;
  assign n197 = x2 & x13;
  assign n198 = n196 & n197;
  assign n199 = n196 | n197;
  assign n200 = ~n198 & n199;
  assign n201 = n472 & n200;
  assign n202 = n472 | n200;
  assign n203 = ~n201 & n202;
  assign n204 = x1 & x14;
  assign n205 = n203 & n204;
  assign n206 = n203 | n204;
  assign n207 = ~n205 & n206;
  assign n208 = n160 & n207;
  assign n209 = n160 | n207;
  assign n210 = ~n208 & n209;
  assign n211 = x0 & x15;
  assign n212 = n210 & n211;
  assign n213 = n210 | n211;
  assign n214 = ~n212 & n213;
  assign n490 = n160 | n205;
  assign n491 = (n205 & n207) | (n205 & n490) | (n207 & n490);
  assign n216 = n198 | n201;
  assign n217 = n191 | n194;
  assign n492 = n184 | n186;
  assign n493 = (n184 & n476) | (n184 & n492) | (n476 & n492);
  assign n221 = x7 & x9;
  assign n497 = n170 & n221;
  assign n726 = (n172 & n221) | (n172 & n497) | (n221 & n497);
  assign n728 = (n478 & n726) | (n478 & n497) | (n726 & n497);
  assign n729 = (n600 & n726) | (n600 & n497) | (n726 & n497);
  assign n605 = (n453 & n728) | (n453 & n729) | (n728 & n729);
  assign n499 = n170 | n221;
  assign n730 = n172 | n499;
  assign n731 = (n478 & n499) | (n478 & n730) | (n499 & n730);
  assign n732 = (n499 & n600) | (n499 & n730) | (n600 & n730);
  assign n608 = (n453 & n731) | (n453 & n732) | (n731 & n732);
  assign n224 = ~n605 & n608;
  assign n225 = x6 & x10;
  assign n226 = n224 & n225;
  assign n227 = n224 | n225;
  assign n228 = ~n226 & n227;
  assign n495 = n177 | n179;
  assign n609 = n228 & n495;
  assign n601 = n132 | n177;
  assign n602 = (n177 & n179) | (n177 & n601) | (n179 & n601);
  assign n610 = n228 & n602;
  assign n611 = (n468 & n609) | (n468 & n610) | (n609 & n610);
  assign n612 = n228 | n495;
  assign n613 = n228 | n602;
  assign n614 = (n468 & n612) | (n468 & n613) | (n612 & n613);
  assign n231 = ~n611 & n614;
  assign n232 = x5 & x11;
  assign n233 = n231 & n232;
  assign n234 = n231 | n232;
  assign n235 = ~n233 & n234;
  assign n236 = n493 & n235;
  assign n237 = n493 | n235;
  assign n238 = ~n236 & n237;
  assign n239 = x4 & x12;
  assign n240 = n238 & n239;
  assign n241 = n238 | n239;
  assign n242 = ~n240 & n241;
  assign n243 = n217 & n242;
  assign n244 = n217 | n242;
  assign n245 = ~n243 & n244;
  assign n246 = x3 & x13;
  assign n247 = n245 & n246;
  assign n248 = n245 | n246;
  assign n249 = ~n247 & n248;
  assign n250 = n216 & n249;
  assign n251 = n216 | n249;
  assign n252 = ~n250 & n251;
  assign n253 = x2 & x14;
  assign n254 = n252 & n253;
  assign n255 = n252 | n253;
  assign n256 = ~n254 & n255;
  assign n257 = n491 & n256;
  assign n258 = n491 | n256;
  assign n259 = ~n257 & n258;
  assign n260 = x1 & x15;
  assign n261 = n259 & n260;
  assign n262 = n259 | n260;
  assign n263 = ~n261 & n262;
  assign n264 = n212 & n263;
  assign n265 = n212 | n263;
  assign n266 = ~n264 & n265;
  assign n733 = n211 | n260;
  assign n734 = (n210 & n260) | (n210 & n733) | (n260 & n733);
  assign n616 = (n212 & n259) | (n212 & n734) | (n259 & n734);
  assign n502 = (n261 & n263) | (n261 & n616) | (n263 & n616);
  assign n503 = n254 | n491;
  assign n504 = (n254 & n256) | (n254 & n503) | (n256 & n503);
  assign n269 = n247 | n250;
  assign n505 = n240 | n242;
  assign n506 = (n217 & n240) | (n217 & n505) | (n240 & n505);
  assign n273 = x7 & x10;
  assign n512 = n221 & n273;
  assign n617 = n170 & n512;
  assign n735 = (n172 & n512) | (n172 & n617) | (n512 & n617);
  assign n736 = n512 & n617;
  assign n737 = (n478 & n735) | (n478 & n736) | (n735 & n736);
  assign n738 = (n600 & n735) | (n600 & n736) | (n735 & n736);
  assign n620 = (n453 & n737) | (n453 & n738) | (n737 & n738);
  assign n515 = n221 | n273;
  assign n621 = (n170 & n273) | (n170 & n515) | (n273 & n515);
  assign n739 = (n172 & n515) | (n172 & n621) | (n515 & n621);
  assign n740 = n515 & n621;
  assign n741 = (n478 & n739) | (n478 & n740) | (n739 & n740);
  assign n742 = (n600 & n739) | (n600 & n740) | (n739 & n740);
  assign n624 = (n453 & n741) | (n453 & n742) | (n741 & n742);
  assign n276 = ~n620 & n624;
  assign n518 = n226 & n276;
  assign n625 = (n228 & n276) | (n228 & n518) | (n276 & n518);
  assign n626 = (n495 & n518) | (n495 & n625) | (n518 & n625);
  assign n627 = (n518 & n602) | (n518 & n625) | (n602 & n625);
  assign n628 = (n468 & n626) | (n468 & n627) | (n626 & n627);
  assign n521 = n226 | n276;
  assign n629 = n228 | n521;
  assign n630 = (n495 & n521) | (n495 & n629) | (n521 & n629);
  assign n631 = (n521 & n602) | (n521 & n629) | (n602 & n629);
  assign n632 = (n468 & n630) | (n468 & n631) | (n630 & n631);
  assign n279 = ~n628 & n632;
  assign n280 = x6 & x11;
  assign n281 = n279 & n280;
  assign n282 = n279 | n280;
  assign n283 = ~n281 & n282;
  assign n507 = n233 | n235;
  assign n633 = n283 & n507;
  assign n634 = n233 & n283;
  assign n635 = (n493 & n633) | (n493 & n634) | (n633 & n634);
  assign n636 = n283 | n507;
  assign n637 = n233 | n283;
  assign n638 = (n493 & n636) | (n493 & n637) | (n636 & n637);
  assign n286 = ~n635 & n638;
  assign n287 = x5 & x12;
  assign n288 = n286 & n287;
  assign n289 = n286 | n287;
  assign n290 = ~n288 & n289;
  assign n291 = n506 & n290;
  assign n292 = n506 | n290;
  assign n293 = ~n291 & n292;
  assign n294 = x4 & x13;
  assign n295 = n293 & n294;
  assign n296 = n293 | n294;
  assign n297 = ~n295 & n296;
  assign n298 = n269 & n297;
  assign n299 = n269 | n297;
  assign n300 = ~n298 & n299;
  assign n301 = x3 & x14;
  assign n302 = n300 & n301;
  assign n303 = n300 | n301;
  assign n304 = ~n302 & n303;
  assign n305 = n504 & n304;
  assign n306 = n504 | n304;
  assign n307 = ~n305 & n306;
  assign n308 = x2 & x15;
  assign n309 = n307 & n308;
  assign n310 = n307 | n308;
  assign n311 = ~n309 & n310;
  assign n312 = n502 & n311;
  assign n313 = n502 | n311;
  assign n314 = ~n312 & n313;
  assign n523 = n309 | n502;
  assign n524 = (n309 & n311) | (n309 & n523) | (n311 & n523);
  assign n525 = n302 | n504;
  assign n526 = (n302 & n304) | (n302 & n525) | (n304 & n525);
  assign n527 = n295 | n297;
  assign n528 = (n269 & n295) | (n269 & n527) | (n295 & n527);
  assign n321 = x7 & x11;
  assign n743 = n321 & n738;
  assign n744 = n321 & n737;
  assign n745 = (n453 & n743) | (n453 & n744) | (n743 & n744);
  assign n534 = (n321 & n628) | (n321 & n745) | (n628 & n745);
  assign n746 = n321 | n738;
  assign n747 = n321 | n737;
  assign n748 = (n453 & n746) | (n453 & n747) | (n746 & n747);
  assign n536 = n628 | n748;
  assign n324 = ~n534 & n536;
  assign n538 = n281 & n324;
  assign n639 = (n283 & n324) | (n283 & n538) | (n324 & n538);
  assign n640 = (n507 & n538) | (n507 & n639) | (n538 & n639);
  assign n641 = (n233 & n538) | (n233 & n639) | (n538 & n639);
  assign n642 = (n493 & n640) | (n493 & n641) | (n640 & n641);
  assign n541 = n281 | n324;
  assign n643 = n283 | n541;
  assign n644 = (n507 & n541) | (n507 & n643) | (n541 & n643);
  assign n645 = (n233 & n541) | (n233 & n643) | (n541 & n643);
  assign n646 = (n493 & n644) | (n493 & n645) | (n644 & n645);
  assign n327 = ~n642 & n646;
  assign n328 = x6 & x12;
  assign n329 = n327 & n328;
  assign n330 = n327 | n328;
  assign n331 = ~n329 & n330;
  assign n529 = n288 | n290;
  assign n647 = n331 & n529;
  assign n648 = n288 & n331;
  assign n649 = (n506 & n647) | (n506 & n648) | (n647 & n648);
  assign n650 = n331 | n529;
  assign n651 = n288 | n331;
  assign n652 = (n506 & n650) | (n506 & n651) | (n650 & n651);
  assign n334 = ~n649 & n652;
  assign n335 = x5 & x13;
  assign n336 = n334 & n335;
  assign n337 = n334 | n335;
  assign n338 = ~n336 & n337;
  assign n339 = n528 & n338;
  assign n340 = n528 | n338;
  assign n341 = ~n339 & n340;
  assign n342 = x4 & x14;
  assign n343 = n341 & n342;
  assign n344 = n341 | n342;
  assign n345 = ~n343 & n344;
  assign n346 = n526 & n345;
  assign n347 = n526 | n345;
  assign n348 = ~n346 & n347;
  assign n349 = x3 & x15;
  assign n350 = n348 & n349;
  assign n351 = n348 | n349;
  assign n352 = ~n350 & n351;
  assign n353 = n524 & n352;
  assign n354 = n524 | n352;
  assign n355 = ~n353 & n354;
  assign n356 = n350 | n353;
  assign n361 = x7 & x12;
  assign n653 = n361 & n745;
  assign n654 = n321 & n361;
  assign n655 = (n628 & n653) | (n628 & n654) | (n653 & n654);
  assign n548 = (n361 & n642) | (n361 & n655) | (n642 & n655);
  assign n656 = n361 | n745;
  assign n657 = n321 | n361;
  assign n658 = (n628 & n656) | (n628 & n657) | (n656 & n657);
  assign n550 = n642 | n658;
  assign n364 = ~n548 & n550;
  assign n552 = n329 & n364;
  assign n659 = (n331 & n364) | (n331 & n552) | (n364 & n552);
  assign n660 = (n529 & n552) | (n529 & n659) | (n552 & n659);
  assign n661 = (n288 & n552) | (n288 & n659) | (n552 & n659);
  assign n662 = (n506 & n660) | (n506 & n661) | (n660 & n661);
  assign n555 = n329 | n364;
  assign n663 = n331 | n555;
  assign n664 = (n529 & n555) | (n529 & n663) | (n555 & n663);
  assign n665 = (n288 & n555) | (n288 & n663) | (n555 & n663);
  assign n666 = (n506 & n664) | (n506 & n665) | (n664 & n665);
  assign n367 = ~n662 & n666;
  assign n368 = x6 & x13;
  assign n369 = n367 & n368;
  assign n370 = n367 | n368;
  assign n371 = ~n369 & n370;
  assign n543 = n336 | n338;
  assign n667 = n371 & n543;
  assign n668 = n336 & n371;
  assign n669 = (n528 & n667) | (n528 & n668) | (n667 & n668);
  assign n670 = n371 | n543;
  assign n671 = n336 | n371;
  assign n672 = (n528 & n670) | (n528 & n671) | (n670 & n671);
  assign n374 = ~n669 & n672;
  assign n375 = x5 & x14;
  assign n376 = n374 & n375;
  assign n377 = n374 | n375;
  assign n378 = ~n376 & n377;
  assign n673 = n343 & n378;
  assign n674 = (n346 & n378) | (n346 & n673) | (n378 & n673);
  assign n675 = n343 | n378;
  assign n676 = n346 | n675;
  assign n381 = ~n674 & n676;
  assign n382 = x4 & x15;
  assign n383 = n381 & n382;
  assign n384 = n381 | n382;
  assign n385 = ~n383 & n384;
  assign n386 = n356 & n385;
  assign n387 = n356 | n385;
  assign n388 = ~n386 & n387;
  assign n677 = n383 | n385;
  assign n678 = (n356 & n383) | (n356 & n677) | (n383 & n677);
  assign n357 = n343 | n346;
  assign n393 = x7 & x13;
  assign n680 = n361 & n393;
  assign n2671 = n680 & n745;
  assign n750 = n393 & n654;
  assign n751 = (n628 & n2671) | (n628 & n750) | (n2671 & n750);
  assign n681 = (n642 & n751) | (n642 & n680) | (n751 & n680);
  assign n562 = (n393 & n662) | (n393 & n681) | (n662 & n681);
  assign n683 = n361 | n393;
  assign n2672 = (n393 & n683) | (n393 & n745) | (n683 & n745);
  assign n753 = n393 | n654;
  assign n754 = (n628 & n2672) | (n628 & n753) | (n2672 & n753);
  assign n684 = (n642 & n754) | (n642 & n683) | (n754 & n683);
  assign n564 = n662 | n684;
  assign n396 = ~n562 & n564;
  assign n566 = n369 & n396;
  assign n685 = (n371 & n396) | (n371 & n566) | (n396 & n566);
  assign n686 = (n543 & n566) | (n543 & n685) | (n566 & n685);
  assign n687 = (n336 & n566) | (n336 & n685) | (n566 & n685);
  assign n688 = (n528 & n686) | (n528 & n687) | (n686 & n687);
  assign n569 = n369 | n396;
  assign n689 = n371 | n569;
  assign n690 = (n543 & n569) | (n543 & n689) | (n569 & n689);
  assign n691 = (n336 & n569) | (n336 & n689) | (n569 & n689);
  assign n692 = (n528 & n690) | (n528 & n691) | (n690 & n691);
  assign n399 = ~n688 & n692;
  assign n400 = x6 & x14;
  assign n401 = n399 & n400;
  assign n402 = n399 | n400;
  assign n403 = ~n401 & n402;
  assign n557 = n376 | n378;
  assign n693 = n403 & n557;
  assign n694 = n376 & n403;
  assign n695 = (n357 & n693) | (n357 & n694) | (n693 & n694);
  assign n696 = n403 | n557;
  assign n697 = n376 | n403;
  assign n698 = (n357 & n696) | (n357 & n697) | (n696 & n697);
  assign n406 = ~n695 & n698;
  assign n407 = x5 & x15;
  assign n408 = n406 & n407;
  assign n409 = n406 | n407;
  assign n410 = ~n408 & n409;
  assign n411 = n678 & n410;
  assign n412 = n678 | n410;
  assign n413 = ~n411 & n412;
  assign n571 = n408 | n410;
  assign n572 = (n678 & n408) | (n678 & n571) | (n408 & n571);
  assign n417 = x7 & x14;
  assign n756 = n417 & n680;
  assign n3429 = n745 & n756;
  assign n700 = n393 & n417;
  assign n3430 = n654 & n700;
  assign n2675 = (n628 & n3429) | (n628 & n3430) | (n3429 & n3430);
  assign n757 = (n642 & n2675) | (n642 & n756) | (n2675 & n756);
  assign n701 = (n662 & n757) | (n662 & n700) | (n757 & n700);
  assign n576 = (n417 & n688) | (n417 & n701) | (n688 & n701);
  assign n759 = n417 | n680;
  assign n3431 = (n417 & n745) | (n417 & n759) | (n745 & n759);
  assign n703 = n393 | n417;
  assign n3432 = (n417 & n654) | (n417 & n703) | (n654 & n703);
  assign n2678 = (n628 & n3431) | (n628 & n3432) | (n3431 & n3432);
  assign n760 = (n642 & n2678) | (n642 & n759) | (n2678 & n759);
  assign n704 = (n662 & n760) | (n662 & n703) | (n760 & n703);
  assign n578 = n688 | n704;
  assign n420 = ~n576 & n578;
  assign n580 = n401 & n420;
  assign n705 = (n403 & n420) | (n403 & n580) | (n420 & n580);
  assign n706 = (n557 & n580) | (n557 & n705) | (n580 & n705);
  assign n707 = (n376 & n580) | (n376 & n705) | (n580 & n705);
  assign n708 = (n357 & n706) | (n357 & n707) | (n706 & n707);
  assign n583 = n401 | n420;
  assign n709 = n403 | n583;
  assign n710 = (n557 & n583) | (n557 & n709) | (n583 & n709);
  assign n711 = (n376 & n583) | (n376 & n709) | (n583 & n709);
  assign n712 = (n357 & n710) | (n357 & n711) | (n710 & n711);
  assign n423 = ~n708 & n712;
  assign n424 = x6 & x15;
  assign n425 = n423 & n424;
  assign n426 = n423 | n424;
  assign n427 = ~n425 & n426;
  assign n428 = n572 & n427;
  assign n429 = n572 | n427;
  assign n430 = ~n428 & n429;
  assign n433 = x7 & x15;
  assign n714 = n417 & n433;
  assign n3436 = n680 & n714;
  assign n3895 = n745 & n3436;
  assign n3434 = n433 & n3430;
  assign n3435 = (n628 & n3895) | (n628 & n3434) | (n3895 & n3434);
  assign n2681 = (n642 & n3435) | (n642 & n3436) | (n3435 & n3436);
  assign n762 = n433 & n700;
  assign n763 = (n662 & n2681) | (n662 & n762) | (n2681 & n762);
  assign n715 = (n688 & n763) | (n688 & n714) | (n763 & n714);
  assign n588 = (n433 & n708) | (n433 & n715) | (n708 & n715);
  assign n717 = n417 | n433;
  assign n3440 = (n433 & n680) | (n433 & n717) | (n680 & n717);
  assign n3896 = (n433 & n745) | (n433 & n3440) | (n745 & n3440);
  assign n3438 = n433 | n3430;
  assign n3439 = (n628 & n3896) | (n628 & n3438) | (n3896 & n3438);
  assign n2684 = (n642 & n3439) | (n642 & n3440) | (n3439 & n3440);
  assign n765 = n433 | n700;
  assign n766 = (n662 & n2684) | (n662 & n765) | (n2684 & n765);
  assign n718 = (n688 & n766) | (n688 & n717) | (n766 & n717);
  assign n590 = n708 | n718;
  assign n436 = ~n588 & n590;
  assign n592 = n425 & n436;
  assign n719 = (n427 & n436) | (n427 & n592) | (n436 & n592);
  assign n593 = (n572 & n719) | (n572 & n592) | (n719 & n592);
  assign n595 = n425 | n436;
  assign n720 = n427 | n595;
  assign n596 = (n572 & n720) | (n572 & n595) | (n720 & n595);
  assign n439 = ~n593 & n596;
  assign n721 = n588 | n719;
  assign n722 = n588 | n592;
  assign n723 = (n572 & n721) | (n572 & n722) | (n721 & n722);
  assign n799 = x16 & x32;
  assign n800 = x17 & x32;
  assign n801 = x16 & x33;
  assign n802 = n800 & n801;
  assign n803 = n800 | n801;
  assign n804 = ~n802 & n803;
  assign n805 = x18 & x32;
  assign n806 = x17 & x33;
  assign n807 = n805 & n806;
  assign n808 = n805 | n806;
  assign n809 = ~n807 & n808;
  assign n810 = n802 & n809;
  assign n811 = n802 | n809;
  assign n812 = ~n810 & n811;
  assign n813 = x16 & x34;
  assign n814 = n812 & n813;
  assign n815 = n812 | n813;
  assign n816 = ~n814 & n815;
  assign n2685 = n802 | n807;
  assign n2686 = (n807 & n809) | (n807 & n2685) | (n809 & n2685);
  assign n818 = x19 & x32;
  assign n819 = x18 & x33;
  assign n820 = n818 & n819;
  assign n821 = n818 | n819;
  assign n822 = ~n820 & n821;
  assign n823 = n2686 & n822;
  assign n824 = n2686 | n822;
  assign n825 = ~n823 & n824;
  assign n826 = x17 & x34;
  assign n827 = n825 & n826;
  assign n828 = n825 | n826;
  assign n829 = ~n827 & n828;
  assign n830 = n814 & n829;
  assign n831 = n814 | n829;
  assign n832 = ~n830 & n831;
  assign n833 = x16 & x35;
  assign n834 = n832 & n833;
  assign n835 = n832 | n833;
  assign n836 = ~n834 & n835;
  assign n2687 = n814 | n827;
  assign n2688 = (n827 & n829) | (n827 & n2687) | (n829 & n2687);
  assign n2689 = n820 | n822;
  assign n2690 = (n820 & n2686) | (n820 & n2689) | (n2686 & n2689);
  assign n839 = x20 & x32;
  assign n840 = x19 & x33;
  assign n841 = n839 & n840;
  assign n842 = n839 | n840;
  assign n843 = ~n841 & n842;
  assign n844 = n2690 & n843;
  assign n845 = n2690 | n843;
  assign n846 = ~n844 & n845;
  assign n847 = x18 & x34;
  assign n848 = n846 & n847;
  assign n849 = n846 | n847;
  assign n850 = ~n848 & n849;
  assign n851 = n2688 & n850;
  assign n852 = n2688 | n850;
  assign n853 = ~n851 & n852;
  assign n854 = x17 & x35;
  assign n855 = n853 & n854;
  assign n856 = n853 | n854;
  assign n857 = ~n855 & n856;
  assign n858 = n834 & n857;
  assign n859 = n834 | n857;
  assign n860 = ~n858 & n859;
  assign n861 = x16 & x36;
  assign n862 = n860 & n861;
  assign n863 = n860 | n861;
  assign n864 = ~n862 & n863;
  assign n2691 = n834 | n855;
  assign n2692 = (n855 & n857) | (n855 & n2691) | (n857 & n2691);
  assign n868 = x21 & x32;
  assign n869 = x20 & x33;
  assign n870 = n868 & n869;
  assign n871 = n868 | n869;
  assign n872 = ~n870 & n871;
  assign n2693 = n841 | n843;
  assign n2695 = n872 & n2693;
  assign n2696 = n841 & n872;
  assign n2697 = (n2690 & n2695) | (n2690 & n2696) | (n2695 & n2696);
  assign n2698 = n872 | n2693;
  assign n2699 = n841 | n872;
  assign n2700 = (n2690 & n2698) | (n2690 & n2699) | (n2698 & n2699);
  assign n875 = ~n2697 & n2700;
  assign n876 = x19 & x34;
  assign n877 = n875 & n876;
  assign n878 = n875 | n876;
  assign n879 = ~n877 & n878;
  assign n2701 = n848 & n879;
  assign n2702 = (n851 & n879) | (n851 & n2701) | (n879 & n2701);
  assign n2703 = n848 | n879;
  assign n2704 = n851 | n2703;
  assign n882 = ~n2702 & n2704;
  assign n883 = x18 & x35;
  assign n884 = n882 & n883;
  assign n885 = n882 | n883;
  assign n886 = ~n884 & n885;
  assign n887 = n2692 & n886;
  assign n888 = n2692 | n886;
  assign n889 = ~n887 & n888;
  assign n890 = x17 & x36;
  assign n891 = n889 & n890;
  assign n892 = n889 | n890;
  assign n893 = ~n891 & n892;
  assign n894 = n862 & n893;
  assign n895 = n862 | n893;
  assign n896 = ~n894 & n895;
  assign n897 = x16 & x37;
  assign n898 = n896 & n897;
  assign n899 = n896 | n897;
  assign n900 = ~n898 & n899;
  assign n2705 = n862 | n891;
  assign n2706 = (n891 & n893) | (n891 & n2705) | (n893 & n2705);
  assign n902 = n884 | n887;
  assign n905 = x22 & x32;
  assign n906 = x21 & x33;
  assign n907 = n905 & n906;
  assign n908 = n905 | n906;
  assign n909 = ~n907 & n908;
  assign n2707 = n870 & n909;
  assign n2708 = (n909 & n2697) | (n909 & n2707) | (n2697 & n2707);
  assign n2709 = n870 | n909;
  assign n2710 = n2697 | n2709;
  assign n912 = ~n2708 & n2710;
  assign n913 = x20 & x34;
  assign n914 = n912 & n913;
  assign n915 = n912 | n913;
  assign n916 = ~n914 & n915;
  assign n2711 = n877 & n916;
  assign n2712 = (n916 & n2702) | (n916 & n2711) | (n2702 & n2711);
  assign n2713 = n877 | n916;
  assign n2714 = n2702 | n2713;
  assign n919 = ~n2712 & n2714;
  assign n920 = x19 & x35;
  assign n921 = n919 & n920;
  assign n922 = n919 | n920;
  assign n923 = ~n921 & n922;
  assign n924 = n902 & n923;
  assign n925 = n902 | n923;
  assign n926 = ~n924 & n925;
  assign n927 = x18 & x36;
  assign n928 = n926 & n927;
  assign n929 = n926 | n927;
  assign n930 = ~n928 & n929;
  assign n931 = n2706 & n930;
  assign n932 = n2706 | n930;
  assign n933 = ~n931 & n932;
  assign n934 = x17 & x37;
  assign n935 = n933 & n934;
  assign n936 = n933 | n934;
  assign n937 = ~n935 & n936;
  assign n938 = n898 & n937;
  assign n939 = n898 | n937;
  assign n940 = ~n938 & n939;
  assign n941 = x16 & x38;
  assign n942 = n940 & n941;
  assign n943 = n940 | n941;
  assign n944 = ~n942 & n943;
  assign n3897 = n897 | n934;
  assign n3898 = (n896 & n934) | (n896 & n3897) | (n934 & n3897);
  assign n3442 = (n898 & n933) | (n898 & n3898) | (n933 & n3898);
  assign n2716 = (n935 & n937) | (n935 & n3442) | (n937 & n3442);
  assign n2717 = n928 | n2706;
  assign n2718 = (n928 & n930) | (n928 & n2717) | (n930 & n2717);
  assign n2719 = n921 | n923;
  assign n2720 = (n902 & n921) | (n902 & n2719) | (n921 & n2719);
  assign n950 = x23 & x32;
  assign n951 = x22 & x33;
  assign n952 = n950 & n951;
  assign n953 = n950 | n951;
  assign n954 = ~n952 & n953;
  assign n3443 = n870 | n907;
  assign n3444 = (n907 & n909) | (n907 & n3443) | (n909 & n3443);
  assign n2724 = n954 & n3444;
  assign n2722 = n907 | n909;
  assign n2725 = n954 & n2722;
  assign n2726 = (n2697 & n2724) | (n2697 & n2725) | (n2724 & n2725);
  assign n2727 = n954 | n3444;
  assign n2728 = n954 | n2722;
  assign n2729 = (n2697 & n2727) | (n2697 & n2728) | (n2727 & n2728);
  assign n957 = ~n2726 & n2729;
  assign n958 = x21 & x34;
  assign n959 = n957 & n958;
  assign n960 = n957 | n958;
  assign n961 = ~n959 & n960;
  assign n2730 = n914 & n961;
  assign n2731 = (n961 & n2712) | (n961 & n2730) | (n2712 & n2730);
  assign n2732 = n914 | n961;
  assign n2733 = n2712 | n2732;
  assign n964 = ~n2731 & n2733;
  assign n965 = x20 & x35;
  assign n966 = n964 & n965;
  assign n967 = n964 | n965;
  assign n968 = ~n966 & n967;
  assign n969 = n2720 & n968;
  assign n970 = n2720 | n968;
  assign n971 = ~n969 & n970;
  assign n972 = x19 & x36;
  assign n973 = n971 & n972;
  assign n974 = n971 | n972;
  assign n975 = ~n973 & n974;
  assign n976 = n2718 & n975;
  assign n977 = n2718 | n975;
  assign n978 = ~n976 & n977;
  assign n979 = x18 & x37;
  assign n980 = n978 & n979;
  assign n981 = n978 | n979;
  assign n982 = ~n980 & n981;
  assign n983 = n2716 & n982;
  assign n984 = n2716 | n982;
  assign n985 = ~n983 & n984;
  assign n986 = x17 & x38;
  assign n987 = n985 & n986;
  assign n988 = n985 | n986;
  assign n989 = ~n987 & n988;
  assign n990 = n942 & n989;
  assign n991 = n942 | n989;
  assign n992 = ~n990 & n991;
  assign n993 = x16 & x39;
  assign n994 = n992 & n993;
  assign n995 = n992 | n993;
  assign n996 = ~n994 & n995;
  assign n2734 = n942 | n987;
  assign n2735 = (n987 & n989) | (n987 & n2734) | (n989 & n2734);
  assign n998 = n980 | n983;
  assign n999 = n973 | n976;
  assign n2736 = n966 | n968;
  assign n2737 = (n966 & n2720) | (n966 & n2736) | (n2720 & n2736);
  assign n1003 = x24 & x32;
  assign n1004 = x23 & x33;
  assign n1005 = n1003 & n1004;
  assign n1006 = n1003 | n1004;
  assign n1007 = ~n1005 & n1006;
  assign n2741 = n952 & n1007;
  assign n3447 = (n1007 & n2725) | (n1007 & n2741) | (n2725 & n2741);
  assign n3448 = (n1007 & n2724) | (n1007 & n2741) | (n2724 & n2741);
  assign n3449 = (n2697 & n3447) | (n2697 & n3448) | (n3447 & n3448);
  assign n2743 = n952 | n1007;
  assign n3450 = n2725 | n2743;
  assign n3451 = n2724 | n2743;
  assign n3452 = (n2697 & n3450) | (n2697 & n3451) | (n3450 & n3451);
  assign n1010 = ~n3449 & n3452;
  assign n1011 = x22 & x34;
  assign n1012 = n1010 & n1011;
  assign n1013 = n1010 | n1011;
  assign n1014 = ~n1012 & n1013;
  assign n2739 = n959 | n961;
  assign n3453 = n1014 & n2739;
  assign n3445 = n914 | n959;
  assign n3446 = (n959 & n961) | (n959 & n3445) | (n961 & n3445);
  assign n3454 = n1014 & n3446;
  assign n3455 = (n2712 & n3453) | (n2712 & n3454) | (n3453 & n3454);
  assign n3456 = n1014 | n2739;
  assign n3457 = n1014 | n3446;
  assign n3458 = (n2712 & n3456) | (n2712 & n3457) | (n3456 & n3457);
  assign n1017 = ~n3455 & n3458;
  assign n1018 = x21 & x35;
  assign n1019 = n1017 & n1018;
  assign n1020 = n1017 | n1018;
  assign n1021 = ~n1019 & n1020;
  assign n1022 = n2737 & n1021;
  assign n1023 = n2737 | n1021;
  assign n1024 = ~n1022 & n1023;
  assign n1025 = x20 & x36;
  assign n1026 = n1024 & n1025;
  assign n1027 = n1024 | n1025;
  assign n1028 = ~n1026 & n1027;
  assign n1029 = n999 & n1028;
  assign n1030 = n999 | n1028;
  assign n1031 = ~n1029 & n1030;
  assign n1032 = x19 & x37;
  assign n1033 = n1031 & n1032;
  assign n1034 = n1031 | n1032;
  assign n1035 = ~n1033 & n1034;
  assign n1036 = n998 & n1035;
  assign n1037 = n998 | n1035;
  assign n1038 = ~n1036 & n1037;
  assign n1039 = x18 & x38;
  assign n1040 = n1038 & n1039;
  assign n1041 = n1038 | n1039;
  assign n1042 = ~n1040 & n1041;
  assign n1043 = n2735 & n1042;
  assign n1044 = n2735 | n1042;
  assign n1045 = ~n1043 & n1044;
  assign n1046 = x17 & x39;
  assign n1047 = n1045 & n1046;
  assign n1048 = n1045 | n1046;
  assign n1049 = ~n1047 & n1048;
  assign n1050 = n994 & n1049;
  assign n1051 = n994 | n1049;
  assign n1052 = ~n1050 & n1051;
  assign n1053 = x16 & x40;
  assign n1054 = n1052 & n1053;
  assign n1055 = n1052 | n1053;
  assign n1056 = ~n1054 & n1055;
  assign n3899 = n993 | n1046;
  assign n3900 = (n992 & n1046) | (n992 & n3899) | (n1046 & n3899);
  assign n3460 = (n994 & n1045) | (n994 & n3900) | (n1045 & n3900);
  assign n2746 = (n1047 & n1049) | (n1047 & n3460) | (n1049 & n3460);
  assign n2747 = n1040 | n2735;
  assign n2748 = (n1040 & n1042) | (n1040 & n2747) | (n1042 & n2747);
  assign n1059 = n1033 | n1036;
  assign n2749 = n1026 | n1028;
  assign n2750 = (n999 & n1026) | (n999 & n2749) | (n1026 & n2749);
  assign n2740 = (n2712 & n3446) | (n2712 & n2739) | (n3446 & n2739);
  assign n1064 = x25 & x32;
  assign n1065 = x24 & x33;
  assign n1066 = n1064 & n1065;
  assign n1067 = n1064 | n1065;
  assign n1068 = ~n1066 & n1067;
  assign n3461 = n952 | n1005;
  assign n3462 = (n1005 & n1007) | (n1005 & n3461) | (n1007 & n3461);
  assign n2758 = n1068 & n3462;
  assign n2756 = n1005 | n1007;
  assign n2759 = n1068 & n2756;
  assign n3463 = (n2725 & n2758) | (n2725 & n2759) | (n2758 & n2759);
  assign n3464 = (n2724 & n2758) | (n2724 & n2759) | (n2758 & n2759);
  assign n3465 = (n2697 & n3463) | (n2697 & n3464) | (n3463 & n3464);
  assign n2761 = n1068 | n3462;
  assign n2762 = n1068 | n2756;
  assign n3466 = (n2725 & n2761) | (n2725 & n2762) | (n2761 & n2762);
  assign n3467 = (n2724 & n2761) | (n2724 & n2762) | (n2761 & n2762);
  assign n3468 = (n2697 & n3466) | (n2697 & n3467) | (n3466 & n3467);
  assign n1071 = ~n3465 & n3468;
  assign n1072 = x23 & x34;
  assign n1073 = n1071 & n1072;
  assign n1074 = n1071 | n1072;
  assign n1075 = ~n1073 & n1074;
  assign n2753 = n1012 | n1014;
  assign n2764 = n1075 & n2753;
  assign n2765 = n1012 & n1075;
  assign n2766 = (n2740 & n2764) | (n2740 & n2765) | (n2764 & n2765);
  assign n2767 = n1075 | n2753;
  assign n2768 = n1012 | n1075;
  assign n2769 = (n2740 & n2767) | (n2740 & n2768) | (n2767 & n2768);
  assign n1078 = ~n2766 & n2769;
  assign n1079 = x22 & x35;
  assign n1080 = n1078 & n1079;
  assign n1081 = n1078 | n1079;
  assign n1082 = ~n1080 & n1081;
  assign n2751 = n1019 | n1021;
  assign n3469 = n1082 & n2751;
  assign n3470 = n1019 & n1082;
  assign n3471 = (n2737 & n3469) | (n2737 & n3470) | (n3469 & n3470);
  assign n3472 = n1082 | n2751;
  assign n3473 = n1019 | n1082;
  assign n3474 = (n2737 & n3472) | (n2737 & n3473) | (n3472 & n3473);
  assign n1085 = ~n3471 & n3474;
  assign n1086 = x21 & x36;
  assign n1087 = n1085 & n1086;
  assign n1088 = n1085 | n1086;
  assign n1089 = ~n1087 & n1088;
  assign n1090 = n2750 & n1089;
  assign n1091 = n2750 | n1089;
  assign n1092 = ~n1090 & n1091;
  assign n1093 = x20 & x37;
  assign n1094 = n1092 & n1093;
  assign n1095 = n1092 | n1093;
  assign n1096 = ~n1094 & n1095;
  assign n1097 = n1059 & n1096;
  assign n1098 = n1059 | n1096;
  assign n1099 = ~n1097 & n1098;
  assign n1100 = x19 & x38;
  assign n1101 = n1099 & n1100;
  assign n1102 = n1099 | n1100;
  assign n1103 = ~n1101 & n1102;
  assign n1104 = n2748 & n1103;
  assign n1105 = n2748 | n1103;
  assign n1106 = ~n1104 & n1105;
  assign n1107 = x18 & x39;
  assign n1108 = n1106 & n1107;
  assign n1109 = n1106 | n1107;
  assign n1110 = ~n1108 & n1109;
  assign n1111 = n2746 & n1110;
  assign n1112 = n2746 | n1110;
  assign n1113 = ~n1111 & n1112;
  assign n1114 = x17 & x40;
  assign n1115 = n1113 & n1114;
  assign n1116 = n1113 | n1114;
  assign n1117 = ~n1115 & n1116;
  assign n1118 = n1054 & n1117;
  assign n1119 = n1054 | n1117;
  assign n1120 = ~n1118 & n1119;
  assign n1121 = x16 & x41;
  assign n1122 = n1120 & n1121;
  assign n1123 = n1120 | n1121;
  assign n1124 = ~n1122 & n1123;
  assign n3901 = n1053 | n1114;
  assign n3902 = (n1052 & n1114) | (n1052 & n3901) | (n1114 & n3901);
  assign n3476 = (n1054 & n1113) | (n1054 & n3902) | (n1113 & n3902);
  assign n2771 = (n1115 & n1117) | (n1115 & n3476) | (n1117 & n3476);
  assign n2772 = n1108 | n2746;
  assign n2773 = (n1108 & n1110) | (n1108 & n2772) | (n1110 & n2772);
  assign n2774 = n1101 | n2748;
  assign n2775 = (n1101 & n1103) | (n1101 & n2774) | (n1103 & n2774);
  assign n2776 = n1094 | n1096;
  assign n2777 = (n1059 & n1094) | (n1059 & n2776) | (n1094 & n2776);
  assign n2752 = (n1019 & n2737) | (n1019 & n2751) | (n2737 & n2751);
  assign n3477 = n1066 | n1068;
  assign n3478 = (n1066 & n3462) | (n1066 & n3477) | (n3462 & n3477);
  assign n3479 = (n1066 & n2756) | (n1066 & n3477) | (n2756 & n3477);
  assign n3480 = (n2725 & n3478) | (n2725 & n3479) | (n3478 & n3479);
  assign n3481 = (n2724 & n3478) | (n2724 & n3479) | (n3478 & n3479);
  assign n3482 = (n2697 & n3480) | (n2697 & n3481) | (n3480 & n3481);
  assign n1133 = x26 & x32;
  assign n1134 = x25 & x33;
  assign n1135 = n1133 & n1134;
  assign n1136 = n1133 | n1134;
  assign n1137 = ~n1135 & n1136;
  assign n1138 = n3482 & n1137;
  assign n1139 = n3482 | n1137;
  assign n1140 = ~n1138 & n1139;
  assign n1141 = x24 & x34;
  assign n1142 = n1140 & n1141;
  assign n1143 = n1140 | n1141;
  assign n1144 = ~n1142 & n1143;
  assign n2785 = n1073 & n1144;
  assign n3483 = (n1144 & n2764) | (n1144 & n2785) | (n2764 & n2785);
  assign n3484 = (n1144 & n2765) | (n1144 & n2785) | (n2765 & n2785);
  assign n3485 = (n2740 & n3483) | (n2740 & n3484) | (n3483 & n3484);
  assign n2787 = n1073 | n1144;
  assign n3486 = n2764 | n2787;
  assign n3487 = n2765 | n2787;
  assign n3488 = (n2740 & n3486) | (n2740 & n3487) | (n3486 & n3487);
  assign n1147 = ~n3485 & n3488;
  assign n1148 = x23 & x35;
  assign n1149 = n1147 & n1148;
  assign n1150 = n1147 | n1148;
  assign n1151 = ~n1149 & n1150;
  assign n2780 = n1080 | n1082;
  assign n2789 = n1151 & n2780;
  assign n2790 = n1080 & n1151;
  assign n2791 = (n2752 & n2789) | (n2752 & n2790) | (n2789 & n2790);
  assign n2792 = n1151 | n2780;
  assign n2793 = n1080 | n1151;
  assign n2794 = (n2752 & n2792) | (n2752 & n2793) | (n2792 & n2793);
  assign n1154 = ~n2791 & n2794;
  assign n1155 = x22 & x36;
  assign n1156 = n1154 & n1155;
  assign n1157 = n1154 | n1155;
  assign n1158 = ~n1156 & n1157;
  assign n2778 = n1087 | n1089;
  assign n3489 = n1158 & n2778;
  assign n3490 = n1087 & n1158;
  assign n3491 = (n2750 & n3489) | (n2750 & n3490) | (n3489 & n3490);
  assign n3492 = n1158 | n2778;
  assign n3493 = n1087 | n1158;
  assign n3494 = (n2750 & n3492) | (n2750 & n3493) | (n3492 & n3493);
  assign n1161 = ~n3491 & n3494;
  assign n1162 = x21 & x37;
  assign n1163 = n1161 & n1162;
  assign n1164 = n1161 | n1162;
  assign n1165 = ~n1163 & n1164;
  assign n1166 = n2777 & n1165;
  assign n1167 = n2777 | n1165;
  assign n1168 = ~n1166 & n1167;
  assign n1169 = x20 & x38;
  assign n1170 = n1168 & n1169;
  assign n1171 = n1168 | n1169;
  assign n1172 = ~n1170 & n1171;
  assign n1173 = n2775 & n1172;
  assign n1174 = n2775 | n1172;
  assign n1175 = ~n1173 & n1174;
  assign n1176 = x19 & x39;
  assign n1177 = n1175 & n1176;
  assign n1178 = n1175 | n1176;
  assign n1179 = ~n1177 & n1178;
  assign n1180 = n2773 & n1179;
  assign n1181 = n2773 | n1179;
  assign n1182 = ~n1180 & n1181;
  assign n1183 = x18 & x40;
  assign n1184 = n1182 & n1183;
  assign n1185 = n1182 | n1183;
  assign n1186 = ~n1184 & n1185;
  assign n1187 = n2771 & n1186;
  assign n1188 = n2771 | n1186;
  assign n1189 = ~n1187 & n1188;
  assign n1190 = x17 & x41;
  assign n1191 = n1189 & n1190;
  assign n1192 = n1189 | n1190;
  assign n1193 = ~n1191 & n1192;
  assign n1194 = n1122 & n1193;
  assign n1195 = n1122 | n1193;
  assign n1196 = ~n1194 & n1195;
  assign n1197 = x16 & x42;
  assign n1198 = n1196 & n1197;
  assign n1199 = n1196 | n1197;
  assign n1200 = ~n1198 & n1199;
  assign n2795 = n1122 | n1191;
  assign n2796 = (n1191 & n1193) | (n1191 & n2795) | (n1193 & n2795);
  assign n1202 = n1184 | n1187;
  assign n1203 = n1177 | n1180;
  assign n2779 = (n1087 & n2750) | (n1087 & n2778) | (n2750 & n2778);
  assign n2802 = n1142 | n1144;
  assign n3495 = n1073 | n1142;
  assign n3496 = (n1142 & n1144) | (n1142 & n3495) | (n1144 & n3495);
  assign n3497 = (n2764 & n2802) | (n2764 & n3496) | (n2802 & n3496);
  assign n3498 = (n2765 & n2802) | (n2765 & n3496) | (n2802 & n3496);
  assign n3499 = (n2740 & n3497) | (n2740 & n3498) | (n3497 & n3498);
  assign n1210 = x27 & x32;
  assign n1211 = x26 & x33;
  assign n1212 = n1210 & n1211;
  assign n1213 = n1210 | n1211;
  assign n1214 = ~n1212 & n1213;
  assign n2804 = n1135 | n1137;
  assign n2806 = n1214 & n2804;
  assign n2807 = n1135 & n1214;
  assign n2808 = (n3482 & n2806) | (n3482 & n2807) | (n2806 & n2807);
  assign n2809 = n1214 | n2804;
  assign n2810 = n1135 | n1214;
  assign n2811 = (n3482 & n2809) | (n3482 & n2810) | (n2809 & n2810);
  assign n1217 = ~n2808 & n2811;
  assign n1218 = x25 & x34;
  assign n1219 = n1217 & n1218;
  assign n1220 = n1217 | n1218;
  assign n1221 = ~n1219 & n1220;
  assign n1222 = n3499 & n1221;
  assign n1223 = n3499 | n1221;
  assign n1224 = ~n1222 & n1223;
  assign n1225 = x24 & x35;
  assign n1226 = n1224 & n1225;
  assign n1227 = n1224 | n1225;
  assign n1228 = ~n1226 & n1227;
  assign n2812 = n1149 & n1228;
  assign n2813 = (n1228 & n2791) | (n1228 & n2812) | (n2791 & n2812);
  assign n2814 = n1149 | n1228;
  assign n2815 = n2791 | n2814;
  assign n1231 = ~n2813 & n2815;
  assign n1232 = x23 & x36;
  assign n1233 = n1231 & n1232;
  assign n1234 = n1231 | n1232;
  assign n1235 = ~n1233 & n1234;
  assign n2799 = n1156 | n1158;
  assign n2816 = n1235 & n2799;
  assign n2817 = n1156 & n1235;
  assign n2818 = (n2779 & n2816) | (n2779 & n2817) | (n2816 & n2817);
  assign n2819 = n1235 | n2799;
  assign n2820 = n1156 | n1235;
  assign n2821 = (n2779 & n2819) | (n2779 & n2820) | (n2819 & n2820);
  assign n1238 = ~n2818 & n2821;
  assign n1239 = x22 & x37;
  assign n1240 = n1238 & n1239;
  assign n1241 = n1238 | n1239;
  assign n1242 = ~n1240 & n1241;
  assign n2797 = n1163 | n1165;
  assign n3500 = n1242 & n2797;
  assign n3501 = n1163 & n1242;
  assign n3502 = (n2777 & n3500) | (n2777 & n3501) | (n3500 & n3501);
  assign n3503 = n1242 | n2797;
  assign n3504 = n1163 | n1242;
  assign n3505 = (n2777 & n3503) | (n2777 & n3504) | (n3503 & n3504);
  assign n1245 = ~n3502 & n3505;
  assign n1246 = x21 & x38;
  assign n1247 = n1245 & n1246;
  assign n1248 = n1245 | n1246;
  assign n1249 = ~n1247 & n1248;
  assign n3506 = n1170 & n1249;
  assign n3507 = (n1173 & n1249) | (n1173 & n3506) | (n1249 & n3506);
  assign n3508 = n1170 | n1249;
  assign n3509 = n1173 | n3508;
  assign n1252 = ~n3507 & n3509;
  assign n1253 = x20 & x39;
  assign n1254 = n1252 & n1253;
  assign n1255 = n1252 | n1253;
  assign n1256 = ~n1254 & n1255;
  assign n1257 = n1203 & n1256;
  assign n1258 = n1203 | n1256;
  assign n1259 = ~n1257 & n1258;
  assign n1260 = x19 & x40;
  assign n1261 = n1259 & n1260;
  assign n1262 = n1259 | n1260;
  assign n1263 = ~n1261 & n1262;
  assign n1264 = n1202 & n1263;
  assign n1265 = n1202 | n1263;
  assign n1266 = ~n1264 & n1265;
  assign n1267 = x18 & x41;
  assign n1268 = n1266 & n1267;
  assign n1269 = n1266 | n1267;
  assign n1270 = ~n1268 & n1269;
  assign n1271 = n2796 & n1270;
  assign n1272 = n2796 | n1270;
  assign n1273 = ~n1271 & n1272;
  assign n1274 = x17 & x42;
  assign n1275 = n1273 & n1274;
  assign n1276 = n1273 | n1274;
  assign n1277 = ~n1275 & n1276;
  assign n1278 = n1198 & n1277;
  assign n1279 = n1198 | n1277;
  assign n1280 = ~n1278 & n1279;
  assign n1281 = x16 & x43;
  assign n1282 = n1280 & n1281;
  assign n1283 = n1280 | n1281;
  assign n1284 = ~n1282 & n1283;
  assign n3903 = n1197 | n1274;
  assign n3904 = (n1196 & n1274) | (n1196 & n3903) | (n1274 & n3903);
  assign n3511 = (n1198 & n1273) | (n1198 & n3904) | (n1273 & n3904);
  assign n2823 = (n1275 & n1277) | (n1275 & n3511) | (n1277 & n3511);
  assign n2824 = n1268 | n2796;
  assign n2825 = (n1268 & n1270) | (n1268 & n2824) | (n1270 & n2824);
  assign n1287 = n1261 | n1264;
  assign n3512 = n1254 | n1256;
  assign n3513 = (n1203 & n1254) | (n1203 & n3512) | (n1254 & n3512);
  assign n1204 = n1170 | n1173;
  assign n2798 = (n1163 & n2777) | (n1163 & n2797) | (n2777 & n2797);
  assign n1295 = x28 & x32;
  assign n1296 = x27 & x33;
  assign n1297 = n1295 & n1296;
  assign n1298 = n1295 | n1296;
  assign n1299 = ~n1297 & n1298;
  assign n3514 = n1212 | n1214;
  assign n3515 = (n1212 & n2804) | (n1212 & n3514) | (n2804 & n3514);
  assign n2835 = n1299 & n3515;
  assign n3516 = n1135 | n1212;
  assign n3517 = (n1212 & n1214) | (n1212 & n3516) | (n1214 & n3516);
  assign n2836 = n1299 & n3517;
  assign n2837 = (n3482 & n2835) | (n3482 & n2836) | (n2835 & n2836);
  assign n2838 = n1299 | n3515;
  assign n2839 = n1299 | n3517;
  assign n2840 = (n3482 & n2838) | (n3482 & n2839) | (n2838 & n2839);
  assign n1302 = ~n2837 & n2840;
  assign n1303 = x26 & x34;
  assign n1304 = n1302 & n1303;
  assign n1305 = n1302 | n1303;
  assign n1306 = ~n1304 & n1305;
  assign n2830 = n1219 | n1221;
  assign n2841 = n1306 & n2830;
  assign n2842 = n1219 & n1306;
  assign n2843 = (n3499 & n2841) | (n3499 & n2842) | (n2841 & n2842);
  assign n2844 = n1306 | n2830;
  assign n2845 = n1219 | n1306;
  assign n2846 = (n3499 & n2844) | (n3499 & n2845) | (n2844 & n2845);
  assign n1309 = ~n2843 & n2846;
  assign n1310 = x25 & x35;
  assign n1311 = n1309 & n1310;
  assign n1312 = n1309 | n1310;
  assign n1313 = ~n1311 & n1312;
  assign n2847 = n1226 & n1313;
  assign n3518 = (n1313 & n2812) | (n1313 & n2847) | (n2812 & n2847);
  assign n3519 = (n1228 & n1313) | (n1228 & n2847) | (n1313 & n2847);
  assign n3520 = (n2791 & n3518) | (n2791 & n3519) | (n3518 & n3519);
  assign n2849 = n1226 | n1313;
  assign n3521 = n2812 | n2849;
  assign n3522 = n1228 | n2849;
  assign n3523 = (n2791 & n3521) | (n2791 & n3522) | (n3521 & n3522);
  assign n1316 = ~n3520 & n3523;
  assign n1317 = x24 & x36;
  assign n1318 = n1316 & n1317;
  assign n1319 = n1316 | n1317;
  assign n1320 = ~n1318 & n1319;
  assign n2851 = n1233 & n1320;
  assign n2852 = (n1320 & n2818) | (n1320 & n2851) | (n2818 & n2851);
  assign n2853 = n1233 | n1320;
  assign n2854 = n2818 | n2853;
  assign n1323 = ~n2852 & n2854;
  assign n1324 = x23 & x37;
  assign n1325 = n1323 & n1324;
  assign n1326 = n1323 | n1324;
  assign n1327 = ~n1325 & n1326;
  assign n2828 = n1240 | n1242;
  assign n2855 = n1327 & n2828;
  assign n2856 = n1240 & n1327;
  assign n2857 = (n2798 & n2855) | (n2798 & n2856) | (n2855 & n2856);
  assign n2858 = n1327 | n2828;
  assign n2859 = n1240 | n1327;
  assign n2860 = (n2798 & n2858) | (n2798 & n2859) | (n2858 & n2859);
  assign n1330 = ~n2857 & n2860;
  assign n1331 = x22 & x38;
  assign n1332 = n1330 & n1331;
  assign n1333 = n1330 | n1331;
  assign n1334 = ~n1332 & n1333;
  assign n2826 = n1247 | n1249;
  assign n3524 = n1334 & n2826;
  assign n3525 = n1247 & n1334;
  assign n3526 = (n1204 & n3524) | (n1204 & n3525) | (n3524 & n3525);
  assign n3527 = n1334 | n2826;
  assign n3528 = n1247 | n1334;
  assign n3529 = (n1204 & n3527) | (n1204 & n3528) | (n3527 & n3528);
  assign n1337 = ~n3526 & n3529;
  assign n1338 = x21 & x39;
  assign n1339 = n1337 & n1338;
  assign n1340 = n1337 | n1338;
  assign n1341 = ~n1339 & n1340;
  assign n1342 = n3513 & n1341;
  assign n1343 = n3513 | n1341;
  assign n1344 = ~n1342 & n1343;
  assign n1345 = x20 & x40;
  assign n1346 = n1344 & n1345;
  assign n1347 = n1344 | n1345;
  assign n1348 = ~n1346 & n1347;
  assign n1349 = n1287 & n1348;
  assign n1350 = n1287 | n1348;
  assign n1351 = ~n1349 & n1350;
  assign n1352 = x19 & x41;
  assign n1353 = n1351 & n1352;
  assign n1354 = n1351 | n1352;
  assign n1355 = ~n1353 & n1354;
  assign n1356 = n2825 & n1355;
  assign n1357 = n2825 | n1355;
  assign n1358 = ~n1356 & n1357;
  assign n1359 = x18 & x42;
  assign n1360 = n1358 & n1359;
  assign n1361 = n1358 | n1359;
  assign n1362 = ~n1360 & n1361;
  assign n1363 = n2823 & n1362;
  assign n1364 = n2823 | n1362;
  assign n1365 = ~n1363 & n1364;
  assign n1366 = x17 & x43;
  assign n1367 = n1365 & n1366;
  assign n1368 = n1365 | n1366;
  assign n1369 = ~n1367 & n1368;
  assign n1370 = n1282 & n1369;
  assign n1371 = n1282 | n1369;
  assign n1372 = ~n1370 & n1371;
  assign n1373 = x16 & x44;
  assign n1374 = n1372 & n1373;
  assign n1375 = n1372 | n1373;
  assign n1376 = ~n1374 & n1375;
  assign n3905 = n1281 | n1366;
  assign n3906 = (n1280 & n1366) | (n1280 & n3905) | (n1366 & n3905);
  assign n3531 = (n1282 & n1365) | (n1282 & n3906) | (n1365 & n3906);
  assign n2862 = (n1367 & n1369) | (n1367 & n3531) | (n1369 & n3531);
  assign n2863 = n1360 | n2823;
  assign n2864 = (n1360 & n1362) | (n1360 & n2863) | (n1362 & n2863);
  assign n2865 = n1353 | n2825;
  assign n2866 = (n1353 & n1355) | (n1353 & n2865) | (n1355 & n2865);
  assign n3532 = n1346 | n1348;
  assign n3533 = (n1287 & n1346) | (n1287 & n3532) | (n1346 & n3532);
  assign n2867 = n1339 | n1341;
  assign n2868 = (n3513 & n1339) | (n3513 & n2867) | (n1339 & n2867);
  assign n2827 = (n1204 & n1247) | (n1204 & n2826) | (n1247 & n2826);
  assign n2872 = n1311 | n1313;
  assign n3534 = n1226 | n1311;
  assign n3535 = (n1311 & n1313) | (n1311 & n3534) | (n1313 & n3534);
  assign n3536 = (n2812 & n2872) | (n2812 & n3535) | (n2872 & n3535);
  assign n3537 = (n1228 & n2872) | (n1228 & n3535) | (n2872 & n3535);
  assign n3538 = (n2791 & n3536) | (n2791 & n3537) | (n3536 & n3537);
  assign n1388 = x29 & x32;
  assign n1389 = x28 & x33;
  assign n1390 = n1388 & n1389;
  assign n1391 = n1388 | n1389;
  assign n1392 = ~n1390 & n1391;
  assign n3543 = n1297 | n1299;
  assign n3907 = n1392 & n3543;
  assign n3908 = n1297 & n1392;
  assign n3909 = (n3515 & n3907) | (n3515 & n3908) | (n3907 & n3908);
  assign n3545 = (n1297 & n3517) | (n1297 & n3543) | (n3517 & n3543);
  assign n3547 = n1392 & n3545;
  assign n3548 = (n3482 & n3909) | (n3482 & n3547) | (n3909 & n3547);
  assign n3910 = n1392 | n3543;
  assign n3911 = n1297 | n1392;
  assign n3912 = (n3515 & n3910) | (n3515 & n3911) | (n3910 & n3911);
  assign n3550 = n1392 | n3545;
  assign n3551 = (n3482 & n3912) | (n3482 & n3550) | (n3912 & n3550);
  assign n1395 = ~n3548 & n3551;
  assign n1396 = x27 & x34;
  assign n1397 = n1395 & n1396;
  assign n1398 = n1395 | n1396;
  assign n1399 = ~n1397 & n1398;
  assign n3539 = n1304 | n1306;
  assign n3540 = (n1304 & n2830) | (n1304 & n3539) | (n2830 & n3539);
  assign n3552 = n1399 & n3540;
  assign n3541 = n1219 | n1304;
  assign n3542 = (n1304 & n1306) | (n1304 & n3541) | (n1306 & n3541);
  assign n3553 = n1399 & n3542;
  assign n3554 = (n3499 & n3552) | (n3499 & n3553) | (n3552 & n3553);
  assign n3555 = n1399 | n3540;
  assign n3556 = n1399 | n3542;
  assign n3557 = (n3499 & n3555) | (n3499 & n3556) | (n3555 & n3556);
  assign n1402 = ~n3554 & n3557;
  assign n1403 = x26 & x35;
  assign n1404 = n1402 & n1403;
  assign n1405 = n1402 | n1403;
  assign n1406 = ~n1404 & n1405;
  assign n1407 = n3538 & n1406;
  assign n1408 = n3538 | n1406;
  assign n1409 = ~n1407 & n1408;
  assign n1410 = x25 & x36;
  assign n1411 = n1409 & n1410;
  assign n1412 = n1409 | n1410;
  assign n1413 = ~n1411 & n1412;
  assign n2880 = n1318 & n1413;
  assign n2881 = (n1413 & n2852) | (n1413 & n2880) | (n2852 & n2880);
  assign n2882 = n1318 | n1413;
  assign n2883 = n2852 | n2882;
  assign n1416 = ~n2881 & n2883;
  assign n1417 = x24 & x37;
  assign n1418 = n1416 & n1417;
  assign n1419 = n1416 | n1417;
  assign n1420 = ~n1418 & n1419;
  assign n2884 = n1325 & n1420;
  assign n2885 = (n1420 & n2857) | (n1420 & n2884) | (n2857 & n2884);
  assign n2886 = n1325 | n1420;
  assign n2887 = n2857 | n2886;
  assign n1423 = ~n2885 & n2887;
  assign n1424 = x23 & x38;
  assign n1425 = n1423 & n1424;
  assign n1426 = n1423 | n1424;
  assign n1427 = ~n1425 & n1426;
  assign n2869 = n1332 | n1334;
  assign n2888 = n1427 & n2869;
  assign n2889 = n1332 & n1427;
  assign n2890 = (n2827 & n2888) | (n2827 & n2889) | (n2888 & n2889);
  assign n2891 = n1427 | n2869;
  assign n2892 = n1332 | n1427;
  assign n2893 = (n2827 & n2891) | (n2827 & n2892) | (n2891 & n2892);
  assign n1430 = ~n2890 & n2893;
  assign n1431 = x22 & x39;
  assign n1432 = n1430 & n1431;
  assign n1433 = n1430 | n1431;
  assign n1434 = ~n1432 & n1433;
  assign n1435 = n2868 & n1434;
  assign n1436 = n2868 | n1434;
  assign n1437 = ~n1435 & n1436;
  assign n1438 = x21 & x40;
  assign n1439 = n1437 & n1438;
  assign n1440 = n1437 | n1438;
  assign n1441 = ~n1439 & n1440;
  assign n1442 = n3533 & n1441;
  assign n1443 = n3533 | n1441;
  assign n1444 = ~n1442 & n1443;
  assign n1445 = x20 & x41;
  assign n1446 = n1444 & n1445;
  assign n1447 = n1444 | n1445;
  assign n1448 = ~n1446 & n1447;
  assign n1449 = n2866 & n1448;
  assign n1450 = n2866 | n1448;
  assign n1451 = ~n1449 & n1450;
  assign n1452 = x19 & x42;
  assign n1453 = n1451 & n1452;
  assign n1454 = n1451 | n1452;
  assign n1455 = ~n1453 & n1454;
  assign n1456 = n2864 & n1455;
  assign n1457 = n2864 | n1455;
  assign n1458 = ~n1456 & n1457;
  assign n1459 = x18 & x43;
  assign n1460 = n1458 & n1459;
  assign n1461 = n1458 | n1459;
  assign n1462 = ~n1460 & n1461;
  assign n1463 = n2862 & n1462;
  assign n1464 = n2862 | n1462;
  assign n1465 = ~n1463 & n1464;
  assign n1466 = x17 & x44;
  assign n1467 = n1465 & n1466;
  assign n1468 = n1465 | n1466;
  assign n1469 = ~n1467 & n1468;
  assign n1470 = n1374 & n1469;
  assign n1471 = n1374 | n1469;
  assign n1472 = ~n1470 & n1471;
  assign n1473 = x16 & x45;
  assign n1474 = n1472 & n1473;
  assign n1475 = n1472 | n1473;
  assign n1476 = ~n1474 & n1475;
  assign n2894 = n1374 | n1467;
  assign n2895 = (n1467 & n1469) | (n1467 & n2894) | (n1469 & n2894);
  assign n2896 = n1460 | n2862;
  assign n2897 = (n1460 & n1462) | (n1460 & n2896) | (n1462 & n2896);
  assign n2898 = n1453 | n2864;
  assign n2899 = (n1453 & n1455) | (n1453 & n2898) | (n1455 & n2898);
  assign n2900 = n1446 | n2866;
  assign n2901 = (n1446 & n1448) | (n1446 & n2900) | (n1448 & n2900);
  assign n2902 = n1439 | n1441;
  assign n2903 = (n3533 & n1439) | (n3533 & n2902) | (n1439 & n2902);
  assign n1489 = x30 & x32;
  assign n1490 = x29 & x33;
  assign n1491 = n1489 & n1490;
  assign n1492 = n1489 | n1490;
  assign n1493 = ~n1491 & n1492;
  assign n2910 = n1390 | n1392;
  assign n2912 = n1493 & n2910;
  assign n2913 = n1390 & n1493;
  assign n3544 = (n1297 & n3515) | (n1297 & n3543) | (n3515 & n3543);
  assign n3558 = (n2912 & n2913) | (n2912 & n3544) | (n2913 & n3544);
  assign n3559 = (n2912 & n2913) | (n2912 & n3545) | (n2913 & n3545);
  assign n3560 = (n3482 & n3558) | (n3482 & n3559) | (n3558 & n3559);
  assign n2915 = n1493 | n2910;
  assign n2916 = n1390 | n1493;
  assign n3561 = (n2915 & n2916) | (n2915 & n3544) | (n2916 & n3544);
  assign n3562 = (n2915 & n2916) | (n2915 & n3545) | (n2916 & n3545);
  assign n3563 = (n3482 & n3561) | (n3482 & n3562) | (n3561 & n3562);
  assign n1496 = ~n3560 & n3563;
  assign n1497 = x28 & x34;
  assign n1498 = n1496 & n1497;
  assign n1499 = n1496 | n1497;
  assign n1500 = ~n1498 & n1499;
  assign n2908 = n1397 | n1399;
  assign n2918 = n1500 & n2908;
  assign n2919 = n1397 & n1500;
  assign n3564 = (n2918 & n2919) | (n2918 & n3540) | (n2919 & n3540);
  assign n3565 = (n2918 & n2919) | (n2918 & n3542) | (n2919 & n3542);
  assign n3566 = (n3499 & n3564) | (n3499 & n3565) | (n3564 & n3565);
  assign n2921 = n1500 | n2908;
  assign n2922 = n1397 | n1500;
  assign n3567 = (n2921 & n2922) | (n2921 & n3540) | (n2922 & n3540);
  assign n3568 = (n2921 & n2922) | (n2921 & n3542) | (n2922 & n3542);
  assign n3569 = (n3499 & n3567) | (n3499 & n3568) | (n3567 & n3568);
  assign n1503 = ~n3566 & n3569;
  assign n1504 = x27 & x35;
  assign n1505 = n1503 & n1504;
  assign n1506 = n1503 | n1504;
  assign n1507 = ~n1505 & n1506;
  assign n2906 = n1404 | n1406;
  assign n2924 = n1507 & n2906;
  assign n2925 = n1404 & n1507;
  assign n2926 = (n3538 & n2924) | (n3538 & n2925) | (n2924 & n2925);
  assign n2927 = n1507 | n2906;
  assign n2928 = n1404 | n1507;
  assign n2929 = (n3538 & n2927) | (n3538 & n2928) | (n2927 & n2928);
  assign n1510 = ~n2926 & n2929;
  assign n1511 = x26 & x36;
  assign n1512 = n1510 & n1511;
  assign n1513 = n1510 | n1511;
  assign n1514 = ~n1512 & n1513;
  assign n2930 = n1411 & n1514;
  assign n3570 = (n1514 & n2880) | (n1514 & n2930) | (n2880 & n2930);
  assign n3571 = (n1413 & n1514) | (n1413 & n2930) | (n1514 & n2930);
  assign n3572 = (n2852 & n3570) | (n2852 & n3571) | (n3570 & n3571);
  assign n2932 = n1411 | n1514;
  assign n3573 = n2880 | n2932;
  assign n3574 = n1413 | n2932;
  assign n3575 = (n2852 & n3573) | (n2852 & n3574) | (n3573 & n3574);
  assign n1517 = ~n3572 & n3575;
  assign n1518 = x25 & x37;
  assign n1519 = n1517 & n1518;
  assign n1520 = n1517 | n1518;
  assign n1521 = ~n1519 & n1520;
  assign n2934 = n1418 & n1521;
  assign n2935 = (n1521 & n2885) | (n1521 & n2934) | (n2885 & n2934);
  assign n2936 = n1418 | n1521;
  assign n2937 = n2885 | n2936;
  assign n1524 = ~n2935 & n2937;
  assign n1525 = x24 & x38;
  assign n1526 = n1524 & n1525;
  assign n1527 = n1524 | n1525;
  assign n1528 = ~n1526 & n1527;
  assign n2938 = n1425 & n1528;
  assign n2939 = (n1528 & n2890) | (n1528 & n2938) | (n2890 & n2938);
  assign n2940 = n1425 | n1528;
  assign n2941 = n2890 | n2940;
  assign n1531 = ~n2939 & n2941;
  assign n1532 = x23 & x39;
  assign n1533 = n1531 & n1532;
  assign n1534 = n1531 | n1532;
  assign n1535 = ~n1533 & n1534;
  assign n2904 = n1432 | n1434;
  assign n2942 = n1535 & n2904;
  assign n2943 = n1432 & n1535;
  assign n2944 = (n2868 & n2942) | (n2868 & n2943) | (n2942 & n2943);
  assign n2945 = n1535 | n2904;
  assign n2946 = n1432 | n1535;
  assign n2947 = (n2868 & n2945) | (n2868 & n2946) | (n2945 & n2946);
  assign n1538 = ~n2944 & n2947;
  assign n1539 = x22 & x40;
  assign n1540 = n1538 & n1539;
  assign n1541 = n1538 | n1539;
  assign n1542 = ~n1540 & n1541;
  assign n1543 = n2903 & n1542;
  assign n1544 = n2903 | n1542;
  assign n1545 = ~n1543 & n1544;
  assign n1546 = x21 & x41;
  assign n1547 = n1545 & n1546;
  assign n1548 = n1545 | n1546;
  assign n1549 = ~n1547 & n1548;
  assign n1550 = n2901 & n1549;
  assign n1551 = n2901 | n1549;
  assign n1552 = ~n1550 & n1551;
  assign n1553 = x20 & x42;
  assign n1554 = n1552 & n1553;
  assign n1555 = n1552 | n1553;
  assign n1556 = ~n1554 & n1555;
  assign n1557 = n2899 & n1556;
  assign n1558 = n2899 | n1556;
  assign n1559 = ~n1557 & n1558;
  assign n1560 = x19 & x43;
  assign n1561 = n1559 & n1560;
  assign n1562 = n1559 | n1560;
  assign n1563 = ~n1561 & n1562;
  assign n1564 = n2897 & n1563;
  assign n1565 = n2897 | n1563;
  assign n1566 = ~n1564 & n1565;
  assign n1567 = x18 & x44;
  assign n1568 = n1566 & n1567;
  assign n1569 = n1566 | n1567;
  assign n1570 = ~n1568 & n1569;
  assign n1571 = n2895 & n1570;
  assign n1572 = n2895 | n1570;
  assign n1573 = ~n1571 & n1572;
  assign n1574 = x17 & x45;
  assign n1575 = n1573 & n1574;
  assign n1576 = n1573 | n1574;
  assign n1577 = ~n1575 & n1576;
  assign n1578 = n1474 & n1577;
  assign n1579 = n1474 | n1577;
  assign n1580 = ~n1578 & n1579;
  assign n1581 = x16 & x46;
  assign n1582 = n1580 & n1581;
  assign n1583 = n1580 | n1581;
  assign n1584 = ~n1582 & n1583;
  assign n3913 = n1473 | n1574;
  assign n3914 = (n1472 & n1574) | (n1472 & n3913) | (n1574 & n3913);
  assign n3577 = (n1474 & n1573) | (n1474 & n3914) | (n1573 & n3914);
  assign n2949 = (n1575 & n1577) | (n1575 & n3577) | (n1577 & n3577);
  assign n3578 = n1568 | n2895;
  assign n3579 = (n1568 & n1570) | (n1568 & n3578) | (n1570 & n3578);
  assign n1587 = n1561 | n1564;
  assign n1588 = n1554 | n1557;
  assign n2953 = n1512 | n1514;
  assign n3580 = n1411 | n1512;
  assign n3581 = (n1512 & n1514) | (n1512 & n3580) | (n1514 & n3580);
  assign n3582 = (n2880 & n2953) | (n2880 & n3581) | (n2953 & n3581);
  assign n3583 = (n1413 & n2953) | (n1413 & n3581) | (n2953 & n3581);
  assign n3584 = (n2852 & n3582) | (n2852 & n3583) | (n3582 & n3583);
  assign n3585 = n1498 | n1500;
  assign n3586 = (n1498 & n2908) | (n1498 & n3585) | (n2908 & n3585);
  assign n3587 = n1397 | n1498;
  assign n3588 = (n1498 & n1500) | (n1498 & n3587) | (n1500 & n3587);
  assign n3589 = (n3540 & n3586) | (n3540 & n3588) | (n3586 & n3588);
  assign n3590 = (n3542 & n3586) | (n3542 & n3588) | (n3586 & n3588);
  assign n3591 = (n3499 & n3589) | (n3499 & n3590) | (n3589 & n3590);
  assign n1598 = x31 & x32;
  assign n1599 = x30 & x33;
  assign n1600 = n1598 & n1599;
  assign n1601 = n1598 | n1599;
  assign n1602 = ~n1600 & n1601;
  assign n3592 = n1491 | n1493;
  assign n3593 = (n1491 & n2910) | (n1491 & n3592) | (n2910 & n3592);
  assign n2961 = n1602 & n3593;
  assign n3594 = n1390 | n1491;
  assign n3595 = (n1491 & n1493) | (n1491 & n3594) | (n1493 & n3594);
  assign n2962 = n1602 & n3595;
  assign n3596 = (n2961 & n2962) | (n2961 & n3544) | (n2962 & n3544);
  assign n3597 = (n2961 & n2962) | (n2961 & n3545) | (n2962 & n3545);
  assign n3598 = (n3482 & n3596) | (n3482 & n3597) | (n3596 & n3597);
  assign n2964 = n1602 | n3593;
  assign n2965 = n1602 | n3595;
  assign n3599 = (n2964 & n2965) | (n2964 & n3544) | (n2965 & n3544);
  assign n3600 = (n2964 & n2965) | (n2964 & n3545) | (n2965 & n3545);
  assign n3601 = (n3482 & n3599) | (n3482 & n3600) | (n3599 & n3600);
  assign n1605 = ~n3598 & n3601;
  assign n1606 = x29 & x34;
  assign n1607 = n1605 & n1606;
  assign n1608 = n1605 | n1606;
  assign n1609 = ~n1607 & n1608;
  assign n1610 = n3591 & n1609;
  assign n1611 = n3591 | n1609;
  assign n1612 = ~n1610 & n1611;
  assign n1613 = x28 & x35;
  assign n1614 = n1612 & n1613;
  assign n1615 = n1612 | n1613;
  assign n1616 = ~n1614 & n1615;
  assign n2967 = n1505 & n1616;
  assign n3602 = (n1616 & n2924) | (n1616 & n2967) | (n2924 & n2967);
  assign n3603 = (n1616 & n2925) | (n1616 & n2967) | (n2925 & n2967);
  assign n3604 = (n3538 & n3602) | (n3538 & n3603) | (n3602 & n3603);
  assign n2969 = n1505 | n1616;
  assign n3605 = n2924 | n2969;
  assign n3606 = n2925 | n2969;
  assign n3607 = (n3538 & n3605) | (n3538 & n3606) | (n3605 & n3606);
  assign n1619 = ~n3604 & n3607;
  assign n1620 = x27 & x36;
  assign n1621 = n1619 & n1620;
  assign n1622 = n1619 | n1620;
  assign n1623 = ~n1621 & n1622;
  assign n1624 = n3584 & n1623;
  assign n1625 = n3584 | n1623;
  assign n1626 = ~n1624 & n1625;
  assign n1627 = x26 & x37;
  assign n1628 = n1626 & n1627;
  assign n1629 = n1626 | n1627;
  assign n1630 = ~n1628 & n1629;
  assign n2971 = n1519 & n1630;
  assign n2972 = (n1630 & n2935) | (n1630 & n2971) | (n2935 & n2971);
  assign n2973 = n1519 | n1630;
  assign n2974 = n2935 | n2973;
  assign n1633 = ~n2972 & n2974;
  assign n1634 = x25 & x38;
  assign n1635 = n1633 & n1634;
  assign n1636 = n1633 | n1634;
  assign n1637 = ~n1635 & n1636;
  assign n2975 = n1526 & n1637;
  assign n2976 = (n1637 & n2939) | (n1637 & n2975) | (n2939 & n2975);
  assign n2977 = n1526 | n1637;
  assign n2978 = n2939 | n2977;
  assign n1640 = ~n2976 & n2978;
  assign n1641 = x24 & x39;
  assign n1642 = n1640 & n1641;
  assign n1643 = n1640 | n1641;
  assign n1644 = ~n1642 & n1643;
  assign n2979 = n1533 & n1644;
  assign n2980 = (n1644 & n2944) | (n1644 & n2979) | (n2944 & n2979);
  assign n2981 = n1533 | n1644;
  assign n2982 = n2944 | n2981;
  assign n1647 = ~n2980 & n2982;
  assign n1648 = x23 & x40;
  assign n1649 = n1647 & n1648;
  assign n1650 = n1647 | n1648;
  assign n1651 = ~n1649 & n1650;
  assign n2950 = n1540 | n1542;
  assign n2983 = n1651 & n2950;
  assign n2984 = n1540 & n1651;
  assign n2985 = (n2903 & n2983) | (n2903 & n2984) | (n2983 & n2984);
  assign n2986 = n1651 | n2950;
  assign n2987 = n1540 | n1651;
  assign n2988 = (n2903 & n2986) | (n2903 & n2987) | (n2986 & n2987);
  assign n1654 = ~n2985 & n2988;
  assign n1655 = x22 & x41;
  assign n1656 = n1654 & n1655;
  assign n1657 = n1654 | n1655;
  assign n1658 = ~n1656 & n1657;
  assign n2989 = n1547 & n1658;
  assign n2990 = (n1550 & n1658) | (n1550 & n2989) | (n1658 & n2989);
  assign n2991 = n1547 | n1658;
  assign n2992 = n1550 | n2991;
  assign n1661 = ~n2990 & n2992;
  assign n1662 = x21 & x42;
  assign n1663 = n1661 & n1662;
  assign n1664 = n1661 | n1662;
  assign n1665 = ~n1663 & n1664;
  assign n1666 = n1588 & n1665;
  assign n1667 = n1588 | n1665;
  assign n1668 = ~n1666 & n1667;
  assign n1669 = x20 & x43;
  assign n1670 = n1668 & n1669;
  assign n1671 = n1668 | n1669;
  assign n1672 = ~n1670 & n1671;
  assign n1673 = n1587 & n1672;
  assign n1674 = n1587 | n1672;
  assign n1675 = ~n1673 & n1674;
  assign n1676 = x19 & x44;
  assign n1677 = n1675 & n1676;
  assign n1678 = n1675 | n1676;
  assign n1679 = ~n1677 & n1678;
  assign n1680 = n3579 & n1679;
  assign n1681 = n3579 | n1679;
  assign n1682 = ~n1680 & n1681;
  assign n1683 = x18 & x45;
  assign n1684 = n1682 & n1683;
  assign n1685 = n1682 | n1683;
  assign n1686 = ~n1684 & n1685;
  assign n1687 = n2949 & n1686;
  assign n1688 = n2949 | n1686;
  assign n1689 = ~n1687 & n1688;
  assign n1690 = x17 & x46;
  assign n1691 = n1689 & n1690;
  assign n1692 = n1689 | n1690;
  assign n1693 = ~n1691 & n1692;
  assign n1694 = n1582 & n1693;
  assign n1695 = n1582 | n1693;
  assign n1696 = ~n1694 & n1695;
  assign n1697 = x16 & x47;
  assign n1698 = n1696 & n1697;
  assign n1699 = n1696 | n1697;
  assign n1700 = ~n1698 & n1699;
  assign n3915 = n1581 | n1690;
  assign n3916 = (n1580 & n1690) | (n1580 & n3915) | (n1690 & n3915);
  assign n3609 = (n1582 & n1689) | (n1582 & n3916) | (n1689 & n3916);
  assign n2994 = (n1691 & n1693) | (n1691 & n3609) | (n1693 & n3609);
  assign n2995 = n1684 | n2949;
  assign n2996 = (n1684 & n1686) | (n1684 & n2995) | (n1686 & n2995);
  assign n3610 = n1677 | n3579;
  assign n3611 = (n1677 & n1679) | (n1677 & n3610) | (n1679 & n3610);
  assign n1704 = n1670 | n1673;
  assign n2997 = n1663 | n1665;
  assign n2998 = (n1588 & n1663) | (n1588 & n2997) | (n1663 & n2997);
  assign n3002 = n1614 | n1616;
  assign n3612 = n1505 | n1614;
  assign n3613 = (n1614 & n1616) | (n1614 & n3612) | (n1616 & n3612);
  assign n3614 = (n2924 & n3002) | (n2924 & n3613) | (n3002 & n3613);
  assign n3615 = (n2925 & n3002) | (n2925 & n3613) | (n3002 & n3613);
  assign n3616 = (n3538 & n3614) | (n3538 & n3615) | (n3614 & n3615);
  assign n1715 = x31 & x33;
  assign n3617 = n1600 | n1602;
  assign n3622 = (n1600 & n3595) | (n1600 & n3617) | (n3595 & n3617);
  assign n3010 = n1715 & n3622;
  assign n3620 = n1600 & n1715;
  assign n3917 = (n1602 & n1715) | (n1602 & n3620) | (n1715 & n3620);
  assign n3621 = (n3593 & n3917) | (n3593 & n3620) | (n3917 & n3620);
  assign n3623 = (n3010 & n3544) | (n3010 & n3621) | (n3544 & n3621);
  assign n3624 = (n3010 & n3545) | (n3010 & n3621) | (n3545 & n3621);
  assign n3625 = (n3482 & n3623) | (n3482 & n3624) | (n3623 & n3624);
  assign n3013 = n1715 | n3622;
  assign n3627 = n1600 | n1715;
  assign n3918 = n1602 | n3627;
  assign n3628 = (n3593 & n3918) | (n3593 & n3627) | (n3918 & n3627);
  assign n3629 = (n3013 & n3544) | (n3013 & n3628) | (n3544 & n3628);
  assign n3630 = (n3013 & n3545) | (n3013 & n3628) | (n3545 & n3628);
  assign n3631 = (n3482 & n3629) | (n3482 & n3630) | (n3629 & n3630);
  assign n1718 = ~n3625 & n3631;
  assign n1719 = x30 & x34;
  assign n1720 = n1718 & n1719;
  assign n1721 = n1718 | n1719;
  assign n1722 = ~n1720 & n1721;
  assign n3004 = n1607 | n1609;
  assign n3015 = n1722 & n3004;
  assign n3016 = n1607 & n1722;
  assign n3017 = (n3591 & n3015) | (n3591 & n3016) | (n3015 & n3016);
  assign n3018 = n1722 | n3004;
  assign n3019 = n1607 | n1722;
  assign n3020 = (n3591 & n3018) | (n3591 & n3019) | (n3018 & n3019);
  assign n1725 = ~n3017 & n3020;
  assign n1726 = x29 & x35;
  assign n1727 = n1725 & n1726;
  assign n1728 = n1725 | n1726;
  assign n1729 = ~n1727 & n1728;
  assign n1730 = n3616 & n1729;
  assign n1731 = n3616 | n1729;
  assign n1732 = ~n1730 & n1731;
  assign n1733 = x28 & x36;
  assign n1734 = n1732 & n1733;
  assign n1735 = n1732 | n1733;
  assign n1736 = ~n1734 & n1735;
  assign n2999 = n1621 | n1623;
  assign n3021 = n1736 & n2999;
  assign n3022 = n1621 & n1736;
  assign n3023 = (n3584 & n3021) | (n3584 & n3022) | (n3021 & n3022);
  assign n3024 = n1736 | n2999;
  assign n3025 = n1621 | n1736;
  assign n3026 = (n3584 & n3024) | (n3584 & n3025) | (n3024 & n3025);
  assign n1739 = ~n3023 & n3026;
  assign n1740 = x27 & x37;
  assign n1741 = n1739 & n1740;
  assign n1742 = n1739 | n1740;
  assign n1743 = ~n1741 & n1742;
  assign n3027 = n1628 & n1743;
  assign n3632 = (n1743 & n2971) | (n1743 & n3027) | (n2971 & n3027);
  assign n3633 = (n1630 & n1743) | (n1630 & n3027) | (n1743 & n3027);
  assign n3634 = (n2935 & n3632) | (n2935 & n3633) | (n3632 & n3633);
  assign n3029 = n1628 | n1743;
  assign n3635 = n2971 | n3029;
  assign n3636 = n1630 | n3029;
  assign n3637 = (n2935 & n3635) | (n2935 & n3636) | (n3635 & n3636);
  assign n1746 = ~n3634 & n3637;
  assign n1747 = x26 & x38;
  assign n1748 = n1746 & n1747;
  assign n1749 = n1746 | n1747;
  assign n1750 = ~n1748 & n1749;
  assign n3031 = n1635 & n1750;
  assign n3032 = (n1750 & n2976) | (n1750 & n3031) | (n2976 & n3031);
  assign n3033 = n1635 | n1750;
  assign n3034 = n2976 | n3033;
  assign n1753 = ~n3032 & n3034;
  assign n1754 = x25 & x39;
  assign n1755 = n1753 & n1754;
  assign n1756 = n1753 | n1754;
  assign n1757 = ~n1755 & n1756;
  assign n3035 = n1642 & n1757;
  assign n3036 = (n1757 & n2980) | (n1757 & n3035) | (n2980 & n3035);
  assign n3037 = n1642 | n1757;
  assign n3038 = n2980 | n3037;
  assign n1760 = ~n3036 & n3038;
  assign n1761 = x24 & x40;
  assign n1762 = n1760 & n1761;
  assign n1763 = n1760 | n1761;
  assign n1764 = ~n1762 & n1763;
  assign n3039 = n1649 & n1764;
  assign n3040 = (n1764 & n2985) | (n1764 & n3039) | (n2985 & n3039);
  assign n3041 = n1649 | n1764;
  assign n3042 = n2985 | n3041;
  assign n1767 = ~n3040 & n3042;
  assign n1768 = x23 & x41;
  assign n1769 = n1767 & n1768;
  assign n1770 = n1767 | n1768;
  assign n1771 = ~n1769 & n1770;
  assign n3043 = n1656 & n1771;
  assign n3044 = (n1771 & n2990) | (n1771 & n3043) | (n2990 & n3043);
  assign n3045 = n1656 | n1771;
  assign n3046 = n2990 | n3045;
  assign n1774 = ~n3044 & n3046;
  assign n1775 = x22 & x42;
  assign n1776 = n1774 & n1775;
  assign n1777 = n1774 | n1775;
  assign n1778 = ~n1776 & n1777;
  assign n1779 = n2998 & n1778;
  assign n1780 = n2998 | n1778;
  assign n1781 = ~n1779 & n1780;
  assign n1782 = x21 & x43;
  assign n1783 = n1781 & n1782;
  assign n1784 = n1781 | n1782;
  assign n1785 = ~n1783 & n1784;
  assign n1786 = n1704 & n1785;
  assign n1787 = n1704 | n1785;
  assign n1788 = ~n1786 & n1787;
  assign n1789 = x20 & x44;
  assign n1790 = n1788 & n1789;
  assign n1791 = n1788 | n1789;
  assign n1792 = ~n1790 & n1791;
  assign n1793 = n3611 & n1792;
  assign n1794 = n3611 | n1792;
  assign n1795 = ~n1793 & n1794;
  assign n1796 = x19 & x45;
  assign n1797 = n1795 & n1796;
  assign n1798 = n1795 | n1796;
  assign n1799 = ~n1797 & n1798;
  assign n1800 = n2996 & n1799;
  assign n1801 = n2996 | n1799;
  assign n1802 = ~n1800 & n1801;
  assign n1803 = x18 & x46;
  assign n1804 = n1802 & n1803;
  assign n1805 = n1802 | n1803;
  assign n1806 = ~n1804 & n1805;
  assign n1807 = n2994 & n1806;
  assign n1808 = n2994 | n1806;
  assign n1809 = ~n1807 & n1808;
  assign n1810 = x17 & x47;
  assign n1811 = n1809 & n1810;
  assign n1812 = n1809 | n1810;
  assign n1813 = ~n1811 & n1812;
  assign n1814 = n1698 & n1813;
  assign n1815 = n1698 | n1813;
  assign n1816 = ~n1814 & n1815;
  assign n3919 = n1697 | n1810;
  assign n3920 = (n1696 & n1810) | (n1696 & n3919) | (n1810 & n3919);
  assign n3639 = (n1698 & n1809) | (n1698 & n3920) | (n1809 & n3920);
  assign n3048 = (n1811 & n1813) | (n1811 & n3639) | (n1813 & n3639);
  assign n3049 = n1804 | n2994;
  assign n3050 = (n1804 & n1806) | (n1804 & n3049) | (n1806 & n3049);
  assign n3051 = n1797 | n2996;
  assign n3052 = (n1797 & n1799) | (n1797 & n3051) | (n1799 & n3051);
  assign n3640 = n1790 | n3611;
  assign n3641 = (n1790 & n1792) | (n1790 & n3640) | (n1792 & n3640);
  assign n3053 = n1783 | n1785;
  assign n3054 = (n1704 & n1783) | (n1704 & n3053) | (n1783 & n3053);
  assign n3055 = n1776 | n1778;
  assign n3056 = (n1776 & n2998) | (n1776 & n3055) | (n2998 & n3055);
  assign n3058 = n1741 | n1743;
  assign n3642 = n1628 | n1741;
  assign n3643 = (n1741 & n1743) | (n1741 & n3642) | (n1743 & n3642);
  assign n3644 = (n2971 & n3058) | (n2971 & n3643) | (n3058 & n3643);
  assign n3645 = (n1630 & n3058) | (n1630 & n3643) | (n3058 & n3643);
  assign n3646 = (n2935 & n3644) | (n2935 & n3645) | (n3644 & n3645);
  assign n1831 = x31 & x34;
  assign n1832 = n3625 & n1831;
  assign n1833 = n3625 | n1831;
  assign n1834 = ~n1832 & n1833;
  assign n3647 = n1720 | n1722;
  assign n3648 = (n1720 & n3004) | (n1720 & n3647) | (n3004 & n3647);
  assign n3065 = n1834 & n3648;
  assign n3649 = n1607 | n1720;
  assign n3650 = (n1720 & n1722) | (n1720 & n3649) | (n1722 & n3649);
  assign n3066 = n1834 & n3650;
  assign n3067 = (n3591 & n3065) | (n3591 & n3066) | (n3065 & n3066);
  assign n3068 = n1834 | n3648;
  assign n3069 = n1834 | n3650;
  assign n3070 = (n3591 & n3068) | (n3591 & n3069) | (n3068 & n3069);
  assign n1837 = ~n3067 & n3070;
  assign n1838 = x30 & x35;
  assign n1839 = n1837 & n1838;
  assign n1840 = n1837 | n1838;
  assign n1841 = ~n1839 & n1840;
  assign n3060 = n1727 | n1729;
  assign n3071 = n1841 & n3060;
  assign n3072 = n1727 & n1841;
  assign n3073 = (n3616 & n3071) | (n3616 & n3072) | (n3071 & n3072);
  assign n3074 = n1841 | n3060;
  assign n3075 = n1727 | n1841;
  assign n3076 = (n3616 & n3074) | (n3616 & n3075) | (n3074 & n3075);
  assign n1844 = ~n3073 & n3076;
  assign n1845 = x29 & x36;
  assign n1846 = n1844 & n1845;
  assign n1847 = n1844 | n1845;
  assign n1848 = ~n1846 & n1847;
  assign n3077 = n1734 & n1848;
  assign n3651 = (n1848 & n3022) | (n1848 & n3077) | (n3022 & n3077);
  assign n3652 = (n1848 & n3021) | (n1848 & n3077) | (n3021 & n3077);
  assign n3653 = (n3584 & n3651) | (n3584 & n3652) | (n3651 & n3652);
  assign n3079 = n1734 | n1848;
  assign n3654 = n3022 | n3079;
  assign n3655 = n3021 | n3079;
  assign n3656 = (n3584 & n3654) | (n3584 & n3655) | (n3654 & n3655);
  assign n1851 = ~n3653 & n3656;
  assign n1852 = x28 & x37;
  assign n1853 = n1851 & n1852;
  assign n1854 = n1851 | n1852;
  assign n1855 = ~n1853 & n1854;
  assign n1856 = n3646 & n1855;
  assign n1857 = n3646 | n1855;
  assign n1858 = ~n1856 & n1857;
  assign n1859 = x27 & x38;
  assign n1860 = n1858 & n1859;
  assign n1861 = n1858 | n1859;
  assign n1862 = ~n1860 & n1861;
  assign n3081 = n1748 & n1862;
  assign n3082 = (n1862 & n3032) | (n1862 & n3081) | (n3032 & n3081);
  assign n3083 = n1748 | n1862;
  assign n3084 = n3032 | n3083;
  assign n1865 = ~n3082 & n3084;
  assign n1866 = x26 & x39;
  assign n1867 = n1865 & n1866;
  assign n1868 = n1865 | n1866;
  assign n1869 = ~n1867 & n1868;
  assign n3085 = n1755 & n1869;
  assign n3086 = (n1869 & n3036) | (n1869 & n3085) | (n3036 & n3085);
  assign n3087 = n1755 | n1869;
  assign n3088 = n3036 | n3087;
  assign n1872 = ~n3086 & n3088;
  assign n1873 = x25 & x40;
  assign n1874 = n1872 & n1873;
  assign n1875 = n1872 | n1873;
  assign n1876 = ~n1874 & n1875;
  assign n3089 = n1762 & n1876;
  assign n3090 = (n1876 & n3040) | (n1876 & n3089) | (n3040 & n3089);
  assign n3091 = n1762 | n1876;
  assign n3092 = n3040 | n3091;
  assign n1879 = ~n3090 & n3092;
  assign n1880 = x24 & x41;
  assign n1881 = n1879 & n1880;
  assign n1882 = n1879 | n1880;
  assign n1883 = ~n1881 & n1882;
  assign n3093 = n1769 & n1883;
  assign n3094 = (n1883 & n3044) | (n1883 & n3093) | (n3044 & n3093);
  assign n3095 = n1769 | n1883;
  assign n3096 = n3044 | n3095;
  assign n1886 = ~n3094 & n3096;
  assign n1887 = x23 & x42;
  assign n1888 = n1886 & n1887;
  assign n1889 = n1886 | n1887;
  assign n1890 = ~n1888 & n1889;
  assign n1891 = n3056 & n1890;
  assign n1892 = n3056 | n1890;
  assign n1893 = ~n1891 & n1892;
  assign n1894 = x22 & x43;
  assign n1895 = n1893 & n1894;
  assign n1896 = n1893 | n1894;
  assign n1897 = ~n1895 & n1896;
  assign n1898 = n3054 & n1897;
  assign n1899 = n3054 | n1897;
  assign n1900 = ~n1898 & n1899;
  assign n1901 = x21 & x44;
  assign n1902 = n1900 & n1901;
  assign n1903 = n1900 | n1901;
  assign n1904 = ~n1902 & n1903;
  assign n1905 = n3641 & n1904;
  assign n1906 = n3641 | n1904;
  assign n1907 = ~n1905 & n1906;
  assign n1908 = x20 & x45;
  assign n1909 = n1907 & n1908;
  assign n1910 = n1907 | n1908;
  assign n1911 = ~n1909 & n1910;
  assign n1912 = n3052 & n1911;
  assign n1913 = n3052 | n1911;
  assign n1914 = ~n1912 & n1913;
  assign n1915 = x19 & x46;
  assign n1916 = n1914 & n1915;
  assign n1917 = n1914 | n1915;
  assign n1918 = ~n1916 & n1917;
  assign n1919 = n3050 & n1918;
  assign n1920 = n3050 | n1918;
  assign n1921 = ~n1919 & n1920;
  assign n1922 = x18 & x47;
  assign n1923 = n1921 & n1922;
  assign n1924 = n1921 | n1922;
  assign n1925 = ~n1923 & n1924;
  assign n1926 = n3048 & n1925;
  assign n1927 = n3048 | n1925;
  assign n1928 = ~n1926 & n1927;
  assign n3097 = n1923 | n3048;
  assign n3098 = (n1923 & n1925) | (n1923 & n3097) | (n1925 & n3097);
  assign n3099 = n1916 | n3050;
  assign n3100 = (n1916 & n1918) | (n1916 & n3099) | (n1918 & n3099);
  assign n3101 = n1909 | n3052;
  assign n3102 = (n1909 & n1911) | (n1909 & n3101) | (n1911 & n3101);
  assign n3103 = n1902 | n1904;
  assign n3104 = (n3641 & n1902) | (n3641 & n3103) | (n1902 & n3103);
  assign n3105 = n1895 | n1897;
  assign n3106 = (n1895 & n3054) | (n1895 & n3105) | (n3054 & n3105);
  assign n3107 = n1888 | n1890;
  assign n3108 = (n1888 & n3056) | (n1888 & n3107) | (n3056 & n3107);
  assign n3112 = n1846 | n1848;
  assign n3657 = n1734 | n1846;
  assign n3658 = (n1846 & n1848) | (n1846 & n3657) | (n1848 & n3657);
  assign n3659 = (n3022 & n3112) | (n3022 & n3658) | (n3112 & n3658);
  assign n3660 = (n3021 & n3112) | (n3021 & n3658) | (n3112 & n3658);
  assign n3661 = (n3584 & n3659) | (n3584 & n3660) | (n3659 & n3660);
  assign n1943 = x31 & x35;
  assign n3666 = n1831 & n1943;
  assign n3667 = n3625 & n3666;
  assign n3921 = (n1834 & n1943) | (n1834 & n3667) | (n1943 & n3667);
  assign n11946 = n1943 & n3666;
  assign n11947 = n3625 & n11946;
  assign n3923 = (n3648 & n3921) | (n3648 & n11947) | (n3921 & n11947);
  assign n3924 = (n3650 & n3921) | (n3650 & n11947) | (n3921 & n11947);
  assign n3670 = (n3591 & n3923) | (n3591 & n3924) | (n3923 & n3924);
  assign n3671 = n1831 | n1943;
  assign n3672 = (n1943 & n3625) | (n1943 & n3671) | (n3625 & n3671);
  assign n3925 = n1834 | n3672;
  assign n3926 = (n3648 & n3672) | (n3648 & n3925) | (n3672 & n3925);
  assign n3927 = (n3650 & n3672) | (n3650 & n3925) | (n3672 & n3925);
  assign n3675 = (n3591 & n3926) | (n3591 & n3927) | (n3926 & n3927);
  assign n1946 = ~n3670 & n3675;
  assign n3662 = n1839 | n1841;
  assign n3663 = (n1839 & n3060) | (n1839 & n3662) | (n3060 & n3662);
  assign n3676 = n1946 & n3663;
  assign n3664 = n1727 | n1839;
  assign n3665 = (n1839 & n1841) | (n1839 & n3664) | (n1841 & n3664);
  assign n3677 = n1946 & n3665;
  assign n3678 = (n3616 & n3676) | (n3616 & n3677) | (n3676 & n3677);
  assign n3679 = n1946 | n3663;
  assign n3680 = n1946 | n3665;
  assign n3681 = (n3616 & n3679) | (n3616 & n3680) | (n3679 & n3680);
  assign n1949 = ~n3678 & n3681;
  assign n1950 = x30 & x36;
  assign n1951 = n1949 & n1950;
  assign n1952 = n1949 | n1950;
  assign n1953 = ~n1951 & n1952;
  assign n1954 = n3661 & n1953;
  assign n1955 = n3661 | n1953;
  assign n1956 = ~n1954 & n1955;
  assign n1957 = x29 & x37;
  assign n1958 = n1956 & n1957;
  assign n1959 = n1956 | n1957;
  assign n1960 = ~n1958 & n1959;
  assign n3109 = n1853 | n1855;
  assign n3121 = n1960 & n3109;
  assign n3122 = n1853 & n1960;
  assign n3123 = (n3646 & n3121) | (n3646 & n3122) | (n3121 & n3122);
  assign n3124 = n1960 | n3109;
  assign n3125 = n1853 | n1960;
  assign n3126 = (n3646 & n3124) | (n3646 & n3125) | (n3124 & n3125);
  assign n1963 = ~n3123 & n3126;
  assign n1964 = x28 & x38;
  assign n1965 = n1963 & n1964;
  assign n1966 = n1963 | n1964;
  assign n1967 = ~n1965 & n1966;
  assign n3127 = n1860 & n1967;
  assign n3682 = (n1967 & n3081) | (n1967 & n3127) | (n3081 & n3127);
  assign n3683 = (n1862 & n1967) | (n1862 & n3127) | (n1967 & n3127);
  assign n3684 = (n3032 & n3682) | (n3032 & n3683) | (n3682 & n3683);
  assign n3129 = n1860 | n1967;
  assign n3685 = n3081 | n3129;
  assign n3686 = n1862 | n3129;
  assign n3687 = (n3032 & n3685) | (n3032 & n3686) | (n3685 & n3686);
  assign n1970 = ~n3684 & n3687;
  assign n1971 = x27 & x39;
  assign n1972 = n1970 & n1971;
  assign n1973 = n1970 | n1971;
  assign n1974 = ~n1972 & n1973;
  assign n3131 = n1867 & n1974;
  assign n3132 = (n1974 & n3086) | (n1974 & n3131) | (n3086 & n3131);
  assign n3133 = n1867 | n1974;
  assign n3134 = n3086 | n3133;
  assign n1977 = ~n3132 & n3134;
  assign n1978 = x26 & x40;
  assign n1979 = n1977 & n1978;
  assign n1980 = n1977 | n1978;
  assign n1981 = ~n1979 & n1980;
  assign n3135 = n1874 & n1981;
  assign n3136 = (n1981 & n3090) | (n1981 & n3135) | (n3090 & n3135);
  assign n3137 = n1874 | n1981;
  assign n3138 = n3090 | n3137;
  assign n1984 = ~n3136 & n3138;
  assign n1985 = x25 & x41;
  assign n1986 = n1984 & n1985;
  assign n1987 = n1984 | n1985;
  assign n1988 = ~n1986 & n1987;
  assign n3139 = n1881 & n1988;
  assign n3140 = (n1988 & n3094) | (n1988 & n3139) | (n3094 & n3139);
  assign n3141 = n1881 | n1988;
  assign n3142 = n3094 | n3141;
  assign n1991 = ~n3140 & n3142;
  assign n1992 = x24 & x42;
  assign n1993 = n1991 & n1992;
  assign n1994 = n1991 | n1992;
  assign n1995 = ~n1993 & n1994;
  assign n1996 = n3108 & n1995;
  assign n1997 = n3108 | n1995;
  assign n1998 = ~n1996 & n1997;
  assign n1999 = x23 & x43;
  assign n2000 = n1998 & n1999;
  assign n2001 = n1998 | n1999;
  assign n2002 = ~n2000 & n2001;
  assign n2003 = n3106 & n2002;
  assign n2004 = n3106 | n2002;
  assign n2005 = ~n2003 & n2004;
  assign n2006 = x22 & x44;
  assign n2007 = n2005 & n2006;
  assign n2008 = n2005 | n2006;
  assign n2009 = ~n2007 & n2008;
  assign n2010 = n3104 & n2009;
  assign n2011 = n3104 | n2009;
  assign n2012 = ~n2010 & n2011;
  assign n2013 = x21 & x45;
  assign n2014 = n2012 & n2013;
  assign n2015 = n2012 | n2013;
  assign n2016 = ~n2014 & n2015;
  assign n2017 = n3102 & n2016;
  assign n2018 = n3102 | n2016;
  assign n2019 = ~n2017 & n2018;
  assign n2020 = x20 & x46;
  assign n2021 = n2019 & n2020;
  assign n2022 = n2019 | n2020;
  assign n2023 = ~n2021 & n2022;
  assign n2024 = n3100 & n2023;
  assign n2025 = n3100 | n2023;
  assign n2026 = ~n2024 & n2025;
  assign n2027 = x19 & x47;
  assign n2028 = n2026 & n2027;
  assign n2029 = n2026 | n2027;
  assign n2030 = ~n2028 & n2029;
  assign n2031 = n3098 & n2030;
  assign n2032 = n3098 | n2030;
  assign n2033 = ~n2031 & n2032;
  assign n2034 = n2028 | n2031;
  assign n2035 = n2021 | n2024;
  assign n2036 = n2014 | n2017;
  assign n3143 = n2007 | n2009;
  assign n3144 = (n2007 & n3104) | (n2007 & n3143) | (n3104 & n3143);
  assign n3145 = n2000 | n2002;
  assign n3146 = (n2000 & n3106) | (n2000 & n3145) | (n3106 & n3145);
  assign n3147 = n1993 | n1995;
  assign n3148 = (n1993 & n3108) | (n1993 & n3147) | (n3108 & n3147);
  assign n3150 = n1965 | n1967;
  assign n3688 = n1860 | n1965;
  assign n3689 = (n1965 & n1967) | (n1965 & n3688) | (n1967 & n3688);
  assign n3690 = (n3081 & n3150) | (n3081 & n3689) | (n3150 & n3689);
  assign n3691 = (n1862 & n3150) | (n1862 & n3689) | (n3150 & n3689);
  assign n3692 = (n3032 & n3690) | (n3032 & n3691) | (n3690 & n3691);
  assign n2047 = x31 & x36;
  assign n17664 = n2047 & n3666;
  assign n17665 = n3625 & n17664;
  assign n15577 = n1943 & n2047;
  assign n15578 = (n1834 & n17665) | (n1834 & n15577) | (n17665 & n15577);
  assign n17666 = n3666 & n15577;
  assign n15580 = n3625 & n17666;
  assign n11950 = (n3648 & n15578) | (n3648 & n15580) | (n15578 & n15580);
  assign n11951 = (n3650 & n15578) | (n3650 & n15580) | (n15578 & n15580);
  assign n3930 = (n3591 & n11950) | (n3591 & n11951) | (n11950 & n11951);
  assign n3694 = (n1946 & n2047) | (n1946 & n3930) | (n2047 & n3930);
  assign n3695 = (n3930 & n3663) | (n3930 & n3694) | (n3663 & n3694);
  assign n3696 = (n3930 & n3665) | (n3930 & n3694) | (n3665 & n3694);
  assign n3697 = (n3616 & n3695) | (n3616 & n3696) | (n3695 & n3696);
  assign n17667 = n2047 | n3666;
  assign n17668 = (n2047 & n3625) | (n2047 & n17667) | (n3625 & n17667);
  assign n15582 = n1943 | n2047;
  assign n15583 = (n1834 & n17668) | (n1834 & n15582) | (n17668 & n15582);
  assign n17669 = (n2047 & n3666) | (n2047 & n15582) | (n3666 & n15582);
  assign n15585 = (n2047 & n3625) | (n2047 & n17669) | (n3625 & n17669);
  assign n11954 = (n3648 & n15583) | (n3648 & n15585) | (n15583 & n15585);
  assign n11955 = (n3650 & n15583) | (n3650 & n15585) | (n15583 & n15585);
  assign n3933 = (n3591 & n11954) | (n3591 & n11955) | (n11954 & n11955);
  assign n3699 = n1946 | n3933;
  assign n3700 = (n3933 & n3663) | (n3933 & n3699) | (n3663 & n3699);
  assign n3701 = (n3933 & n3665) | (n3933 & n3699) | (n3665 & n3699);
  assign n3702 = (n3616 & n3700) | (n3616 & n3701) | (n3700 & n3701);
  assign n2050 = ~n3697 & n3702;
  assign n3163 = n1951 & n2050;
  assign n3703 = (n1953 & n2050) | (n1953 & n3163) | (n2050 & n3163);
  assign n3164 = (n3661 & n3703) | (n3661 & n3163) | (n3703 & n3163);
  assign n3166 = n1951 | n2050;
  assign n3704 = n1953 | n3166;
  assign n3167 = (n3661 & n3704) | (n3661 & n3166) | (n3704 & n3166);
  assign n2053 = ~n3164 & n3167;
  assign n2054 = x30 & x37;
  assign n2055 = n2053 & n2054;
  assign n2056 = n2053 | n2054;
  assign n2057 = ~n2055 & n2056;
  assign n3168 = n1958 & n2057;
  assign n3705 = (n2057 & n3122) | (n2057 & n3168) | (n3122 & n3168);
  assign n3706 = (n2057 & n3121) | (n2057 & n3168) | (n3121 & n3168);
  assign n3707 = (n3646 & n3705) | (n3646 & n3706) | (n3705 & n3706);
  assign n3170 = n1958 | n2057;
  assign n3708 = n3122 | n3170;
  assign n3709 = n3121 | n3170;
  assign n3710 = (n3646 & n3708) | (n3646 & n3709) | (n3708 & n3709);
  assign n2060 = ~n3707 & n3710;
  assign n2061 = x29 & x38;
  assign n2062 = n2060 & n2061;
  assign n2063 = n2060 | n2061;
  assign n2064 = ~n2062 & n2063;
  assign n2065 = n3692 & n2064;
  assign n2066 = n3692 | n2064;
  assign n2067 = ~n2065 & n2066;
  assign n2068 = x28 & x39;
  assign n2069 = n2067 & n2068;
  assign n2070 = n2067 | n2068;
  assign n2071 = ~n2069 & n2070;
  assign n3172 = n1972 & n2071;
  assign n3173 = (n2071 & n3132) | (n2071 & n3172) | (n3132 & n3172);
  assign n3174 = n1972 | n2071;
  assign n3175 = n3132 | n3174;
  assign n2074 = ~n3173 & n3175;
  assign n2075 = x27 & x40;
  assign n2076 = n2074 & n2075;
  assign n2077 = n2074 | n2075;
  assign n2078 = ~n2076 & n2077;
  assign n3176 = n1979 & n2078;
  assign n3177 = (n2078 & n3136) | (n2078 & n3176) | (n3136 & n3176);
  assign n3178 = n1979 | n2078;
  assign n3179 = n3136 | n3178;
  assign n2081 = ~n3177 & n3179;
  assign n2082 = x26 & x41;
  assign n2083 = n2081 & n2082;
  assign n2084 = n2081 | n2082;
  assign n2085 = ~n2083 & n2084;
  assign n3180 = n1986 & n2085;
  assign n3181 = (n2085 & n3140) | (n2085 & n3180) | (n3140 & n3180);
  assign n3182 = n1986 | n2085;
  assign n3183 = n3140 | n3182;
  assign n2088 = ~n3181 & n3183;
  assign n2089 = x25 & x42;
  assign n2090 = n2088 & n2089;
  assign n2091 = n2088 | n2089;
  assign n2092 = ~n2090 & n2091;
  assign n2093 = n3148 & n2092;
  assign n2094 = n3148 | n2092;
  assign n2095 = ~n2093 & n2094;
  assign n2096 = x24 & x43;
  assign n2097 = n2095 & n2096;
  assign n2098 = n2095 | n2096;
  assign n2099 = ~n2097 & n2098;
  assign n2100 = n3146 & n2099;
  assign n2101 = n3146 | n2099;
  assign n2102 = ~n2100 & n2101;
  assign n2103 = x23 & x44;
  assign n2104 = n2102 & n2103;
  assign n2105 = n2102 | n2103;
  assign n2106 = ~n2104 & n2105;
  assign n2107 = n3144 & n2106;
  assign n2108 = n3144 | n2106;
  assign n2109 = ~n2107 & n2108;
  assign n2110 = x22 & x45;
  assign n2111 = n2109 & n2110;
  assign n2112 = n2109 | n2110;
  assign n2113 = ~n2111 & n2112;
  assign n2114 = n2036 & n2113;
  assign n2115 = n2036 | n2113;
  assign n2116 = ~n2114 & n2115;
  assign n2117 = x21 & x46;
  assign n2118 = n2116 & n2117;
  assign n2119 = n2116 | n2117;
  assign n2120 = ~n2118 & n2119;
  assign n2121 = n2035 & n2120;
  assign n2122 = n2035 | n2120;
  assign n2123 = ~n2121 & n2122;
  assign n2124 = x20 & x47;
  assign n2125 = n2123 & n2124;
  assign n2126 = n2123 | n2124;
  assign n2127 = ~n2125 & n2126;
  assign n2128 = n2034 & n2127;
  assign n2129 = n2034 | n2127;
  assign n2130 = ~n2128 & n2129;
  assign n2131 = n2125 | n2128;
  assign n2132 = n2118 | n2121;
  assign n3184 = n2111 | n2113;
  assign n3185 = (n2036 & n2111) | (n2036 & n3184) | (n2111 & n3184);
  assign n3186 = n2104 | n2106;
  assign n3187 = (n2104 & n3144) | (n2104 & n3186) | (n3144 & n3186);
  assign n3188 = n2097 | n2099;
  assign n3189 = (n2097 & n3146) | (n2097 & n3188) | (n3146 & n3188);
  assign n3190 = n2090 | n2092;
  assign n3191 = (n2090 & n3148) | (n2090 & n3190) | (n3148 & n3190);
  assign n3195 = n2055 | n2057;
  assign n3711 = n1958 | n2055;
  assign n3712 = (n2055 & n2057) | (n2055 & n3711) | (n2057 & n3711);
  assign n3713 = (n3122 & n3195) | (n3122 & n3712) | (n3195 & n3712);
  assign n3714 = (n3121 & n3195) | (n3121 & n3712) | (n3195 & n3712);
  assign n3715 = (n3646 & n3713) | (n3646 & n3714) | (n3713 & n3714);
  assign n2143 = x31 & x37;
  assign n3197 = n2143 & n3697;
  assign n3716 = (n2143 & n3197) | (n2143 & n3703) | (n3197 & n3703);
  assign n3934 = (n2050 & n2143) | (n2050 & n3197) | (n2143 & n3197);
  assign n11956 = n2143 & n3697;
  assign n3936 = (n1951 & n3934) | (n1951 & n11956) | (n3934 & n11956);
  assign n3718 = (n3661 & n3716) | (n3661 & n3936) | (n3716 & n3936);
  assign n3199 = n2143 | n3697;
  assign n3719 = n3199 | n3703;
  assign n3937 = n2050 | n3199;
  assign n3938 = (n1951 & n3199) | (n1951 & n3937) | (n3199 & n3937);
  assign n3721 = (n3661 & n3719) | (n3661 & n3938) | (n3719 & n3938);
  assign n2146 = ~n3718 & n3721;
  assign n2147 = n3715 & n2146;
  assign n2148 = n3715 | n2146;
  assign n2149 = ~n2147 & n2148;
  assign n2150 = x30 & x38;
  assign n2151 = n2149 & n2150;
  assign n2152 = n2149 | n2150;
  assign n2153 = ~n2151 & n2152;
  assign n3192 = n2062 | n2064;
  assign n3201 = n2153 & n3192;
  assign n3202 = n2062 & n2153;
  assign n3203 = (n3692 & n3201) | (n3692 & n3202) | (n3201 & n3202);
  assign n3204 = n2153 | n3192;
  assign n3205 = n2062 | n2153;
  assign n3206 = (n3692 & n3204) | (n3692 & n3205) | (n3204 & n3205);
  assign n2156 = ~n3203 & n3206;
  assign n2157 = x29 & x39;
  assign n2158 = n2156 & n2157;
  assign n2159 = n2156 | n2157;
  assign n2160 = ~n2158 & n2159;
  assign n3207 = n2069 & n2160;
  assign n3722 = (n2160 & n3172) | (n2160 & n3207) | (n3172 & n3207);
  assign n3723 = (n2071 & n2160) | (n2071 & n3207) | (n2160 & n3207);
  assign n3724 = (n3132 & n3722) | (n3132 & n3723) | (n3722 & n3723);
  assign n3209 = n2069 | n2160;
  assign n3725 = n3172 | n3209;
  assign n3726 = n2071 | n3209;
  assign n3727 = (n3132 & n3725) | (n3132 & n3726) | (n3725 & n3726);
  assign n2163 = ~n3724 & n3727;
  assign n2164 = x28 & x40;
  assign n2165 = n2163 & n2164;
  assign n2166 = n2163 | n2164;
  assign n2167 = ~n2165 & n2166;
  assign n3211 = n2076 & n2167;
  assign n3212 = (n2167 & n3177) | (n2167 & n3211) | (n3177 & n3211);
  assign n3213 = n2076 | n2167;
  assign n3214 = n3177 | n3213;
  assign n2170 = ~n3212 & n3214;
  assign n2171 = x27 & x41;
  assign n2172 = n2170 & n2171;
  assign n2173 = n2170 | n2171;
  assign n2174 = ~n2172 & n2173;
  assign n3215 = n2083 & n2174;
  assign n3216 = (n2174 & n3181) | (n2174 & n3215) | (n3181 & n3215);
  assign n3217 = n2083 | n2174;
  assign n3218 = n3181 | n3217;
  assign n2177 = ~n3216 & n3218;
  assign n2178 = x26 & x42;
  assign n2179 = n2177 & n2178;
  assign n2180 = n2177 | n2178;
  assign n2181 = ~n2179 & n2180;
  assign n2182 = n3191 & n2181;
  assign n2183 = n3191 | n2181;
  assign n2184 = ~n2182 & n2183;
  assign n2185 = x25 & x43;
  assign n2186 = n2184 & n2185;
  assign n2187 = n2184 | n2185;
  assign n2188 = ~n2186 & n2187;
  assign n2189 = n3189 & n2188;
  assign n2190 = n3189 | n2188;
  assign n2191 = ~n2189 & n2190;
  assign n2192 = x24 & x44;
  assign n2193 = n2191 & n2192;
  assign n2194 = n2191 | n2192;
  assign n2195 = ~n2193 & n2194;
  assign n2196 = n3187 & n2195;
  assign n2197 = n3187 | n2195;
  assign n2198 = ~n2196 & n2197;
  assign n2199 = x23 & x45;
  assign n2200 = n2198 & n2199;
  assign n2201 = n2198 | n2199;
  assign n2202 = ~n2200 & n2201;
  assign n2203 = n3185 & n2202;
  assign n2204 = n3185 | n2202;
  assign n2205 = ~n2203 & n2204;
  assign n2206 = x22 & x46;
  assign n2207 = n2205 & n2206;
  assign n2208 = n2205 | n2206;
  assign n2209 = ~n2207 & n2208;
  assign n2210 = n2132 & n2209;
  assign n2211 = n2132 | n2209;
  assign n2212 = ~n2210 & n2211;
  assign n2213 = x21 & x47;
  assign n2214 = n2212 & n2213;
  assign n2215 = n2212 | n2213;
  assign n2216 = ~n2214 & n2215;
  assign n2217 = n2131 & n2216;
  assign n2218 = n2131 | n2216;
  assign n2219 = ~n2217 & n2218;
  assign n2220 = n2214 | n2217;
  assign n3219 = n2207 | n2209;
  assign n3220 = (n2132 & n2207) | (n2132 & n3219) | (n2207 & n3219);
  assign n3221 = n2200 | n2202;
  assign n3222 = (n2200 & n3185) | (n2200 & n3221) | (n3185 & n3221);
  assign n3223 = n2193 | n2195;
  assign n3224 = (n2193 & n3187) | (n2193 & n3223) | (n3187 & n3223);
  assign n3225 = n2186 | n2188;
  assign n3226 = (n2186 & n3189) | (n2186 & n3225) | (n3189 & n3225);
  assign n3227 = n2179 | n2181;
  assign n3228 = (n2179 & n3191) | (n2179 & n3227) | (n3191 & n3227);
  assign n3230 = n2158 | n2160;
  assign n3728 = n2069 | n2158;
  assign n3729 = (n2158 & n2160) | (n2158 & n3728) | (n2160 & n3728);
  assign n3730 = (n3172 & n3230) | (n3172 & n3729) | (n3230 & n3729);
  assign n3731 = (n2071 & n3230) | (n2071 & n3729) | (n3230 & n3729);
  assign n3732 = (n3132 & n3730) | (n3132 & n3731) | (n3730 & n3731);
  assign n2231 = x31 & x38;
  assign n3942 = n2143 & n2231;
  assign n11957 = n3697 & n3942;
  assign n3943 = (n3703 & n11957) | (n3703 & n3942) | (n11957 & n3942);
  assign n3939 = n2231 & n3936;
  assign n3940 = (n3661 & n3943) | (n3661 & n3939) | (n3943 & n3939);
  assign n3734 = (n2146 & n2231) | (n2146 & n3940) | (n2231 & n3940);
  assign n3736 = n2231 & n3936;
  assign n3737 = (n3661 & n3943) | (n3661 & n3736) | (n3943 & n3736);
  assign n3236 = (n3715 & n3734) | (n3715 & n3737) | (n3734 & n3737);
  assign n3947 = n2143 | n2231;
  assign n11958 = (n2231 & n3697) | (n2231 & n3947) | (n3697 & n3947);
  assign n3948 = (n3703 & n11958) | (n3703 & n3947) | (n11958 & n3947);
  assign n3944 = n2231 | n3936;
  assign n3945 = (n3661 & n3948) | (n3661 & n3944) | (n3948 & n3944);
  assign n3739 = n2146 | n3945;
  assign n3741 = n2231 | n3936;
  assign n3742 = (n3661 & n3948) | (n3661 & n3741) | (n3948 & n3741);
  assign n3239 = (n3715 & n3739) | (n3715 & n3742) | (n3739 & n3742);
  assign n2234 = ~n3236 & n3239;
  assign n3240 = n2151 & n2234;
  assign n3743 = (n2234 & n3202) | (n2234 & n3240) | (n3202 & n3240);
  assign n3744 = (n2234 & n3201) | (n2234 & n3240) | (n3201 & n3240);
  assign n3745 = (n3692 & n3743) | (n3692 & n3744) | (n3743 & n3744);
  assign n3242 = n2151 | n2234;
  assign n3746 = n3202 | n3242;
  assign n3747 = n3201 | n3242;
  assign n3748 = (n3692 & n3746) | (n3692 & n3747) | (n3746 & n3747);
  assign n2237 = ~n3745 & n3748;
  assign n2238 = x30 & x39;
  assign n2239 = n2237 & n2238;
  assign n2240 = n2237 | n2238;
  assign n2241 = ~n2239 & n2240;
  assign n2242 = n3732 & n2241;
  assign n2243 = n3732 | n2241;
  assign n2244 = ~n2242 & n2243;
  assign n2245 = x29 & x40;
  assign n2246 = n2244 & n2245;
  assign n2247 = n2244 | n2245;
  assign n2248 = ~n2246 & n2247;
  assign n3244 = n2165 & n2248;
  assign n3245 = (n2248 & n3212) | (n2248 & n3244) | (n3212 & n3244);
  assign n3246 = n2165 | n2248;
  assign n3247 = n3212 | n3246;
  assign n2251 = ~n3245 & n3247;
  assign n2252 = x28 & x41;
  assign n2253 = n2251 & n2252;
  assign n2254 = n2251 | n2252;
  assign n2255 = ~n2253 & n2254;
  assign n3248 = n2172 & n2255;
  assign n3249 = (n2255 & n3216) | (n2255 & n3248) | (n3216 & n3248);
  assign n3250 = n2172 | n2255;
  assign n3251 = n3216 | n3250;
  assign n2258 = ~n3249 & n3251;
  assign n2259 = x27 & x42;
  assign n2260 = n2258 & n2259;
  assign n2261 = n2258 | n2259;
  assign n2262 = ~n2260 & n2261;
  assign n2263 = n3228 & n2262;
  assign n2264 = n3228 | n2262;
  assign n2265 = ~n2263 & n2264;
  assign n2266 = x26 & x43;
  assign n2267 = n2265 & n2266;
  assign n2268 = n2265 | n2266;
  assign n2269 = ~n2267 & n2268;
  assign n2270 = n3226 & n2269;
  assign n2271 = n3226 | n2269;
  assign n2272 = ~n2270 & n2271;
  assign n2273 = x25 & x44;
  assign n2274 = n2272 & n2273;
  assign n2275 = n2272 | n2273;
  assign n2276 = ~n2274 & n2275;
  assign n2277 = n3224 & n2276;
  assign n2278 = n3224 | n2276;
  assign n2279 = ~n2277 & n2278;
  assign n2280 = x24 & x45;
  assign n2281 = n2279 & n2280;
  assign n2282 = n2279 | n2280;
  assign n2283 = ~n2281 & n2282;
  assign n2284 = n3222 & n2283;
  assign n2285 = n3222 | n2283;
  assign n2286 = ~n2284 & n2285;
  assign n2287 = x23 & x46;
  assign n2288 = n2286 & n2287;
  assign n2289 = n2286 | n2287;
  assign n2290 = ~n2288 & n2289;
  assign n2291 = n3220 & n2290;
  assign n2292 = n3220 | n2290;
  assign n2293 = ~n2291 & n2292;
  assign n2294 = x22 & x47;
  assign n2295 = n2293 & n2294;
  assign n2296 = n2293 | n2294;
  assign n2297 = ~n2295 & n2296;
  assign n2298 = n2220 & n2297;
  assign n2299 = n2220 | n2297;
  assign n2300 = ~n2298 & n2299;
  assign n3252 = n2295 | n2297;
  assign n3253 = (n2220 & n2295) | (n2220 & n3252) | (n2295 & n3252);
  assign n3254 = n2288 | n2290;
  assign n3255 = (n2288 & n3220) | (n2288 & n3254) | (n3220 & n3254);
  assign n3256 = n2281 | n2283;
  assign n3257 = (n2281 & n3222) | (n2281 & n3256) | (n3222 & n3256);
  assign n3258 = n2274 | n2276;
  assign n3259 = (n2274 & n3224) | (n2274 & n3258) | (n3224 & n3258);
  assign n3260 = n2267 | n2269;
  assign n3261 = (n2267 & n3226) | (n2267 & n3260) | (n3226 & n3260);
  assign n3262 = n2260 | n2262;
  assign n3263 = (n2260 & n3228) | (n2260 & n3262) | (n3228 & n3262);
  assign n2311 = x31 & x39;
  assign n3267 = n2234 | n3236;
  assign n3749 = (n2151 & n3236) | (n2151 & n3267) | (n3236 & n3267);
  assign n3269 = n2311 & n3749;
  assign n15589 = n2311 & n3942;
  assign n17670 = n3697 & n15589;
  assign n15590 = (n3703 & n17670) | (n3703 & n15589) | (n17670 & n15589);
  assign n11960 = n2231 & n2311;
  assign n15591 = n3936 & n11960;
  assign n15587 = (n3661 & n15590) | (n3661 & n15591) | (n15590 & n15591);
  assign n11961 = (n2146 & n15587) | (n2146 & n11960) | (n15587 & n11960);
  assign n11964 = (n3661 & n15590) | (n3661 & n15591) | (n15590 & n15591);
  assign n3951 = (n3715 & n11961) | (n3715 & n11964) | (n11961 & n11964);
  assign n3751 = (n2234 & n2311) | (n2234 & n3951) | (n2311 & n3951);
  assign n3752 = (n3202 & n3269) | (n3202 & n3751) | (n3269 & n3751);
  assign n3753 = (n3201 & n3269) | (n3201 & n3751) | (n3269 & n3751);
  assign n3754 = (n3692 & n3752) | (n3692 & n3753) | (n3752 & n3753);
  assign n3272 = n2311 | n3749;
  assign n15595 = n2311 | n3942;
  assign n17671 = (n2311 & n3697) | (n2311 & n15595) | (n3697 & n15595);
  assign n15596 = (n3703 & n17671) | (n3703 & n15595) | (n17671 & n15595);
  assign n11966 = n2231 | n2311;
  assign n15597 = (n2311 & n3936) | (n2311 & n11966) | (n3936 & n11966);
  assign n15593 = (n3661 & n15596) | (n3661 & n15597) | (n15596 & n15597);
  assign n11967 = (n2146 & n15593) | (n2146 & n11966) | (n15593 & n11966);
  assign n11970 = (n3661 & n15596) | (n3661 & n15597) | (n15596 & n15597);
  assign n3954 = (n3715 & n11967) | (n3715 & n11970) | (n11967 & n11970);
  assign n3756 = n2234 | n3954;
  assign n3757 = (n3202 & n3272) | (n3202 & n3756) | (n3272 & n3756);
  assign n3758 = (n3201 & n3272) | (n3201 & n3756) | (n3272 & n3756);
  assign n3759 = (n3692 & n3757) | (n3692 & n3758) | (n3757 & n3758);
  assign n2314 = ~n3754 & n3759;
  assign n3276 = n2239 & n2314;
  assign n3760 = (n2241 & n2314) | (n2241 & n3276) | (n2314 & n3276);
  assign n3277 = (n3732 & n3760) | (n3732 & n3276) | (n3760 & n3276);
  assign n3279 = n2239 | n2314;
  assign n3761 = n2241 | n3279;
  assign n3280 = (n3732 & n3761) | (n3732 & n3279) | (n3761 & n3279);
  assign n2317 = ~n3277 & n3280;
  assign n2318 = x30 & x40;
  assign n2319 = n2317 & n2318;
  assign n2320 = n2317 | n2318;
  assign n2321 = ~n2319 & n2320;
  assign n3281 = n2246 & n2321;
  assign n3762 = (n2321 & n3244) | (n2321 & n3281) | (n3244 & n3281);
  assign n3763 = (n2248 & n2321) | (n2248 & n3281) | (n2321 & n3281);
  assign n3764 = (n3212 & n3762) | (n3212 & n3763) | (n3762 & n3763);
  assign n3283 = n2246 | n2321;
  assign n3765 = n3244 | n3283;
  assign n3766 = n2248 | n3283;
  assign n3767 = (n3212 & n3765) | (n3212 & n3766) | (n3765 & n3766);
  assign n2324 = ~n3764 & n3767;
  assign n2325 = x29 & x41;
  assign n2326 = n2324 & n2325;
  assign n2327 = n2324 | n2325;
  assign n2328 = ~n2326 & n2327;
  assign n3285 = n2253 & n2328;
  assign n3286 = (n2328 & n3249) | (n2328 & n3285) | (n3249 & n3285);
  assign n3287 = n2253 | n2328;
  assign n3288 = n3249 | n3287;
  assign n2331 = ~n3286 & n3288;
  assign n2332 = x28 & x42;
  assign n2333 = n2331 & n2332;
  assign n2334 = n2331 | n2332;
  assign n2335 = ~n2333 & n2334;
  assign n2336 = n3263 & n2335;
  assign n2337 = n3263 | n2335;
  assign n2338 = ~n2336 & n2337;
  assign n2339 = x27 & x43;
  assign n2340 = n2338 & n2339;
  assign n2341 = n2338 | n2339;
  assign n2342 = ~n2340 & n2341;
  assign n2343 = n3261 & n2342;
  assign n2344 = n3261 | n2342;
  assign n2345 = ~n2343 & n2344;
  assign n2346 = x26 & x44;
  assign n2347 = n2345 & n2346;
  assign n2348 = n2345 | n2346;
  assign n2349 = ~n2347 & n2348;
  assign n2350 = n3259 & n2349;
  assign n2351 = n3259 | n2349;
  assign n2352 = ~n2350 & n2351;
  assign n2353 = x25 & x45;
  assign n2354 = n2352 & n2353;
  assign n2355 = n2352 | n2353;
  assign n2356 = ~n2354 & n2355;
  assign n2357 = n3257 & n2356;
  assign n2358 = n3257 | n2356;
  assign n2359 = ~n2357 & n2358;
  assign n2360 = x24 & x46;
  assign n2361 = n2359 & n2360;
  assign n2362 = n2359 | n2360;
  assign n2363 = ~n2361 & n2362;
  assign n2364 = n3255 & n2363;
  assign n2365 = n3255 | n2363;
  assign n2366 = ~n2364 & n2365;
  assign n2367 = x23 & x47;
  assign n2368 = n2366 & n2367;
  assign n2369 = n2366 | n2367;
  assign n2370 = ~n2368 & n2369;
  assign n2371 = n3253 & n2370;
  assign n2372 = n3253 | n2370;
  assign n2373 = ~n2371 & n2372;
  assign n3289 = n2368 | n2370;
  assign n3290 = (n2368 & n3253) | (n2368 & n3289) | (n3253 & n3289);
  assign n3291 = n2361 | n2363;
  assign n3292 = (n2361 & n3255) | (n2361 & n3291) | (n3255 & n3291);
  assign n3293 = n2354 | n2356;
  assign n3294 = (n2354 & n3257) | (n2354 & n3293) | (n3257 & n3293);
  assign n3295 = n2347 | n2349;
  assign n3296 = (n2347 & n3259) | (n2347 & n3295) | (n3259 & n3295);
  assign n3297 = n2340 | n2342;
  assign n3298 = (n2340 & n3261) | (n2340 & n3297) | (n3261 & n3297);
  assign n3299 = n2333 | n2335;
  assign n3300 = (n2333 & n3263) | (n2333 & n3299) | (n3263 & n3299);
  assign n3302 = n2319 | n2321;
  assign n3768 = n2246 | n2319;
  assign n3769 = (n2319 & n2321) | (n2319 & n3768) | (n2321 & n3768);
  assign n3770 = (n3244 & n3302) | (n3244 & n3769) | (n3302 & n3769);
  assign n3771 = (n2248 & n3302) | (n2248 & n3769) | (n3302 & n3769);
  assign n3772 = (n3212 & n3770) | (n3212 & n3771) | (n3770 & n3771);
  assign n2383 = x31 & x40;
  assign n3304 = n2383 & n3754;
  assign n3773 = (n2383 & n3304) | (n2383 & n3760) | (n3304 & n3760);
  assign n3955 = (n2314 & n2383) | (n2314 & n3304) | (n2383 & n3304);
  assign n11971 = n2383 & n3754;
  assign n3957 = (n2239 & n3955) | (n2239 & n11971) | (n3955 & n11971);
  assign n3775 = (n3732 & n3773) | (n3732 & n3957) | (n3773 & n3957);
  assign n3306 = n2383 | n3754;
  assign n3776 = n3306 | n3760;
  assign n3958 = n2314 | n3306;
  assign n3959 = (n2239 & n3306) | (n2239 & n3958) | (n3306 & n3958);
  assign n3778 = (n3732 & n3776) | (n3732 & n3959) | (n3776 & n3959);
  assign n2386 = ~n3775 & n3778;
  assign n2387 = n3772 & n2386;
  assign n2388 = n3772 | n2386;
  assign n2389 = ~n2387 & n2388;
  assign n2390 = x30 & x41;
  assign n2391 = n2389 & n2390;
  assign n2392 = n2389 | n2390;
  assign n2393 = ~n2391 & n2392;
  assign n3308 = n2326 & n2393;
  assign n3309 = (n2393 & n3286) | (n2393 & n3308) | (n3286 & n3308);
  assign n3310 = n2326 | n2393;
  assign n3311 = n3286 | n3310;
  assign n2396 = ~n3309 & n3311;
  assign n2397 = x29 & x42;
  assign n2398 = n2396 & n2397;
  assign n2399 = n2396 | n2397;
  assign n2400 = ~n2398 & n2399;
  assign n2401 = n3300 & n2400;
  assign n2402 = n3300 | n2400;
  assign n2403 = ~n2401 & n2402;
  assign n2404 = x28 & x43;
  assign n2405 = n2403 & n2404;
  assign n2406 = n2403 | n2404;
  assign n2407 = ~n2405 & n2406;
  assign n2408 = n3298 & n2407;
  assign n2409 = n3298 | n2407;
  assign n2410 = ~n2408 & n2409;
  assign n2411 = x27 & x44;
  assign n2412 = n2410 & n2411;
  assign n2413 = n2410 | n2411;
  assign n2414 = ~n2412 & n2413;
  assign n2415 = n3296 & n2414;
  assign n2416 = n3296 | n2414;
  assign n2417 = ~n2415 & n2416;
  assign n2418 = x26 & x45;
  assign n2419 = n2417 & n2418;
  assign n2420 = n2417 | n2418;
  assign n2421 = ~n2419 & n2420;
  assign n2422 = n3294 & n2421;
  assign n2423 = n3294 | n2421;
  assign n2424 = ~n2422 & n2423;
  assign n2425 = x25 & x46;
  assign n2426 = n2424 & n2425;
  assign n2427 = n2424 | n2425;
  assign n2428 = ~n2426 & n2427;
  assign n2429 = n3292 & n2428;
  assign n2430 = n3292 | n2428;
  assign n2431 = ~n2429 & n2430;
  assign n2432 = x24 & x47;
  assign n2433 = n2431 & n2432;
  assign n2434 = n2431 | n2432;
  assign n2435 = ~n2433 & n2434;
  assign n2436 = n3290 & n2435;
  assign n2437 = n3290 | n2435;
  assign n2438 = ~n2436 & n2437;
  assign n3312 = n2433 | n2435;
  assign n3313 = (n2433 & n3290) | (n2433 & n3312) | (n3290 & n3312);
  assign n3314 = n2426 | n2428;
  assign n3315 = (n2426 & n3292) | (n2426 & n3314) | (n3292 & n3314);
  assign n3316 = n2419 | n2421;
  assign n3317 = (n2419 & n3294) | (n2419 & n3316) | (n3294 & n3316);
  assign n3318 = n2412 | n2414;
  assign n3319 = (n2412 & n3296) | (n2412 & n3318) | (n3296 & n3318);
  assign n3320 = n2405 | n2407;
  assign n3321 = (n2405 & n3298) | (n2405 & n3320) | (n3298 & n3320);
  assign n3322 = n2398 | n2400;
  assign n3323 = (n2398 & n3300) | (n2398 & n3322) | (n3300 & n3322);
  assign n2447 = x31 & x41;
  assign n3963 = n2383 & n2447;
  assign n11972 = n3754 & n3963;
  assign n3964 = (n3760 & n11972) | (n3760 & n3963) | (n11972 & n3963);
  assign n3960 = n2447 & n3957;
  assign n3961 = (n3732 & n3964) | (n3732 & n3960) | (n3964 & n3960);
  assign n3780 = (n2386 & n2447) | (n2386 & n3961) | (n2447 & n3961);
  assign n3782 = n2447 & n3957;
  assign n3783 = (n3732 & n3964) | (n3732 & n3782) | (n3964 & n3782);
  assign n3328 = (n3772 & n3780) | (n3772 & n3783) | (n3780 & n3783);
  assign n3968 = n2383 | n2447;
  assign n11973 = (n2447 & n3754) | (n2447 & n3968) | (n3754 & n3968);
  assign n3969 = (n3760 & n11973) | (n3760 & n3968) | (n11973 & n3968);
  assign n3965 = n2447 | n3957;
  assign n3966 = (n3732 & n3969) | (n3732 & n3965) | (n3969 & n3965);
  assign n3785 = n2386 | n3966;
  assign n3787 = n2447 | n3957;
  assign n3788 = (n3732 & n3969) | (n3732 & n3787) | (n3969 & n3787);
  assign n3331 = (n3772 & n3785) | (n3772 & n3788) | (n3785 & n3788);
  assign n2450 = ~n3328 & n3331;
  assign n3332 = n2391 & n2450;
  assign n3789 = (n2450 & n3308) | (n2450 & n3332) | (n3308 & n3332);
  assign n3790 = (n2393 & n2450) | (n2393 & n3332) | (n2450 & n3332);
  assign n3791 = (n3286 & n3789) | (n3286 & n3790) | (n3789 & n3790);
  assign n3334 = n2391 | n2450;
  assign n3792 = n3308 | n3334;
  assign n3793 = n2393 | n3334;
  assign n3794 = (n3286 & n3792) | (n3286 & n3793) | (n3792 & n3793);
  assign n2453 = ~n3791 & n3794;
  assign n2454 = x30 & x42;
  assign n2455 = n2453 & n2454;
  assign n2456 = n2453 | n2454;
  assign n2457 = ~n2455 & n2456;
  assign n2458 = n3323 & n2457;
  assign n2459 = n3323 | n2457;
  assign n2460 = ~n2458 & n2459;
  assign n2461 = x29 & x43;
  assign n2462 = n2460 & n2461;
  assign n2463 = n2460 | n2461;
  assign n2464 = ~n2462 & n2463;
  assign n2465 = n3321 & n2464;
  assign n2466 = n3321 | n2464;
  assign n2467 = ~n2465 & n2466;
  assign n2468 = x28 & x44;
  assign n2469 = n2467 & n2468;
  assign n2470 = n2467 | n2468;
  assign n2471 = ~n2469 & n2470;
  assign n2472 = n3319 & n2471;
  assign n2473 = n3319 | n2471;
  assign n2474 = ~n2472 & n2473;
  assign n2475 = x27 & x45;
  assign n2476 = n2474 & n2475;
  assign n2477 = n2474 | n2475;
  assign n2478 = ~n2476 & n2477;
  assign n2479 = n3317 & n2478;
  assign n2480 = n3317 | n2478;
  assign n2481 = ~n2479 & n2480;
  assign n2482 = x26 & x46;
  assign n2483 = n2481 & n2482;
  assign n2484 = n2481 | n2482;
  assign n2485 = ~n2483 & n2484;
  assign n2486 = n3315 & n2485;
  assign n2487 = n3315 | n2485;
  assign n2488 = ~n2486 & n2487;
  assign n2489 = x25 & x47;
  assign n2490 = n2488 & n2489;
  assign n2491 = n2488 | n2489;
  assign n2492 = ~n2490 & n2491;
  assign n2493 = n3313 & n2492;
  assign n2494 = n3313 | n2492;
  assign n2495 = ~n2493 & n2494;
  assign n3336 = n2490 | n2492;
  assign n3337 = (n2490 & n3313) | (n2490 & n3336) | (n3313 & n3336);
  assign n3338 = n2483 | n2485;
  assign n3339 = (n2483 & n3315) | (n2483 & n3338) | (n3315 & n3338);
  assign n3340 = n2476 | n2478;
  assign n3341 = (n2476 & n3317) | (n2476 & n3340) | (n3317 & n3340);
  assign n3342 = n2469 | n2471;
  assign n3343 = (n2469 & n3319) | (n2469 & n3342) | (n3319 & n3342);
  assign n3344 = n2462 | n2464;
  assign n3345 = (n2462 & n3321) | (n2462 & n3344) | (n3321 & n3344);
  assign n2503 = x31 & x42;
  assign n3349 = n2450 | n3328;
  assign n3795 = (n2391 & n3328) | (n2391 & n3349) | (n3328 & n3349);
  assign n3351 = n2503 & n3795;
  assign n15601 = n2503 & n3963;
  assign n17672 = n3754 & n15601;
  assign n15602 = (n3760 & n17672) | (n3760 & n15601) | (n17672 & n15601);
  assign n11975 = n2447 & n2503;
  assign n15603 = n3957 & n11975;
  assign n15599 = (n3732 & n15602) | (n3732 & n15603) | (n15602 & n15603);
  assign n11976 = (n2386 & n15599) | (n2386 & n11975) | (n15599 & n11975);
  assign n11979 = (n3732 & n15602) | (n3732 & n15603) | (n15602 & n15603);
  assign n3972 = (n3772 & n11976) | (n3772 & n11979) | (n11976 & n11979);
  assign n3797 = (n2450 & n2503) | (n2450 & n3972) | (n2503 & n3972);
  assign n3798 = (n3308 & n3351) | (n3308 & n3797) | (n3351 & n3797);
  assign n3799 = (n2393 & n3351) | (n2393 & n3797) | (n3351 & n3797);
  assign n3800 = (n3286 & n3798) | (n3286 & n3799) | (n3798 & n3799);
  assign n3354 = n2503 | n3795;
  assign n15607 = n2503 | n3963;
  assign n17673 = (n2503 & n3754) | (n2503 & n15607) | (n3754 & n15607);
  assign n15608 = (n3760 & n17673) | (n3760 & n15607) | (n17673 & n15607);
  assign n11981 = n2447 | n2503;
  assign n15609 = (n2503 & n3957) | (n2503 & n11981) | (n3957 & n11981);
  assign n15605 = (n3732 & n15608) | (n3732 & n15609) | (n15608 & n15609);
  assign n11982 = (n2386 & n15605) | (n2386 & n11981) | (n15605 & n11981);
  assign n11985 = (n3732 & n15608) | (n3732 & n15609) | (n15608 & n15609);
  assign n3975 = (n3772 & n11982) | (n3772 & n11985) | (n11982 & n11985);
  assign n3802 = n2450 | n3975;
  assign n3803 = (n3308 & n3354) | (n3308 & n3802) | (n3354 & n3802);
  assign n3804 = (n2393 & n3354) | (n2393 & n3802) | (n3354 & n3802);
  assign n3805 = (n3286 & n3803) | (n3286 & n3804) | (n3803 & n3804);
  assign n2506 = ~n3800 & n3805;
  assign n3807 = n2455 & n2506;
  assign n3976 = (n2457 & n2506) | (n2457 & n3807) | (n2506 & n3807);
  assign n3808 = (n3323 & n3976) | (n3323 & n3807) | (n3976 & n3807);
  assign n3810 = n2455 | n2506;
  assign n3977 = n2457 | n3810;
  assign n3811 = (n3323 & n3977) | (n3323 & n3810) | (n3977 & n3810);
  assign n2509 = ~n3808 & n3811;
  assign n2510 = x30 & x43;
  assign n2511 = n2509 & n2510;
  assign n2512 = n2509 | n2510;
  assign n2513 = ~n2511 & n2512;
  assign n2514 = n3345 & n2513;
  assign n2515 = n3345 | n2513;
  assign n2516 = ~n2514 & n2515;
  assign n2517 = x29 & x44;
  assign n2518 = n2516 & n2517;
  assign n2519 = n2516 | n2517;
  assign n2520 = ~n2518 & n2519;
  assign n2521 = n3343 & n2520;
  assign n2522 = n3343 | n2520;
  assign n2523 = ~n2521 & n2522;
  assign n2524 = x28 & x45;
  assign n2525 = n2523 & n2524;
  assign n2526 = n2523 | n2524;
  assign n2527 = ~n2525 & n2526;
  assign n2528 = n3341 & n2527;
  assign n2529 = n3341 | n2527;
  assign n2530 = ~n2528 & n2529;
  assign n2531 = x27 & x46;
  assign n2532 = n2530 & n2531;
  assign n2533 = n2530 | n2531;
  assign n2534 = ~n2532 & n2533;
  assign n2535 = n3339 & n2534;
  assign n2536 = n3339 | n2534;
  assign n2537 = ~n2535 & n2536;
  assign n2538 = x26 & x47;
  assign n2539 = n2537 & n2538;
  assign n2540 = n2537 | n2538;
  assign n2541 = ~n2539 & n2540;
  assign n2542 = n3337 & n2541;
  assign n2543 = n3337 | n2541;
  assign n2544 = ~n2542 & n2543;
  assign n3357 = n2539 | n2541;
  assign n3358 = (n2539 & n3337) | (n2539 & n3357) | (n3337 & n3357);
  assign n3359 = n2532 | n2534;
  assign n3360 = (n2532 & n3339) | (n2532 & n3359) | (n3339 & n3359);
  assign n3361 = n2525 | n2527;
  assign n3362 = (n2525 & n3341) | (n2525 & n3361) | (n3341 & n3361);
  assign n3363 = n2518 | n2520;
  assign n3364 = (n2518 & n3343) | (n2518 & n3363) | (n3343 & n3363);
  assign n2551 = x31 & x43;
  assign n3370 = n2551 & n3800;
  assign n3812 = n2551 & n3800;
  assign n3813 = (n2506 & n2551) | (n2506 & n3812) | (n2551 & n3812);
  assign n3815 = (n2455 & n3370) | (n2455 & n3813) | (n3370 & n3813);
  assign n3978 = n3370 | n3813;
  assign n3979 = (n2457 & n3815) | (n2457 & n3978) | (n3815 & n3978);
  assign n3816 = (n3323 & n3979) | (n3323 & n3815) | (n3979 & n3815);
  assign n3373 = n2551 | n3800;
  assign n3817 = n2551 | n3800;
  assign n3818 = n2506 | n3817;
  assign n3820 = (n2455 & n3373) | (n2455 & n3818) | (n3373 & n3818);
  assign n3980 = n3373 | n3818;
  assign n3981 = (n2457 & n3820) | (n2457 & n3980) | (n3820 & n3980);
  assign n3821 = (n3323 & n3981) | (n3323 & n3820) | (n3981 & n3820);
  assign n2554 = ~n3816 & n3821;
  assign n3823 = n2511 & n2554;
  assign n3982 = (n2513 & n2554) | (n2513 & n3823) | (n2554 & n3823);
  assign n3824 = (n3345 & n3982) | (n3345 & n3823) | (n3982 & n3823);
  assign n3826 = n2511 | n2554;
  assign n3983 = n2513 | n3826;
  assign n3827 = (n3345 & n3983) | (n3345 & n3826) | (n3983 & n3826);
  assign n2557 = ~n3824 & n3827;
  assign n2558 = x30 & x44;
  assign n2559 = n2557 & n2558;
  assign n2560 = n2557 | n2558;
  assign n2561 = ~n2559 & n2560;
  assign n2562 = n3364 & n2561;
  assign n2563 = n3364 | n2561;
  assign n2564 = ~n2562 & n2563;
  assign n2565 = x29 & x45;
  assign n2566 = n2564 & n2565;
  assign n2567 = n2564 | n2565;
  assign n2568 = ~n2566 & n2567;
  assign n2569 = n3362 & n2568;
  assign n2570 = n3362 | n2568;
  assign n2571 = ~n2569 & n2570;
  assign n2572 = x28 & x46;
  assign n2573 = n2571 & n2572;
  assign n2574 = n2571 | n2572;
  assign n2575 = ~n2573 & n2574;
  assign n2576 = n3360 & n2575;
  assign n2577 = n3360 | n2575;
  assign n2578 = ~n2576 & n2577;
  assign n2579 = x27 & x47;
  assign n2580 = n2578 & n2579;
  assign n2581 = n2578 | n2579;
  assign n2582 = ~n2580 & n2581;
  assign n2583 = n3358 & n2582;
  assign n2584 = n3358 | n2582;
  assign n2585 = ~n2583 & n2584;
  assign n3375 = n2580 | n2582;
  assign n3376 = (n2580 & n3358) | (n2580 & n3375) | (n3358 & n3375);
  assign n3377 = n2573 | n2575;
  assign n3378 = (n2573 & n3360) | (n2573 & n3377) | (n3360 & n3377);
  assign n3379 = n2566 | n2568;
  assign n3380 = (n2566 & n3362) | (n2566 & n3379) | (n3362 & n3379);
  assign n2591 = x31 & x44;
  assign n3984 = n2591 & n3979;
  assign n3985 = n2591 & n3815;
  assign n3986 = (n3323 & n3984) | (n3323 & n3985) | (n3984 & n3985);
  assign n3829 = (n2554 & n2591) | (n2554 & n3986) | (n2591 & n3986);
  assign n3987 = (n2511 & n3829) | (n2511 & n3986) | (n3829 & n3986);
  assign n11986 = n2591 | n3986;
  assign n11987 = (n2554 & n3986) | (n2554 & n11986) | (n3986 & n11986);
  assign n3989 = (n2513 & n3987) | (n2513 & n11987) | (n3987 & n11987);
  assign n3831 = (n2511 & n3986) | (n2511 & n3829) | (n3986 & n3829);
  assign n3832 = (n3345 & n3989) | (n3345 & n3831) | (n3989 & n3831);
  assign n3990 = n2591 | n3979;
  assign n3991 = n2591 | n3815;
  assign n3992 = (n3323 & n3990) | (n3323 & n3991) | (n3990 & n3991);
  assign n3834 = n2554 | n3992;
  assign n3993 = (n2511 & n3834) | (n2511 & n3992) | (n3834 & n3992);
  assign n11988 = n2554 | n3992;
  assign n3995 = (n2513 & n3993) | (n2513 & n11988) | (n3993 & n11988);
  assign n3836 = (n2511 & n3992) | (n2511 & n3834) | (n3992 & n3834);
  assign n3837 = (n3345 & n3995) | (n3345 & n3836) | (n3995 & n3836);
  assign n2594 = ~n3832 & n3837;
  assign n3839 = n2559 & n2594;
  assign n3996 = (n2561 & n2594) | (n2561 & n3839) | (n2594 & n3839);
  assign n3840 = (n3364 & n3996) | (n3364 & n3839) | (n3996 & n3839);
  assign n3842 = n2559 | n2594;
  assign n3997 = n2561 | n3842;
  assign n3843 = (n3364 & n3997) | (n3364 & n3842) | (n3997 & n3842);
  assign n2597 = ~n3840 & n3843;
  assign n2598 = x30 & x45;
  assign n2599 = n2597 & n2598;
  assign n2600 = n2597 | n2598;
  assign n2601 = ~n2599 & n2600;
  assign n2602 = n3380 & n2601;
  assign n2603 = n3380 | n2601;
  assign n2604 = ~n2602 & n2603;
  assign n2605 = x29 & x46;
  assign n2606 = n2604 & n2605;
  assign n2607 = n2604 | n2605;
  assign n2608 = ~n2606 & n2607;
  assign n2609 = n3378 & n2608;
  assign n2610 = n3378 | n2608;
  assign n2611 = ~n2609 & n2610;
  assign n2612 = x28 & x47;
  assign n2613 = n2611 & n2612;
  assign n2614 = n2611 | n2612;
  assign n2615 = ~n2613 & n2614;
  assign n2616 = n3376 & n2615;
  assign n2617 = n3376 | n2615;
  assign n2618 = ~n2616 & n2617;
  assign n3391 = n2613 | n2615;
  assign n3392 = (n2613 & n3376) | (n2613 & n3391) | (n3376 & n3391);
  assign n3393 = n2606 | n2608;
  assign n3394 = (n2606 & n3378) | (n2606 & n3393) | (n3378 & n3393);
  assign n2623 = x31 & x45;
  assign n3998 = n2623 & n3989;
  assign n3999 = n2623 & n3831;
  assign n4000 = (n3345 & n3998) | (n3345 & n3999) | (n3998 & n3999);
  assign n3845 = (n2594 & n2623) | (n2594 & n4000) | (n2623 & n4000);
  assign n4001 = (n2559 & n3845) | (n2559 & n4000) | (n3845 & n4000);
  assign n11989 = n2623 | n4000;
  assign n11990 = (n2594 & n4000) | (n2594 & n11989) | (n4000 & n11989);
  assign n4003 = (n2561 & n4001) | (n2561 & n11990) | (n4001 & n11990);
  assign n3847 = (n2559 & n4000) | (n2559 & n3845) | (n4000 & n3845);
  assign n3848 = (n3364 & n4003) | (n3364 & n3847) | (n4003 & n3847);
  assign n4004 = n2623 | n3989;
  assign n4005 = n2623 | n3831;
  assign n4006 = (n3345 & n4004) | (n3345 & n4005) | (n4004 & n4005);
  assign n3850 = n2594 | n4006;
  assign n4007 = (n2559 & n3850) | (n2559 & n4006) | (n3850 & n4006);
  assign n11991 = n2594 | n4006;
  assign n4009 = (n2561 & n4007) | (n2561 & n11991) | (n4007 & n11991);
  assign n3852 = (n2559 & n4006) | (n2559 & n3850) | (n4006 & n3850);
  assign n3853 = (n3364 & n4009) | (n3364 & n3852) | (n4009 & n3852);
  assign n2626 = ~n3848 & n3853;
  assign n3855 = n2599 & n2626;
  assign n4010 = (n2601 & n2626) | (n2601 & n3855) | (n2626 & n3855);
  assign n3856 = (n3380 & n4010) | (n3380 & n3855) | (n4010 & n3855);
  assign n3858 = n2599 | n2626;
  assign n4011 = n2601 | n3858;
  assign n3859 = (n3380 & n4011) | (n3380 & n3858) | (n4011 & n3858);
  assign n2629 = ~n3856 & n3859;
  assign n2630 = x30 & x46;
  assign n2631 = n2629 & n2630;
  assign n2632 = n2629 | n2630;
  assign n2633 = ~n2631 & n2632;
  assign n2634 = n3394 & n2633;
  assign n2635 = n3394 | n2633;
  assign n2636 = ~n2634 & n2635;
  assign n2637 = x29 & x47;
  assign n2638 = n2636 & n2637;
  assign n2639 = n2636 | n2637;
  assign n2640 = ~n2638 & n2639;
  assign n2641 = n3392 & n2640;
  assign n2642 = n3392 | n2640;
  assign n2643 = ~n2641 & n2642;
  assign n3405 = n2638 | n2640;
  assign n3406 = (n2638 & n3392) | (n2638 & n3405) | (n3392 & n3405);
  assign n2647 = x31 & x46;
  assign n4012 = n2647 & n4003;
  assign n4013 = n2647 & n3847;
  assign n4014 = (n3364 & n4012) | (n3364 & n4013) | (n4012 & n4013);
  assign n3861 = (n2626 & n2647) | (n2626 & n4014) | (n2647 & n4014);
  assign n4015 = (n2599 & n3861) | (n2599 & n4014) | (n3861 & n4014);
  assign n11992 = n2647 | n4014;
  assign n11993 = (n2626 & n4014) | (n2626 & n11992) | (n4014 & n11992);
  assign n4017 = (n2601 & n4015) | (n2601 & n11993) | (n4015 & n11993);
  assign n3863 = (n2599 & n4014) | (n2599 & n3861) | (n4014 & n3861);
  assign n3864 = (n3380 & n4017) | (n3380 & n3863) | (n4017 & n3863);
  assign n4018 = n2647 | n4003;
  assign n4019 = n2647 | n3847;
  assign n4020 = (n3364 & n4018) | (n3364 & n4019) | (n4018 & n4019);
  assign n3866 = n2626 | n4020;
  assign n4021 = (n2599 & n3866) | (n2599 & n4020) | (n3866 & n4020);
  assign n11994 = n2626 | n4020;
  assign n4023 = (n2601 & n4021) | (n2601 & n11994) | (n4021 & n11994);
  assign n3868 = (n2599 & n4020) | (n2599 & n3866) | (n4020 & n3866);
  assign n3869 = (n3380 & n4023) | (n3380 & n3868) | (n4023 & n3868);
  assign n2650 = ~n3864 & n3869;
  assign n3871 = n2631 & n2650;
  assign n4024 = (n2633 & n2650) | (n2633 & n3871) | (n2650 & n3871);
  assign n3872 = (n3394 & n4024) | (n3394 & n3871) | (n4024 & n3871);
  assign n3874 = n2631 | n2650;
  assign n4025 = n2633 | n3874;
  assign n3875 = (n3394 & n4025) | (n3394 & n3874) | (n4025 & n3874);
  assign n2653 = ~n3872 & n3875;
  assign n2654 = x30 & x47;
  assign n2655 = n2653 & n2654;
  assign n2656 = n2653 | n2654;
  assign n2657 = ~n2655 & n2656;
  assign n2658 = n3406 & n2657;
  assign n2659 = n3406 | n2657;
  assign n2660 = ~n2658 & n2659;
  assign n2663 = x31 & x47;
  assign n4026 = n2663 & n4017;
  assign n4027 = n2663 & n3863;
  assign n4028 = (n3380 & n4026) | (n3380 & n4027) | (n4026 & n4027);
  assign n3877 = (n2650 & n2663) | (n2650 & n4028) | (n2663 & n4028);
  assign n4029 = (n2631 & n3877) | (n2631 & n4028) | (n3877 & n4028);
  assign n11995 = n2663 | n4028;
  assign n11996 = (n2650 & n4028) | (n2650 & n11995) | (n4028 & n11995);
  assign n4031 = (n2633 & n4029) | (n2633 & n11996) | (n4029 & n11996);
  assign n3879 = (n2631 & n4028) | (n2631 & n3877) | (n4028 & n3877);
  assign n3880 = (n3394 & n4031) | (n3394 & n3879) | (n4031 & n3879);
  assign n4032 = n2663 | n4017;
  assign n4033 = n2663 | n3863;
  assign n4034 = (n3380 & n4032) | (n3380 & n4033) | (n4032 & n4033);
  assign n3882 = n2650 | n4034;
  assign n4035 = (n2631 & n3882) | (n2631 & n4034) | (n3882 & n4034);
  assign n11997 = n2650 | n4034;
  assign n4037 = (n2633 & n4035) | (n2633 & n11997) | (n4035 & n11997);
  assign n3884 = (n2631 & n4034) | (n2631 & n3882) | (n4034 & n3882);
  assign n3885 = (n3394 & n4037) | (n3394 & n3884) | (n4037 & n3884);
  assign n2666 = ~n3880 & n3885;
  assign n3887 = n2655 & n2666;
  assign n4038 = (n2657 & n2666) | (n2657 & n3887) | (n2666 & n3887);
  assign n3888 = (n3406 & n4038) | (n3406 & n3887) | (n4038 & n3887);
  assign n3890 = n2655 | n2666;
  assign n4039 = n2657 | n3890;
  assign n3891 = (n3406 & n4039) | (n3406 & n3890) | (n4039 & n3890);
  assign n2669 = ~n3888 & n3891;
  assign n3427 = n2666 | n3880;
  assign n3893 = (n2655 & n3427) | (n2655 & n3880) | (n3427 & n3880);
  assign n11998 = n2666 | n3880;
  assign n4041 = (n2657 & n3893) | (n2657 & n11998) | (n3893 & n11998);
  assign n3894 = (n3406 & n4041) | (n3406 & n3893) | (n4041 & n3893);
  assign n4106 = x48 & x80;
  assign n4107 = x49 & x80;
  assign n4108 = x48 & x81;
  assign n4109 = n4107 & n4108;
  assign n4110 = n4107 | n4108;
  assign n4111 = ~n4109 & n4110;
  assign n4112 = x50 & x80;
  assign n4113 = x49 & x81;
  assign n4114 = n4112 & n4113;
  assign n4115 = n4112 | n4113;
  assign n4116 = ~n4114 & n4115;
  assign n4117 = n4109 & n4116;
  assign n4118 = n4109 | n4116;
  assign n4119 = ~n4117 & n4118;
  assign n4120 = x48 & x82;
  assign n4121 = n4119 & n4120;
  assign n4122 = n4119 | n4120;
  assign n4123 = ~n4121 & n4122;
  assign n11999 = n4109 | n4114;
  assign n12000 = (n4114 & n4116) | (n4114 & n11999) | (n4116 & n11999);
  assign n4125 = x51 & x80;
  assign n4126 = x50 & x81;
  assign n4127 = n4125 & n4126;
  assign n4128 = n4125 | n4126;
  assign n4129 = ~n4127 & n4128;
  assign n4130 = n12000 & n4129;
  assign n4131 = n12000 | n4129;
  assign n4132 = ~n4130 & n4131;
  assign n4133 = x49 & x82;
  assign n4134 = n4132 & n4133;
  assign n4135 = n4132 | n4133;
  assign n4136 = ~n4134 & n4135;
  assign n4137 = n4121 & n4136;
  assign n4138 = n4121 | n4136;
  assign n4139 = ~n4137 & n4138;
  assign n4140 = x48 & x83;
  assign n4141 = n4139 & n4140;
  assign n4142 = n4139 | n4140;
  assign n4143 = ~n4141 & n4142;
  assign n12001 = n4121 | n4134;
  assign n12002 = (n4134 & n4136) | (n4134 & n12001) | (n4136 & n12001);
  assign n12003 = n4127 | n4129;
  assign n12004 = (n4127 & n12000) | (n4127 & n12003) | (n12000 & n12003);
  assign n4146 = x52 & x80;
  assign n4147 = x51 & x81;
  assign n4148 = n4146 & n4147;
  assign n4149 = n4146 | n4147;
  assign n4150 = ~n4148 & n4149;
  assign n4151 = n12004 & n4150;
  assign n4152 = n12004 | n4150;
  assign n4153 = ~n4151 & n4152;
  assign n4154 = x50 & x82;
  assign n4155 = n4153 & n4154;
  assign n4156 = n4153 | n4154;
  assign n4157 = ~n4155 & n4156;
  assign n4158 = n12002 & n4157;
  assign n4159 = n12002 | n4157;
  assign n4160 = ~n4158 & n4159;
  assign n4161 = x49 & x83;
  assign n4162 = n4160 & n4161;
  assign n4163 = n4160 | n4161;
  assign n4164 = ~n4162 & n4163;
  assign n4165 = n4141 & n4164;
  assign n4166 = n4141 | n4164;
  assign n4167 = ~n4165 & n4166;
  assign n4168 = x48 & x84;
  assign n4169 = n4167 & n4168;
  assign n4170 = n4167 | n4168;
  assign n4171 = ~n4169 & n4170;
  assign n12005 = n4141 | n4162;
  assign n12006 = (n4162 & n4164) | (n4162 & n12005) | (n4164 & n12005);
  assign n4175 = x53 & x80;
  assign n4176 = x52 & x81;
  assign n4177 = n4175 & n4176;
  assign n4178 = n4175 | n4176;
  assign n4179 = ~n4177 & n4178;
  assign n12007 = n4148 | n4150;
  assign n12009 = n4179 & n12007;
  assign n12010 = n4148 & n4179;
  assign n12011 = (n12004 & n12009) | (n12004 & n12010) | (n12009 & n12010);
  assign n12012 = n4179 | n12007;
  assign n12013 = n4148 | n4179;
  assign n12014 = (n12004 & n12012) | (n12004 & n12013) | (n12012 & n12013);
  assign n4182 = ~n12011 & n12014;
  assign n4183 = x51 & x82;
  assign n4184 = n4182 & n4183;
  assign n4185 = n4182 | n4183;
  assign n4186 = ~n4184 & n4185;
  assign n12015 = n4155 & n4186;
  assign n12016 = (n4158 & n4186) | (n4158 & n12015) | (n4186 & n12015);
  assign n12017 = n4155 | n4186;
  assign n12018 = n4158 | n12017;
  assign n4189 = ~n12016 & n12018;
  assign n4190 = x50 & x83;
  assign n4191 = n4189 & n4190;
  assign n4192 = n4189 | n4190;
  assign n4193 = ~n4191 & n4192;
  assign n4194 = n12006 & n4193;
  assign n4195 = n12006 | n4193;
  assign n4196 = ~n4194 & n4195;
  assign n4197 = x49 & x84;
  assign n4198 = n4196 & n4197;
  assign n4199 = n4196 | n4197;
  assign n4200 = ~n4198 & n4199;
  assign n4201 = n4169 & n4200;
  assign n4202 = n4169 | n4200;
  assign n4203 = ~n4201 & n4202;
  assign n4204 = x48 & x85;
  assign n4205 = n4203 & n4204;
  assign n4206 = n4203 | n4204;
  assign n4207 = ~n4205 & n4206;
  assign n12019 = n4169 | n4198;
  assign n12020 = (n4198 & n4200) | (n4198 & n12019) | (n4200 & n12019);
  assign n4209 = n4191 | n4194;
  assign n4212 = x54 & x80;
  assign n4213 = x53 & x81;
  assign n4214 = n4212 & n4213;
  assign n4215 = n4212 | n4213;
  assign n4216 = ~n4214 & n4215;
  assign n12021 = n4177 & n4216;
  assign n12022 = (n4216 & n12011) | (n4216 & n12021) | (n12011 & n12021);
  assign n12023 = n4177 | n4216;
  assign n12024 = n12011 | n12023;
  assign n4219 = ~n12022 & n12024;
  assign n4220 = x52 & x82;
  assign n4221 = n4219 & n4220;
  assign n4222 = n4219 | n4220;
  assign n4223 = ~n4221 & n4222;
  assign n12025 = n4184 & n4223;
  assign n12026 = (n4223 & n12016) | (n4223 & n12025) | (n12016 & n12025);
  assign n12027 = n4184 | n4223;
  assign n12028 = n12016 | n12027;
  assign n4226 = ~n12026 & n12028;
  assign n4227 = x51 & x83;
  assign n4228 = n4226 & n4227;
  assign n4229 = n4226 | n4227;
  assign n4230 = ~n4228 & n4229;
  assign n4231 = n4209 & n4230;
  assign n4232 = n4209 | n4230;
  assign n4233 = ~n4231 & n4232;
  assign n4234 = x50 & x84;
  assign n4235 = n4233 & n4234;
  assign n4236 = n4233 | n4234;
  assign n4237 = ~n4235 & n4236;
  assign n4238 = n12020 & n4237;
  assign n4239 = n12020 | n4237;
  assign n4240 = ~n4238 & n4239;
  assign n4241 = x49 & x85;
  assign n4242 = n4240 & n4241;
  assign n4243 = n4240 | n4241;
  assign n4244 = ~n4242 & n4243;
  assign n4245 = n4205 & n4244;
  assign n4246 = n4205 | n4244;
  assign n4247 = ~n4245 & n4246;
  assign n4248 = x48 & x86;
  assign n4249 = n4247 & n4248;
  assign n4250 = n4247 | n4248;
  assign n4251 = ~n4249 & n4250;
  assign n17674 = n4204 | n4241;
  assign n17675 = (n4203 & n4241) | (n4203 & n17674) | (n4241 & n17674);
  assign n15611 = (n4205 & n4240) | (n4205 & n17675) | (n4240 & n17675);
  assign n12030 = (n4242 & n4244) | (n4242 & n15611) | (n4244 & n15611);
  assign n12031 = n4235 | n12020;
  assign n12032 = (n4235 & n4237) | (n4235 & n12031) | (n4237 & n12031);
  assign n12033 = n4228 | n4230;
  assign n12034 = (n4209 & n4228) | (n4209 & n12033) | (n4228 & n12033);
  assign n4257 = x55 & x80;
  assign n4258 = x54 & x81;
  assign n4259 = n4257 & n4258;
  assign n4260 = n4257 | n4258;
  assign n4261 = ~n4259 & n4260;
  assign n15612 = n4177 | n4214;
  assign n15613 = (n4214 & n4216) | (n4214 & n15612) | (n4216 & n15612);
  assign n12038 = n4261 & n15613;
  assign n12036 = n4214 | n4216;
  assign n12039 = n4261 & n12036;
  assign n12040 = (n12011 & n12038) | (n12011 & n12039) | (n12038 & n12039);
  assign n12041 = n4261 | n15613;
  assign n12042 = n4261 | n12036;
  assign n12043 = (n12011 & n12041) | (n12011 & n12042) | (n12041 & n12042);
  assign n4264 = ~n12040 & n12043;
  assign n4265 = x53 & x82;
  assign n4266 = n4264 & n4265;
  assign n4267 = n4264 | n4265;
  assign n4268 = ~n4266 & n4267;
  assign n12044 = n4221 & n4268;
  assign n12045 = (n4268 & n12026) | (n4268 & n12044) | (n12026 & n12044);
  assign n12046 = n4221 | n4268;
  assign n12047 = n12026 | n12046;
  assign n4271 = ~n12045 & n12047;
  assign n4272 = x52 & x83;
  assign n4273 = n4271 & n4272;
  assign n4274 = n4271 | n4272;
  assign n4275 = ~n4273 & n4274;
  assign n4276 = n12034 & n4275;
  assign n4277 = n12034 | n4275;
  assign n4278 = ~n4276 & n4277;
  assign n4279 = x51 & x84;
  assign n4280 = n4278 & n4279;
  assign n4281 = n4278 | n4279;
  assign n4282 = ~n4280 & n4281;
  assign n4283 = n12032 & n4282;
  assign n4284 = n12032 | n4282;
  assign n4285 = ~n4283 & n4284;
  assign n4286 = x50 & x85;
  assign n4287 = n4285 & n4286;
  assign n4288 = n4285 | n4286;
  assign n4289 = ~n4287 & n4288;
  assign n4290 = n12030 & n4289;
  assign n4291 = n12030 | n4289;
  assign n4292 = ~n4290 & n4291;
  assign n4293 = x49 & x86;
  assign n4294 = n4292 & n4293;
  assign n4295 = n4292 | n4293;
  assign n4296 = ~n4294 & n4295;
  assign n4297 = n4249 & n4296;
  assign n4298 = n4249 | n4296;
  assign n4299 = ~n4297 & n4298;
  assign n4300 = x48 & x87;
  assign n4301 = n4299 & n4300;
  assign n4302 = n4299 | n4300;
  assign n4303 = ~n4301 & n4302;
  assign n12048 = n4249 | n4294;
  assign n12049 = (n4294 & n4296) | (n4294 & n12048) | (n4296 & n12048);
  assign n4305 = n4287 | n4290;
  assign n4306 = n4280 | n4283;
  assign n12050 = n4273 | n4275;
  assign n12051 = (n4273 & n12034) | (n4273 & n12050) | (n12034 & n12050);
  assign n4310 = x56 & x80;
  assign n4311 = x55 & x81;
  assign n4312 = n4310 & n4311;
  assign n4313 = n4310 | n4311;
  assign n4314 = ~n4312 & n4313;
  assign n12055 = n4259 & n4314;
  assign n15616 = (n4314 & n12039) | (n4314 & n12055) | (n12039 & n12055);
  assign n15617 = (n4314 & n12038) | (n4314 & n12055) | (n12038 & n12055);
  assign n15618 = (n12011 & n15616) | (n12011 & n15617) | (n15616 & n15617);
  assign n12057 = n4259 | n4314;
  assign n15619 = n12039 | n12057;
  assign n15620 = n12038 | n12057;
  assign n15621 = (n12011 & n15619) | (n12011 & n15620) | (n15619 & n15620);
  assign n4317 = ~n15618 & n15621;
  assign n4318 = x54 & x82;
  assign n4319 = n4317 & n4318;
  assign n4320 = n4317 | n4318;
  assign n4321 = ~n4319 & n4320;
  assign n12053 = n4266 | n4268;
  assign n15622 = n4321 & n12053;
  assign n15614 = n4221 | n4266;
  assign n15615 = (n4266 & n4268) | (n4266 & n15614) | (n4268 & n15614);
  assign n15623 = n4321 & n15615;
  assign n15624 = (n12026 & n15622) | (n12026 & n15623) | (n15622 & n15623);
  assign n15625 = n4321 | n12053;
  assign n15626 = n4321 | n15615;
  assign n15627 = (n12026 & n15625) | (n12026 & n15626) | (n15625 & n15626);
  assign n4324 = ~n15624 & n15627;
  assign n4325 = x53 & x83;
  assign n4326 = n4324 & n4325;
  assign n4327 = n4324 | n4325;
  assign n4328 = ~n4326 & n4327;
  assign n4329 = n12051 & n4328;
  assign n4330 = n12051 | n4328;
  assign n4331 = ~n4329 & n4330;
  assign n4332 = x52 & x84;
  assign n4333 = n4331 & n4332;
  assign n4334 = n4331 | n4332;
  assign n4335 = ~n4333 & n4334;
  assign n4336 = n4306 & n4335;
  assign n4337 = n4306 | n4335;
  assign n4338 = ~n4336 & n4337;
  assign n4339 = x51 & x85;
  assign n4340 = n4338 & n4339;
  assign n4341 = n4338 | n4339;
  assign n4342 = ~n4340 & n4341;
  assign n4343 = n4305 & n4342;
  assign n4344 = n4305 | n4342;
  assign n4345 = ~n4343 & n4344;
  assign n4346 = x50 & x86;
  assign n4347 = n4345 & n4346;
  assign n4348 = n4345 | n4346;
  assign n4349 = ~n4347 & n4348;
  assign n4350 = n12049 & n4349;
  assign n4351 = n12049 | n4349;
  assign n4352 = ~n4350 & n4351;
  assign n4353 = x49 & x87;
  assign n4354 = n4352 & n4353;
  assign n4355 = n4352 | n4353;
  assign n4356 = ~n4354 & n4355;
  assign n4357 = n4301 & n4356;
  assign n4358 = n4301 | n4356;
  assign n4359 = ~n4357 & n4358;
  assign n4360 = x48 & x88;
  assign n4361 = n4359 & n4360;
  assign n4362 = n4359 | n4360;
  assign n4363 = ~n4361 & n4362;
  assign n17676 = n4300 | n4353;
  assign n17677 = (n4299 & n4353) | (n4299 & n17676) | (n4353 & n17676);
  assign n15629 = (n4301 & n4352) | (n4301 & n17677) | (n4352 & n17677);
  assign n12060 = (n4354 & n4356) | (n4354 & n15629) | (n4356 & n15629);
  assign n12061 = n4347 | n12049;
  assign n12062 = (n4347 & n4349) | (n4347 & n12061) | (n4349 & n12061);
  assign n4366 = n4340 | n4343;
  assign n12063 = n4333 | n4335;
  assign n12064 = (n4306 & n4333) | (n4306 & n12063) | (n4333 & n12063);
  assign n12054 = (n12026 & n15615) | (n12026 & n12053) | (n15615 & n12053);
  assign n4371 = x57 & x80;
  assign n4372 = x56 & x81;
  assign n4373 = n4371 & n4372;
  assign n4374 = n4371 | n4372;
  assign n4375 = ~n4373 & n4374;
  assign n15630 = n4259 | n4312;
  assign n15631 = (n4312 & n4314) | (n4312 & n15630) | (n4314 & n15630);
  assign n12072 = n4375 & n15631;
  assign n12070 = n4312 | n4314;
  assign n12073 = n4375 & n12070;
  assign n15632 = (n12039 & n12072) | (n12039 & n12073) | (n12072 & n12073);
  assign n15633 = (n12038 & n12072) | (n12038 & n12073) | (n12072 & n12073);
  assign n15634 = (n12011 & n15632) | (n12011 & n15633) | (n15632 & n15633);
  assign n12075 = n4375 | n15631;
  assign n12076 = n4375 | n12070;
  assign n15635 = (n12039 & n12075) | (n12039 & n12076) | (n12075 & n12076);
  assign n15636 = (n12038 & n12075) | (n12038 & n12076) | (n12075 & n12076);
  assign n15637 = (n12011 & n15635) | (n12011 & n15636) | (n15635 & n15636);
  assign n4378 = ~n15634 & n15637;
  assign n4379 = x55 & x82;
  assign n4380 = n4378 & n4379;
  assign n4381 = n4378 | n4379;
  assign n4382 = ~n4380 & n4381;
  assign n12067 = n4319 | n4321;
  assign n12078 = n4382 & n12067;
  assign n12079 = n4319 & n4382;
  assign n12080 = (n12054 & n12078) | (n12054 & n12079) | (n12078 & n12079);
  assign n12081 = n4382 | n12067;
  assign n12082 = n4319 | n4382;
  assign n12083 = (n12054 & n12081) | (n12054 & n12082) | (n12081 & n12082);
  assign n4385 = ~n12080 & n12083;
  assign n4386 = x54 & x83;
  assign n4387 = n4385 & n4386;
  assign n4388 = n4385 | n4386;
  assign n4389 = ~n4387 & n4388;
  assign n12065 = n4326 | n4328;
  assign n15638 = n4389 & n12065;
  assign n15639 = n4326 & n4389;
  assign n15640 = (n12051 & n15638) | (n12051 & n15639) | (n15638 & n15639);
  assign n15641 = n4389 | n12065;
  assign n15642 = n4326 | n4389;
  assign n15643 = (n12051 & n15641) | (n12051 & n15642) | (n15641 & n15642);
  assign n4392 = ~n15640 & n15643;
  assign n4393 = x53 & x84;
  assign n4394 = n4392 & n4393;
  assign n4395 = n4392 | n4393;
  assign n4396 = ~n4394 & n4395;
  assign n4397 = n12064 & n4396;
  assign n4398 = n12064 | n4396;
  assign n4399 = ~n4397 & n4398;
  assign n4400 = x52 & x85;
  assign n4401 = n4399 & n4400;
  assign n4402 = n4399 | n4400;
  assign n4403 = ~n4401 & n4402;
  assign n4404 = n4366 & n4403;
  assign n4405 = n4366 | n4403;
  assign n4406 = ~n4404 & n4405;
  assign n4407 = x51 & x86;
  assign n4408 = n4406 & n4407;
  assign n4409 = n4406 | n4407;
  assign n4410 = ~n4408 & n4409;
  assign n4411 = n12062 & n4410;
  assign n4412 = n12062 | n4410;
  assign n4413 = ~n4411 & n4412;
  assign n4414 = x50 & x87;
  assign n4415 = n4413 & n4414;
  assign n4416 = n4413 | n4414;
  assign n4417 = ~n4415 & n4416;
  assign n4418 = n12060 & n4417;
  assign n4419 = n12060 | n4417;
  assign n4420 = ~n4418 & n4419;
  assign n4421 = x49 & x88;
  assign n4422 = n4420 & n4421;
  assign n4423 = n4420 | n4421;
  assign n4424 = ~n4422 & n4423;
  assign n4425 = n4361 & n4424;
  assign n4426 = n4361 | n4424;
  assign n4427 = ~n4425 & n4426;
  assign n4428 = x48 & x89;
  assign n4429 = n4427 & n4428;
  assign n4430 = n4427 | n4428;
  assign n4431 = ~n4429 & n4430;
  assign n17678 = n4360 | n4421;
  assign n17679 = (n4359 & n4421) | (n4359 & n17678) | (n4421 & n17678);
  assign n15645 = (n4361 & n4420) | (n4361 & n17679) | (n4420 & n17679);
  assign n12085 = (n4422 & n4424) | (n4422 & n15645) | (n4424 & n15645);
  assign n12086 = n4415 | n12060;
  assign n12087 = (n4415 & n4417) | (n4415 & n12086) | (n4417 & n12086);
  assign n12088 = n4408 | n12062;
  assign n12089 = (n4408 & n4410) | (n4408 & n12088) | (n4410 & n12088);
  assign n12090 = n4401 | n4403;
  assign n12091 = (n4366 & n4401) | (n4366 & n12090) | (n4401 & n12090);
  assign n12066 = (n4326 & n12051) | (n4326 & n12065) | (n12051 & n12065);
  assign n15646 = n4373 | n4375;
  assign n15647 = (n4373 & n15631) | (n4373 & n15646) | (n15631 & n15646);
  assign n15648 = (n4373 & n12070) | (n4373 & n15646) | (n12070 & n15646);
  assign n15649 = (n12039 & n15647) | (n12039 & n15648) | (n15647 & n15648);
  assign n15650 = (n12038 & n15647) | (n12038 & n15648) | (n15647 & n15648);
  assign n15651 = (n12011 & n15649) | (n12011 & n15650) | (n15649 & n15650);
  assign n4440 = x58 & x80;
  assign n4441 = x57 & x81;
  assign n4442 = n4440 & n4441;
  assign n4443 = n4440 | n4441;
  assign n4444 = ~n4442 & n4443;
  assign n4445 = n15651 & n4444;
  assign n4446 = n15651 | n4444;
  assign n4447 = ~n4445 & n4446;
  assign n4448 = x56 & x82;
  assign n4449 = n4447 & n4448;
  assign n4450 = n4447 | n4448;
  assign n4451 = ~n4449 & n4450;
  assign n12099 = n4380 & n4451;
  assign n15652 = (n4451 & n12078) | (n4451 & n12099) | (n12078 & n12099);
  assign n15653 = (n4451 & n12079) | (n4451 & n12099) | (n12079 & n12099);
  assign n15654 = (n12054 & n15652) | (n12054 & n15653) | (n15652 & n15653);
  assign n12101 = n4380 | n4451;
  assign n15655 = n12078 | n12101;
  assign n15656 = n12079 | n12101;
  assign n15657 = (n12054 & n15655) | (n12054 & n15656) | (n15655 & n15656);
  assign n4454 = ~n15654 & n15657;
  assign n4455 = x55 & x83;
  assign n4456 = n4454 & n4455;
  assign n4457 = n4454 | n4455;
  assign n4458 = ~n4456 & n4457;
  assign n12094 = n4387 | n4389;
  assign n12103 = n4458 & n12094;
  assign n12104 = n4387 & n4458;
  assign n12105 = (n12066 & n12103) | (n12066 & n12104) | (n12103 & n12104);
  assign n12106 = n4458 | n12094;
  assign n12107 = n4387 | n4458;
  assign n12108 = (n12066 & n12106) | (n12066 & n12107) | (n12106 & n12107);
  assign n4461 = ~n12105 & n12108;
  assign n4462 = x54 & x84;
  assign n4463 = n4461 & n4462;
  assign n4464 = n4461 | n4462;
  assign n4465 = ~n4463 & n4464;
  assign n12092 = n4394 | n4396;
  assign n15658 = n4465 & n12092;
  assign n15659 = n4394 & n4465;
  assign n15660 = (n12064 & n15658) | (n12064 & n15659) | (n15658 & n15659);
  assign n15661 = n4465 | n12092;
  assign n15662 = n4394 | n4465;
  assign n15663 = (n12064 & n15661) | (n12064 & n15662) | (n15661 & n15662);
  assign n4468 = ~n15660 & n15663;
  assign n4469 = x53 & x85;
  assign n4470 = n4468 & n4469;
  assign n4471 = n4468 | n4469;
  assign n4472 = ~n4470 & n4471;
  assign n4473 = n12091 & n4472;
  assign n4474 = n12091 | n4472;
  assign n4475 = ~n4473 & n4474;
  assign n4476 = x52 & x86;
  assign n4477 = n4475 & n4476;
  assign n4478 = n4475 | n4476;
  assign n4479 = ~n4477 & n4478;
  assign n4480 = n12089 & n4479;
  assign n4481 = n12089 | n4479;
  assign n4482 = ~n4480 & n4481;
  assign n4483 = x51 & x87;
  assign n4484 = n4482 & n4483;
  assign n4485 = n4482 | n4483;
  assign n4486 = ~n4484 & n4485;
  assign n4487 = n12087 & n4486;
  assign n4488 = n12087 | n4486;
  assign n4489 = ~n4487 & n4488;
  assign n4490 = x50 & x88;
  assign n4491 = n4489 & n4490;
  assign n4492 = n4489 | n4490;
  assign n4493 = ~n4491 & n4492;
  assign n4494 = n12085 & n4493;
  assign n4495 = n12085 | n4493;
  assign n4496 = ~n4494 & n4495;
  assign n4497 = x49 & x89;
  assign n4498 = n4496 & n4497;
  assign n4499 = n4496 | n4497;
  assign n4500 = ~n4498 & n4499;
  assign n4501 = n4429 & n4500;
  assign n4502 = n4429 | n4500;
  assign n4503 = ~n4501 & n4502;
  assign n4504 = x48 & x90;
  assign n4505 = n4503 & n4504;
  assign n4506 = n4503 | n4504;
  assign n4507 = ~n4505 & n4506;
  assign n12109 = n4429 | n4498;
  assign n12110 = (n4498 & n4500) | (n4498 & n12109) | (n4500 & n12109);
  assign n4509 = n4491 | n4494;
  assign n4510 = n4484 | n4487;
  assign n12093 = (n4394 & n12064) | (n4394 & n12092) | (n12064 & n12092);
  assign n12116 = n4449 | n4451;
  assign n15664 = n4380 | n4449;
  assign n15665 = (n4449 & n4451) | (n4449 & n15664) | (n4451 & n15664);
  assign n15666 = (n12078 & n12116) | (n12078 & n15665) | (n12116 & n15665);
  assign n15667 = (n12079 & n12116) | (n12079 & n15665) | (n12116 & n15665);
  assign n15668 = (n12054 & n15666) | (n12054 & n15667) | (n15666 & n15667);
  assign n4517 = x59 & x80;
  assign n4518 = x58 & x81;
  assign n4519 = n4517 & n4518;
  assign n4520 = n4517 | n4518;
  assign n4521 = ~n4519 & n4520;
  assign n12118 = n4442 | n4444;
  assign n12120 = n4521 & n12118;
  assign n12121 = n4442 & n4521;
  assign n12122 = (n15651 & n12120) | (n15651 & n12121) | (n12120 & n12121);
  assign n12123 = n4521 | n12118;
  assign n12124 = n4442 | n4521;
  assign n12125 = (n15651 & n12123) | (n15651 & n12124) | (n12123 & n12124);
  assign n4524 = ~n12122 & n12125;
  assign n4525 = x57 & x82;
  assign n4526 = n4524 & n4525;
  assign n4527 = n4524 | n4525;
  assign n4528 = ~n4526 & n4527;
  assign n4529 = n15668 & n4528;
  assign n4530 = n15668 | n4528;
  assign n4531 = ~n4529 & n4530;
  assign n4532 = x56 & x83;
  assign n4533 = n4531 & n4532;
  assign n4534 = n4531 | n4532;
  assign n4535 = ~n4533 & n4534;
  assign n12126 = n4456 & n4535;
  assign n12127 = (n4535 & n12105) | (n4535 & n12126) | (n12105 & n12126);
  assign n12128 = n4456 | n4535;
  assign n12129 = n12105 | n12128;
  assign n4538 = ~n12127 & n12129;
  assign n4539 = x55 & x84;
  assign n4540 = n4538 & n4539;
  assign n4541 = n4538 | n4539;
  assign n4542 = ~n4540 & n4541;
  assign n12113 = n4463 | n4465;
  assign n12130 = n4542 & n12113;
  assign n12131 = n4463 & n4542;
  assign n12132 = (n12093 & n12130) | (n12093 & n12131) | (n12130 & n12131);
  assign n12133 = n4542 | n12113;
  assign n12134 = n4463 | n4542;
  assign n12135 = (n12093 & n12133) | (n12093 & n12134) | (n12133 & n12134);
  assign n4545 = ~n12132 & n12135;
  assign n4546 = x54 & x85;
  assign n4547 = n4545 & n4546;
  assign n4548 = n4545 | n4546;
  assign n4549 = ~n4547 & n4548;
  assign n12111 = n4470 | n4472;
  assign n15669 = n4549 & n12111;
  assign n15670 = n4470 & n4549;
  assign n15671 = (n12091 & n15669) | (n12091 & n15670) | (n15669 & n15670);
  assign n15672 = n4549 | n12111;
  assign n15673 = n4470 | n4549;
  assign n15674 = (n12091 & n15672) | (n12091 & n15673) | (n15672 & n15673);
  assign n4552 = ~n15671 & n15674;
  assign n4553 = x53 & x86;
  assign n4554 = n4552 & n4553;
  assign n4555 = n4552 | n4553;
  assign n4556 = ~n4554 & n4555;
  assign n15675 = n4477 & n4556;
  assign n15676 = (n4480 & n4556) | (n4480 & n15675) | (n4556 & n15675);
  assign n15677 = n4477 | n4556;
  assign n15678 = n4480 | n15677;
  assign n4559 = ~n15676 & n15678;
  assign n4560 = x52 & x87;
  assign n4561 = n4559 & n4560;
  assign n4562 = n4559 | n4560;
  assign n4563 = ~n4561 & n4562;
  assign n4564 = n4510 & n4563;
  assign n4565 = n4510 | n4563;
  assign n4566 = ~n4564 & n4565;
  assign n4567 = x51 & x88;
  assign n4568 = n4566 & n4567;
  assign n4569 = n4566 | n4567;
  assign n4570 = ~n4568 & n4569;
  assign n4571 = n4509 & n4570;
  assign n4572 = n4509 | n4570;
  assign n4573 = ~n4571 & n4572;
  assign n4574 = x50 & x89;
  assign n4575 = n4573 & n4574;
  assign n4576 = n4573 | n4574;
  assign n4577 = ~n4575 & n4576;
  assign n4578 = n12110 & n4577;
  assign n4579 = n12110 | n4577;
  assign n4580 = ~n4578 & n4579;
  assign n4581 = x49 & x90;
  assign n4582 = n4580 & n4581;
  assign n4583 = n4580 | n4581;
  assign n4584 = ~n4582 & n4583;
  assign n4585 = n4505 & n4584;
  assign n4586 = n4505 | n4584;
  assign n4587 = ~n4585 & n4586;
  assign n4588 = x48 & x91;
  assign n4589 = n4587 & n4588;
  assign n4590 = n4587 | n4588;
  assign n4591 = ~n4589 & n4590;
  assign n17680 = n4504 | n4581;
  assign n17681 = (n4503 & n4581) | (n4503 & n17680) | (n4581 & n17680);
  assign n15680 = (n4505 & n4580) | (n4505 & n17681) | (n4580 & n17681);
  assign n12137 = (n4582 & n4584) | (n4582 & n15680) | (n4584 & n15680);
  assign n12138 = n4575 | n12110;
  assign n12139 = (n4575 & n4577) | (n4575 & n12138) | (n4577 & n12138);
  assign n4594 = n4568 | n4571;
  assign n15681 = n4561 | n4563;
  assign n15682 = (n4510 & n4561) | (n4510 & n15681) | (n4561 & n15681);
  assign n4511 = n4477 | n4480;
  assign n12112 = (n4470 & n12091) | (n4470 & n12111) | (n12091 & n12111);
  assign n4602 = x60 & x80;
  assign n4603 = x59 & x81;
  assign n4604 = n4602 & n4603;
  assign n4605 = n4602 | n4603;
  assign n4606 = ~n4604 & n4605;
  assign n15683 = n4519 | n4521;
  assign n15684 = (n4519 & n12118) | (n4519 & n15683) | (n12118 & n15683);
  assign n12149 = n4606 & n15684;
  assign n15685 = n4442 | n4519;
  assign n15686 = (n4519 & n4521) | (n4519 & n15685) | (n4521 & n15685);
  assign n12150 = n4606 & n15686;
  assign n12151 = (n15651 & n12149) | (n15651 & n12150) | (n12149 & n12150);
  assign n12152 = n4606 | n15684;
  assign n12153 = n4606 | n15686;
  assign n12154 = (n15651 & n12152) | (n15651 & n12153) | (n12152 & n12153);
  assign n4609 = ~n12151 & n12154;
  assign n4610 = x58 & x82;
  assign n4611 = n4609 & n4610;
  assign n4612 = n4609 | n4610;
  assign n4613 = ~n4611 & n4612;
  assign n12144 = n4526 | n4528;
  assign n12155 = n4613 & n12144;
  assign n12156 = n4526 & n4613;
  assign n12157 = (n15668 & n12155) | (n15668 & n12156) | (n12155 & n12156);
  assign n12158 = n4613 | n12144;
  assign n12159 = n4526 | n4613;
  assign n12160 = (n15668 & n12158) | (n15668 & n12159) | (n12158 & n12159);
  assign n4616 = ~n12157 & n12160;
  assign n4617 = x57 & x83;
  assign n4618 = n4616 & n4617;
  assign n4619 = n4616 | n4617;
  assign n4620 = ~n4618 & n4619;
  assign n12161 = n4533 & n4620;
  assign n15687 = (n4620 & n12126) | (n4620 & n12161) | (n12126 & n12161);
  assign n15688 = (n4535 & n4620) | (n4535 & n12161) | (n4620 & n12161);
  assign n15689 = (n12105 & n15687) | (n12105 & n15688) | (n15687 & n15688);
  assign n12163 = n4533 | n4620;
  assign n15690 = n12126 | n12163;
  assign n15691 = n4535 | n12163;
  assign n15692 = (n12105 & n15690) | (n12105 & n15691) | (n15690 & n15691);
  assign n4623 = ~n15689 & n15692;
  assign n4624 = x56 & x84;
  assign n4625 = n4623 & n4624;
  assign n4626 = n4623 | n4624;
  assign n4627 = ~n4625 & n4626;
  assign n12165 = n4540 & n4627;
  assign n12166 = (n4627 & n12132) | (n4627 & n12165) | (n12132 & n12165);
  assign n12167 = n4540 | n4627;
  assign n12168 = n12132 | n12167;
  assign n4630 = ~n12166 & n12168;
  assign n4631 = x55 & x85;
  assign n4632 = n4630 & n4631;
  assign n4633 = n4630 | n4631;
  assign n4634 = ~n4632 & n4633;
  assign n12142 = n4547 | n4549;
  assign n12169 = n4634 & n12142;
  assign n12170 = n4547 & n4634;
  assign n12171 = (n12112 & n12169) | (n12112 & n12170) | (n12169 & n12170);
  assign n12172 = n4634 | n12142;
  assign n12173 = n4547 | n4634;
  assign n12174 = (n12112 & n12172) | (n12112 & n12173) | (n12172 & n12173);
  assign n4637 = ~n12171 & n12174;
  assign n4638 = x54 & x86;
  assign n4639 = n4637 & n4638;
  assign n4640 = n4637 | n4638;
  assign n4641 = ~n4639 & n4640;
  assign n12140 = n4554 | n4556;
  assign n15693 = n4641 & n12140;
  assign n15694 = n4554 & n4641;
  assign n15695 = (n4511 & n15693) | (n4511 & n15694) | (n15693 & n15694);
  assign n15696 = n4641 | n12140;
  assign n15697 = n4554 | n4641;
  assign n15698 = (n4511 & n15696) | (n4511 & n15697) | (n15696 & n15697);
  assign n4644 = ~n15695 & n15698;
  assign n4645 = x53 & x87;
  assign n4646 = n4644 & n4645;
  assign n4647 = n4644 | n4645;
  assign n4648 = ~n4646 & n4647;
  assign n4649 = n15682 & n4648;
  assign n4650 = n15682 | n4648;
  assign n4651 = ~n4649 & n4650;
  assign n4652 = x52 & x88;
  assign n4653 = n4651 & n4652;
  assign n4654 = n4651 | n4652;
  assign n4655 = ~n4653 & n4654;
  assign n4656 = n4594 & n4655;
  assign n4657 = n4594 | n4655;
  assign n4658 = ~n4656 & n4657;
  assign n4659 = x51 & x89;
  assign n4660 = n4658 & n4659;
  assign n4661 = n4658 | n4659;
  assign n4662 = ~n4660 & n4661;
  assign n4663 = n12139 & n4662;
  assign n4664 = n12139 | n4662;
  assign n4665 = ~n4663 & n4664;
  assign n4666 = x50 & x90;
  assign n4667 = n4665 & n4666;
  assign n4668 = n4665 | n4666;
  assign n4669 = ~n4667 & n4668;
  assign n4670 = n12137 & n4669;
  assign n4671 = n12137 | n4669;
  assign n4672 = ~n4670 & n4671;
  assign n4673 = x49 & x91;
  assign n4674 = n4672 & n4673;
  assign n4675 = n4672 | n4673;
  assign n4676 = ~n4674 & n4675;
  assign n4677 = n4589 & n4676;
  assign n4678 = n4589 | n4676;
  assign n4679 = ~n4677 & n4678;
  assign n4680 = x48 & x92;
  assign n4681 = n4679 & n4680;
  assign n4682 = n4679 | n4680;
  assign n4683 = ~n4681 & n4682;
  assign n17682 = n4588 | n4673;
  assign n17683 = (n4587 & n4673) | (n4587 & n17682) | (n4673 & n17682);
  assign n15700 = (n4589 & n4672) | (n4589 & n17683) | (n4672 & n17683);
  assign n12176 = (n4674 & n4676) | (n4674 & n15700) | (n4676 & n15700);
  assign n12177 = n4667 | n12137;
  assign n12178 = (n4667 & n4669) | (n4667 & n12177) | (n4669 & n12177);
  assign n12179 = n4660 | n12139;
  assign n12180 = (n4660 & n4662) | (n4660 & n12179) | (n4662 & n12179);
  assign n15701 = n4653 | n4655;
  assign n15702 = (n4594 & n4653) | (n4594 & n15701) | (n4653 & n15701);
  assign n12181 = n4646 | n4648;
  assign n12182 = (n15682 & n4646) | (n15682 & n12181) | (n4646 & n12181);
  assign n12141 = (n4511 & n4554) | (n4511 & n12140) | (n4554 & n12140);
  assign n12186 = n4618 | n4620;
  assign n15703 = n4533 | n4618;
  assign n15704 = (n4618 & n4620) | (n4618 & n15703) | (n4620 & n15703);
  assign n15705 = (n12126 & n12186) | (n12126 & n15704) | (n12186 & n15704);
  assign n15706 = (n4535 & n12186) | (n4535 & n15704) | (n12186 & n15704);
  assign n15707 = (n12105 & n15705) | (n12105 & n15706) | (n15705 & n15706);
  assign n4695 = x61 & x80;
  assign n4696 = x60 & x81;
  assign n4697 = n4695 & n4696;
  assign n4698 = n4695 | n4696;
  assign n4699 = ~n4697 & n4698;
  assign n15712 = n4604 | n4606;
  assign n17684 = n4699 & n15712;
  assign n17685 = n4604 & n4699;
  assign n17686 = (n15684 & n17684) | (n15684 & n17685) | (n17684 & n17685);
  assign n15714 = (n4604 & n15686) | (n4604 & n15712) | (n15686 & n15712);
  assign n15716 = n4699 & n15714;
  assign n15717 = (n15651 & n17686) | (n15651 & n15716) | (n17686 & n15716);
  assign n17687 = n4699 | n15712;
  assign n17688 = n4604 | n4699;
  assign n17689 = (n15684 & n17687) | (n15684 & n17688) | (n17687 & n17688);
  assign n15719 = n4699 | n15714;
  assign n15720 = (n15651 & n17689) | (n15651 & n15719) | (n17689 & n15719);
  assign n4702 = ~n15717 & n15720;
  assign n4703 = x59 & x82;
  assign n4704 = n4702 & n4703;
  assign n4705 = n4702 | n4703;
  assign n4706 = ~n4704 & n4705;
  assign n15708 = n4611 | n4613;
  assign n15709 = (n4611 & n12144) | (n4611 & n15708) | (n12144 & n15708);
  assign n15721 = n4706 & n15709;
  assign n15710 = n4526 | n4611;
  assign n15711 = (n4611 & n4613) | (n4611 & n15710) | (n4613 & n15710);
  assign n15722 = n4706 & n15711;
  assign n15723 = (n15668 & n15721) | (n15668 & n15722) | (n15721 & n15722);
  assign n15724 = n4706 | n15709;
  assign n15725 = n4706 | n15711;
  assign n15726 = (n15668 & n15724) | (n15668 & n15725) | (n15724 & n15725);
  assign n4709 = ~n15723 & n15726;
  assign n4710 = x58 & x83;
  assign n4711 = n4709 & n4710;
  assign n4712 = n4709 | n4710;
  assign n4713 = ~n4711 & n4712;
  assign n4714 = n15707 & n4713;
  assign n4715 = n15707 | n4713;
  assign n4716 = ~n4714 & n4715;
  assign n4717 = x57 & x84;
  assign n4718 = n4716 & n4717;
  assign n4719 = n4716 | n4717;
  assign n4720 = ~n4718 & n4719;
  assign n12194 = n4625 & n4720;
  assign n12195 = (n4720 & n12166) | (n4720 & n12194) | (n12166 & n12194);
  assign n12196 = n4625 | n4720;
  assign n12197 = n12166 | n12196;
  assign n4723 = ~n12195 & n12197;
  assign n4724 = x56 & x85;
  assign n4725 = n4723 & n4724;
  assign n4726 = n4723 | n4724;
  assign n4727 = ~n4725 & n4726;
  assign n12198 = n4632 & n4727;
  assign n12199 = (n4727 & n12171) | (n4727 & n12198) | (n12171 & n12198);
  assign n12200 = n4632 | n4727;
  assign n12201 = n12171 | n12200;
  assign n4730 = ~n12199 & n12201;
  assign n4731 = x55 & x86;
  assign n4732 = n4730 & n4731;
  assign n4733 = n4730 | n4731;
  assign n4734 = ~n4732 & n4733;
  assign n12183 = n4639 | n4641;
  assign n12202 = n4734 & n12183;
  assign n12203 = n4639 & n4734;
  assign n12204 = (n12141 & n12202) | (n12141 & n12203) | (n12202 & n12203);
  assign n12205 = n4734 | n12183;
  assign n12206 = n4639 | n4734;
  assign n12207 = (n12141 & n12205) | (n12141 & n12206) | (n12205 & n12206);
  assign n4737 = ~n12204 & n12207;
  assign n4738 = x54 & x87;
  assign n4739 = n4737 & n4738;
  assign n4740 = n4737 | n4738;
  assign n4741 = ~n4739 & n4740;
  assign n4742 = n12182 & n4741;
  assign n4743 = n12182 | n4741;
  assign n4744 = ~n4742 & n4743;
  assign n4745 = x53 & x88;
  assign n4746 = n4744 & n4745;
  assign n4747 = n4744 | n4745;
  assign n4748 = ~n4746 & n4747;
  assign n4749 = n15702 & n4748;
  assign n4750 = n15702 | n4748;
  assign n4751 = ~n4749 & n4750;
  assign n4752 = x52 & x89;
  assign n4753 = n4751 & n4752;
  assign n4754 = n4751 | n4752;
  assign n4755 = ~n4753 & n4754;
  assign n4756 = n12180 & n4755;
  assign n4757 = n12180 | n4755;
  assign n4758 = ~n4756 & n4757;
  assign n4759 = x51 & x90;
  assign n4760 = n4758 & n4759;
  assign n4761 = n4758 | n4759;
  assign n4762 = ~n4760 & n4761;
  assign n4763 = n12178 & n4762;
  assign n4764 = n12178 | n4762;
  assign n4765 = ~n4763 & n4764;
  assign n4766 = x50 & x91;
  assign n4767 = n4765 & n4766;
  assign n4768 = n4765 | n4766;
  assign n4769 = ~n4767 & n4768;
  assign n4770 = n12176 & n4769;
  assign n4771 = n12176 | n4769;
  assign n4772 = ~n4770 & n4771;
  assign n4773 = x49 & x92;
  assign n4774 = n4772 & n4773;
  assign n4775 = n4772 | n4773;
  assign n4776 = ~n4774 & n4775;
  assign n4777 = n4681 & n4776;
  assign n4778 = n4681 | n4776;
  assign n4779 = ~n4777 & n4778;
  assign n4780 = x48 & x93;
  assign n4781 = n4779 & n4780;
  assign n4782 = n4779 | n4780;
  assign n4783 = ~n4781 & n4782;
  assign n12208 = n4681 | n4774;
  assign n12209 = (n4774 & n4776) | (n4774 & n12208) | (n4776 & n12208);
  assign n12210 = n4767 | n12176;
  assign n12211 = (n4767 & n4769) | (n4767 & n12210) | (n4769 & n12210);
  assign n12212 = n4760 | n12178;
  assign n12213 = (n4760 & n4762) | (n4760 & n12212) | (n4762 & n12212);
  assign n12214 = n4753 | n12180;
  assign n12215 = (n4753 & n4755) | (n4753 & n12214) | (n4755 & n12214);
  assign n12216 = n4746 | n4748;
  assign n12217 = (n15702 & n4746) | (n15702 & n12216) | (n4746 & n12216);
  assign n4796 = x62 & x80;
  assign n4797 = x61 & x81;
  assign n4798 = n4796 & n4797;
  assign n4799 = n4796 | n4797;
  assign n4800 = ~n4798 & n4799;
  assign n12224 = n4697 | n4699;
  assign n12226 = n4800 & n12224;
  assign n12227 = n4697 & n4800;
  assign n15713 = (n4604 & n15684) | (n4604 & n15712) | (n15684 & n15712);
  assign n15727 = (n12226 & n12227) | (n12226 & n15713) | (n12227 & n15713);
  assign n15728 = (n12226 & n12227) | (n12226 & n15714) | (n12227 & n15714);
  assign n15729 = (n15651 & n15727) | (n15651 & n15728) | (n15727 & n15728);
  assign n12229 = n4800 | n12224;
  assign n12230 = n4697 | n4800;
  assign n15730 = (n12229 & n12230) | (n12229 & n15713) | (n12230 & n15713);
  assign n15731 = (n12229 & n12230) | (n12229 & n15714) | (n12230 & n15714);
  assign n15732 = (n15651 & n15730) | (n15651 & n15731) | (n15730 & n15731);
  assign n4803 = ~n15729 & n15732;
  assign n4804 = x60 & x82;
  assign n4805 = n4803 & n4804;
  assign n4806 = n4803 | n4804;
  assign n4807 = ~n4805 & n4806;
  assign n12222 = n4704 | n4706;
  assign n12232 = n4807 & n12222;
  assign n12233 = n4704 & n4807;
  assign n15733 = (n12232 & n12233) | (n12232 & n15709) | (n12233 & n15709);
  assign n15734 = (n12232 & n12233) | (n12232 & n15711) | (n12233 & n15711);
  assign n15735 = (n15668 & n15733) | (n15668 & n15734) | (n15733 & n15734);
  assign n12235 = n4807 | n12222;
  assign n12236 = n4704 | n4807;
  assign n15736 = (n12235 & n12236) | (n12235 & n15709) | (n12236 & n15709);
  assign n15737 = (n12235 & n12236) | (n12235 & n15711) | (n12236 & n15711);
  assign n15738 = (n15668 & n15736) | (n15668 & n15737) | (n15736 & n15737);
  assign n4810 = ~n15735 & n15738;
  assign n4811 = x59 & x83;
  assign n4812 = n4810 & n4811;
  assign n4813 = n4810 | n4811;
  assign n4814 = ~n4812 & n4813;
  assign n12220 = n4711 | n4713;
  assign n12238 = n4814 & n12220;
  assign n12239 = n4711 & n4814;
  assign n12240 = (n15707 & n12238) | (n15707 & n12239) | (n12238 & n12239);
  assign n12241 = n4814 | n12220;
  assign n12242 = n4711 | n4814;
  assign n12243 = (n15707 & n12241) | (n15707 & n12242) | (n12241 & n12242);
  assign n4817 = ~n12240 & n12243;
  assign n4818 = x58 & x84;
  assign n4819 = n4817 & n4818;
  assign n4820 = n4817 | n4818;
  assign n4821 = ~n4819 & n4820;
  assign n12244 = n4718 & n4821;
  assign n15739 = (n4821 & n12194) | (n4821 & n12244) | (n12194 & n12244);
  assign n15740 = (n4720 & n4821) | (n4720 & n12244) | (n4821 & n12244);
  assign n15741 = (n12166 & n15739) | (n12166 & n15740) | (n15739 & n15740);
  assign n12246 = n4718 | n4821;
  assign n15742 = n12194 | n12246;
  assign n15743 = n4720 | n12246;
  assign n15744 = (n12166 & n15742) | (n12166 & n15743) | (n15742 & n15743);
  assign n4824 = ~n15741 & n15744;
  assign n4825 = x57 & x85;
  assign n4826 = n4824 & n4825;
  assign n4827 = n4824 | n4825;
  assign n4828 = ~n4826 & n4827;
  assign n12248 = n4725 & n4828;
  assign n12249 = (n4828 & n12199) | (n4828 & n12248) | (n12199 & n12248);
  assign n12250 = n4725 | n4828;
  assign n12251 = n12199 | n12250;
  assign n4831 = ~n12249 & n12251;
  assign n4832 = x56 & x86;
  assign n4833 = n4831 & n4832;
  assign n4834 = n4831 | n4832;
  assign n4835 = ~n4833 & n4834;
  assign n12252 = n4732 & n4835;
  assign n12253 = (n4835 & n12204) | (n4835 & n12252) | (n12204 & n12252);
  assign n12254 = n4732 | n4835;
  assign n12255 = n12204 | n12254;
  assign n4838 = ~n12253 & n12255;
  assign n4839 = x55 & x87;
  assign n4840 = n4838 & n4839;
  assign n4841 = n4838 | n4839;
  assign n4842 = ~n4840 & n4841;
  assign n12218 = n4739 | n4741;
  assign n12256 = n4842 & n12218;
  assign n12257 = n4739 & n4842;
  assign n12258 = (n12182 & n12256) | (n12182 & n12257) | (n12256 & n12257);
  assign n12259 = n4842 | n12218;
  assign n12260 = n4739 | n4842;
  assign n12261 = (n12182 & n12259) | (n12182 & n12260) | (n12259 & n12260);
  assign n4845 = ~n12258 & n12261;
  assign n4846 = x54 & x88;
  assign n4847 = n4845 & n4846;
  assign n4848 = n4845 | n4846;
  assign n4849 = ~n4847 & n4848;
  assign n4850 = n12217 & n4849;
  assign n4851 = n12217 | n4849;
  assign n4852 = ~n4850 & n4851;
  assign n4853 = x53 & x89;
  assign n4854 = n4852 & n4853;
  assign n4855 = n4852 | n4853;
  assign n4856 = ~n4854 & n4855;
  assign n4857 = n12215 & n4856;
  assign n4858 = n12215 | n4856;
  assign n4859 = ~n4857 & n4858;
  assign n4860 = x52 & x90;
  assign n4861 = n4859 & n4860;
  assign n4862 = n4859 | n4860;
  assign n4863 = ~n4861 & n4862;
  assign n4864 = n12213 & n4863;
  assign n4865 = n12213 | n4863;
  assign n4866 = ~n4864 & n4865;
  assign n4867 = x51 & x91;
  assign n4868 = n4866 & n4867;
  assign n4869 = n4866 | n4867;
  assign n4870 = ~n4868 & n4869;
  assign n4871 = n12211 & n4870;
  assign n4872 = n12211 | n4870;
  assign n4873 = ~n4871 & n4872;
  assign n4874 = x50 & x92;
  assign n4875 = n4873 & n4874;
  assign n4876 = n4873 | n4874;
  assign n4877 = ~n4875 & n4876;
  assign n4878 = n12209 & n4877;
  assign n4879 = n12209 | n4877;
  assign n4880 = ~n4878 & n4879;
  assign n4881 = x49 & x93;
  assign n4882 = n4880 & n4881;
  assign n4883 = n4880 | n4881;
  assign n4884 = ~n4882 & n4883;
  assign n4885 = n4781 & n4884;
  assign n4886 = n4781 | n4884;
  assign n4887 = ~n4885 & n4886;
  assign n4888 = x48 & x94;
  assign n4889 = n4887 & n4888;
  assign n4890 = n4887 | n4888;
  assign n4891 = ~n4889 & n4890;
  assign n17690 = n4780 | n4881;
  assign n17691 = (n4779 & n4881) | (n4779 & n17690) | (n4881 & n17690);
  assign n15746 = (n4781 & n4880) | (n4781 & n17691) | (n4880 & n17691);
  assign n12263 = (n4882 & n4884) | (n4882 & n15746) | (n4884 & n15746);
  assign n15747 = n4875 | n12209;
  assign n15748 = (n4875 & n4877) | (n4875 & n15747) | (n4877 & n15747);
  assign n4894 = n4868 | n4871;
  assign n4895 = n4861 | n4864;
  assign n12267 = n4819 | n4821;
  assign n15749 = n4718 | n4819;
  assign n15750 = (n4819 & n4821) | (n4819 & n15749) | (n4821 & n15749);
  assign n15751 = (n12194 & n12267) | (n12194 & n15750) | (n12267 & n15750);
  assign n15752 = (n4720 & n12267) | (n4720 & n15750) | (n12267 & n15750);
  assign n15753 = (n12166 & n15751) | (n12166 & n15752) | (n15751 & n15752);
  assign n15754 = n4805 | n4807;
  assign n15755 = (n4805 & n12222) | (n4805 & n15754) | (n12222 & n15754);
  assign n15756 = n4704 | n4805;
  assign n15757 = (n4805 & n4807) | (n4805 & n15756) | (n4807 & n15756);
  assign n15758 = (n15709 & n15755) | (n15709 & n15757) | (n15755 & n15757);
  assign n15759 = (n15711 & n15755) | (n15711 & n15757) | (n15755 & n15757);
  assign n15760 = (n15668 & n15758) | (n15668 & n15759) | (n15758 & n15759);
  assign n4905 = x63 & x80;
  assign n4906 = x62 & x81;
  assign n4907 = n4905 & n4906;
  assign n4908 = n4905 | n4906;
  assign n4909 = ~n4907 & n4908;
  assign n15761 = n4798 | n4800;
  assign n15762 = (n4798 & n12224) | (n4798 & n15761) | (n12224 & n15761);
  assign n12275 = n4909 & n15762;
  assign n15763 = n4697 | n4798;
  assign n15764 = (n4798 & n4800) | (n4798 & n15763) | (n4800 & n15763);
  assign n12276 = n4909 & n15764;
  assign n15765 = (n12275 & n12276) | (n12275 & n15713) | (n12276 & n15713);
  assign n15766 = (n12275 & n12276) | (n12275 & n15714) | (n12276 & n15714);
  assign n15767 = (n15651 & n15765) | (n15651 & n15766) | (n15765 & n15766);
  assign n12278 = n4909 | n15762;
  assign n12279 = n4909 | n15764;
  assign n15768 = (n12278 & n12279) | (n12278 & n15713) | (n12279 & n15713);
  assign n15769 = (n12278 & n12279) | (n12278 & n15714) | (n12279 & n15714);
  assign n15770 = (n15651 & n15768) | (n15651 & n15769) | (n15768 & n15769);
  assign n4912 = ~n15767 & n15770;
  assign n4913 = x61 & x82;
  assign n4914 = n4912 & n4913;
  assign n4915 = n4912 | n4913;
  assign n4916 = ~n4914 & n4915;
  assign n4917 = n15760 & n4916;
  assign n4918 = n15760 | n4916;
  assign n4919 = ~n4917 & n4918;
  assign n4920 = x60 & x83;
  assign n4921 = n4919 & n4920;
  assign n4922 = n4919 | n4920;
  assign n4923 = ~n4921 & n4922;
  assign n12281 = n4812 & n4923;
  assign n15771 = (n4923 & n12238) | (n4923 & n12281) | (n12238 & n12281);
  assign n15772 = (n4923 & n12239) | (n4923 & n12281) | (n12239 & n12281);
  assign n15773 = (n15707 & n15771) | (n15707 & n15772) | (n15771 & n15772);
  assign n12283 = n4812 | n4923;
  assign n15774 = n12238 | n12283;
  assign n15775 = n12239 | n12283;
  assign n15776 = (n15707 & n15774) | (n15707 & n15775) | (n15774 & n15775);
  assign n4926 = ~n15773 & n15776;
  assign n4927 = x59 & x84;
  assign n4928 = n4926 & n4927;
  assign n4929 = n4926 | n4927;
  assign n4930 = ~n4928 & n4929;
  assign n4931 = n15753 & n4930;
  assign n4932 = n15753 | n4930;
  assign n4933 = ~n4931 & n4932;
  assign n4934 = x58 & x85;
  assign n4935 = n4933 & n4934;
  assign n4936 = n4933 | n4934;
  assign n4937 = ~n4935 & n4936;
  assign n12285 = n4826 & n4937;
  assign n12286 = (n4937 & n12249) | (n4937 & n12285) | (n12249 & n12285);
  assign n12287 = n4826 | n4937;
  assign n12288 = n12249 | n12287;
  assign n4940 = ~n12286 & n12288;
  assign n4941 = x57 & x86;
  assign n4942 = n4940 & n4941;
  assign n4943 = n4940 | n4941;
  assign n4944 = ~n4942 & n4943;
  assign n12289 = n4833 & n4944;
  assign n12290 = (n4944 & n12253) | (n4944 & n12289) | (n12253 & n12289);
  assign n12291 = n4833 | n4944;
  assign n12292 = n12253 | n12291;
  assign n4947 = ~n12290 & n12292;
  assign n4948 = x56 & x87;
  assign n4949 = n4947 & n4948;
  assign n4950 = n4947 | n4948;
  assign n4951 = ~n4949 & n4950;
  assign n12293 = n4840 & n4951;
  assign n12294 = (n4951 & n12258) | (n4951 & n12293) | (n12258 & n12293);
  assign n12295 = n4840 | n4951;
  assign n12296 = n12258 | n12295;
  assign n4954 = ~n12294 & n12296;
  assign n4955 = x55 & x88;
  assign n4956 = n4954 & n4955;
  assign n4957 = n4954 | n4955;
  assign n4958 = ~n4956 & n4957;
  assign n12264 = n4847 | n4849;
  assign n12297 = n4958 & n12264;
  assign n12298 = n4847 & n4958;
  assign n12299 = (n12217 & n12297) | (n12217 & n12298) | (n12297 & n12298);
  assign n12300 = n4958 | n12264;
  assign n12301 = n4847 | n4958;
  assign n12302 = (n12217 & n12300) | (n12217 & n12301) | (n12300 & n12301);
  assign n4961 = ~n12299 & n12302;
  assign n4962 = x54 & x89;
  assign n4963 = n4961 & n4962;
  assign n4964 = n4961 | n4962;
  assign n4965 = ~n4963 & n4964;
  assign n12303 = n4854 & n4965;
  assign n12304 = (n4857 & n4965) | (n4857 & n12303) | (n4965 & n12303);
  assign n12305 = n4854 | n4965;
  assign n12306 = n4857 | n12305;
  assign n4968 = ~n12304 & n12306;
  assign n4969 = x53 & x90;
  assign n4970 = n4968 & n4969;
  assign n4971 = n4968 | n4969;
  assign n4972 = ~n4970 & n4971;
  assign n4973 = n4895 & n4972;
  assign n4974 = n4895 | n4972;
  assign n4975 = ~n4973 & n4974;
  assign n4976 = x52 & x91;
  assign n4977 = n4975 & n4976;
  assign n4978 = n4975 | n4976;
  assign n4979 = ~n4977 & n4978;
  assign n4980 = n4894 & n4979;
  assign n4981 = n4894 | n4979;
  assign n4982 = ~n4980 & n4981;
  assign n4983 = x51 & x92;
  assign n4984 = n4982 & n4983;
  assign n4985 = n4982 | n4983;
  assign n4986 = ~n4984 & n4985;
  assign n4987 = n15748 & n4986;
  assign n4988 = n15748 | n4986;
  assign n4989 = ~n4987 & n4988;
  assign n4990 = x50 & x93;
  assign n4991 = n4989 & n4990;
  assign n4992 = n4989 | n4990;
  assign n4993 = ~n4991 & n4992;
  assign n4994 = n12263 & n4993;
  assign n4995 = n12263 | n4993;
  assign n4996 = ~n4994 & n4995;
  assign n4997 = x49 & x94;
  assign n4998 = n4996 & n4997;
  assign n4999 = n4996 | n4997;
  assign n5000 = ~n4998 & n4999;
  assign n5001 = n4889 & n5000;
  assign n5002 = n4889 | n5000;
  assign n5003 = ~n5001 & n5002;
  assign n5004 = x48 & x95;
  assign n5005 = n5003 & n5004;
  assign n5006 = n5003 | n5004;
  assign n5007 = ~n5005 & n5006;
  assign n17692 = n4888 | n4997;
  assign n17693 = (n4887 & n4997) | (n4887 & n17692) | (n4997 & n17692);
  assign n15778 = (n4889 & n4996) | (n4889 & n17693) | (n4996 & n17693);
  assign n12308 = (n4998 & n5000) | (n4998 & n15778) | (n5000 & n15778);
  assign n12309 = n4991 | n12263;
  assign n12310 = (n4991 & n4993) | (n4991 & n12309) | (n4993 & n12309);
  assign n15779 = n4984 | n15748;
  assign n15780 = (n4984 & n4986) | (n4984 & n15779) | (n4986 & n15779);
  assign n5011 = n4977 | n4980;
  assign n12311 = n4970 | n4972;
  assign n12312 = (n4895 & n4970) | (n4895 & n12311) | (n4970 & n12311);
  assign n12316 = n4921 | n4923;
  assign n15781 = n4812 | n4921;
  assign n15782 = (n4921 & n4923) | (n4921 & n15781) | (n4923 & n15781);
  assign n15783 = (n12238 & n12316) | (n12238 & n15782) | (n12316 & n15782);
  assign n15784 = (n12239 & n12316) | (n12239 & n15782) | (n12316 & n15782);
  assign n15785 = (n15707 & n15783) | (n15707 & n15784) | (n15783 & n15784);
  assign n5022 = x64 & x80;
  assign n5023 = x63 & x81;
  assign n5024 = n5022 & n5023;
  assign n5025 = n5022 | n5023;
  assign n5026 = ~n5024 & n5025;
  assign n15786 = n4907 | n4909;
  assign n15791 = (n4907 & n15764) | (n4907 & n15786) | (n15764 & n15786);
  assign n12324 = n5026 & n15791;
  assign n15788 = n5026 & n15786;
  assign n15789 = n4907 & n5026;
  assign n15790 = (n15762 & n15788) | (n15762 & n15789) | (n15788 & n15789);
  assign n15792 = (n12324 & n15713) | (n12324 & n15790) | (n15713 & n15790);
  assign n15793 = (n12324 & n15714) | (n12324 & n15790) | (n15714 & n15790);
  assign n15794 = (n15651 & n15792) | (n15651 & n15793) | (n15792 & n15793);
  assign n12327 = n5026 | n15791;
  assign n15795 = n5026 | n15786;
  assign n15796 = n4907 | n5026;
  assign n15797 = (n15762 & n15795) | (n15762 & n15796) | (n15795 & n15796);
  assign n15798 = (n12327 & n15713) | (n12327 & n15797) | (n15713 & n15797);
  assign n15799 = (n12327 & n15714) | (n12327 & n15797) | (n15714 & n15797);
  assign n15800 = (n15651 & n15798) | (n15651 & n15799) | (n15798 & n15799);
  assign n5029 = ~n15794 & n15800;
  assign n5030 = x62 & x82;
  assign n5031 = n5029 & n5030;
  assign n5032 = n5029 | n5030;
  assign n5033 = ~n5031 & n5032;
  assign n12318 = n4914 | n4916;
  assign n12329 = n5033 & n12318;
  assign n12330 = n4914 & n5033;
  assign n12331 = (n15760 & n12329) | (n15760 & n12330) | (n12329 & n12330);
  assign n12332 = n5033 | n12318;
  assign n12333 = n4914 | n5033;
  assign n12334 = (n15760 & n12332) | (n15760 & n12333) | (n12332 & n12333);
  assign n5036 = ~n12331 & n12334;
  assign n5037 = x61 & x83;
  assign n5038 = n5036 & n5037;
  assign n5039 = n5036 | n5037;
  assign n5040 = ~n5038 & n5039;
  assign n5041 = n15785 & n5040;
  assign n5042 = n15785 | n5040;
  assign n5043 = ~n5041 & n5042;
  assign n5044 = x60 & x84;
  assign n5045 = n5043 & n5044;
  assign n5046 = n5043 | n5044;
  assign n5047 = ~n5045 & n5046;
  assign n12313 = n4928 | n4930;
  assign n12335 = n5047 & n12313;
  assign n12336 = n4928 & n5047;
  assign n12337 = (n15753 & n12335) | (n15753 & n12336) | (n12335 & n12336);
  assign n12338 = n5047 | n12313;
  assign n12339 = n4928 | n5047;
  assign n12340 = (n15753 & n12338) | (n15753 & n12339) | (n12338 & n12339);
  assign n5050 = ~n12337 & n12340;
  assign n5051 = x59 & x85;
  assign n5052 = n5050 & n5051;
  assign n5053 = n5050 | n5051;
  assign n5054 = ~n5052 & n5053;
  assign n12341 = n4935 & n5054;
  assign n15801 = (n5054 & n12285) | (n5054 & n12341) | (n12285 & n12341);
  assign n15802 = (n4937 & n5054) | (n4937 & n12341) | (n5054 & n12341);
  assign n15803 = (n12249 & n15801) | (n12249 & n15802) | (n15801 & n15802);
  assign n12343 = n4935 | n5054;
  assign n15804 = n12285 | n12343;
  assign n15805 = n4937 | n12343;
  assign n15806 = (n12249 & n15804) | (n12249 & n15805) | (n15804 & n15805);
  assign n5057 = ~n15803 & n15806;
  assign n5058 = x58 & x86;
  assign n5059 = n5057 & n5058;
  assign n5060 = n5057 | n5058;
  assign n5061 = ~n5059 & n5060;
  assign n12345 = n4942 & n5061;
  assign n12346 = (n5061 & n12290) | (n5061 & n12345) | (n12290 & n12345);
  assign n12347 = n4942 | n5061;
  assign n12348 = n12290 | n12347;
  assign n5064 = ~n12346 & n12348;
  assign n5065 = x57 & x87;
  assign n5066 = n5064 & n5065;
  assign n5067 = n5064 | n5065;
  assign n5068 = ~n5066 & n5067;
  assign n12349 = n4949 & n5068;
  assign n12350 = (n5068 & n12294) | (n5068 & n12349) | (n12294 & n12349);
  assign n12351 = n4949 | n5068;
  assign n12352 = n12294 | n12351;
  assign n5071 = ~n12350 & n12352;
  assign n5072 = x56 & x88;
  assign n5073 = n5071 & n5072;
  assign n5074 = n5071 | n5072;
  assign n5075 = ~n5073 & n5074;
  assign n12353 = n4956 & n5075;
  assign n12354 = (n5075 & n12299) | (n5075 & n12353) | (n12299 & n12353);
  assign n12355 = n4956 | n5075;
  assign n12356 = n12299 | n12355;
  assign n5078 = ~n12354 & n12356;
  assign n5079 = x55 & x89;
  assign n5080 = n5078 & n5079;
  assign n5081 = n5078 | n5079;
  assign n5082 = ~n5080 & n5081;
  assign n12357 = n4963 & n5082;
  assign n12358 = (n5082 & n12304) | (n5082 & n12357) | (n12304 & n12357);
  assign n12359 = n4963 | n5082;
  assign n12360 = n12304 | n12359;
  assign n5085 = ~n12358 & n12360;
  assign n5086 = x54 & x90;
  assign n5087 = n5085 & n5086;
  assign n5088 = n5085 | n5086;
  assign n5089 = ~n5087 & n5088;
  assign n5090 = n12312 & n5089;
  assign n5091 = n12312 | n5089;
  assign n5092 = ~n5090 & n5091;
  assign n5093 = x53 & x91;
  assign n5094 = n5092 & n5093;
  assign n5095 = n5092 | n5093;
  assign n5096 = ~n5094 & n5095;
  assign n5097 = n5011 & n5096;
  assign n5098 = n5011 | n5096;
  assign n5099 = ~n5097 & n5098;
  assign n5100 = x52 & x92;
  assign n5101 = n5099 & n5100;
  assign n5102 = n5099 | n5100;
  assign n5103 = ~n5101 & n5102;
  assign n5104 = n15780 & n5103;
  assign n5105 = n15780 | n5103;
  assign n5106 = ~n5104 & n5105;
  assign n5107 = x51 & x93;
  assign n5108 = n5106 & n5107;
  assign n5109 = n5106 | n5107;
  assign n5110 = ~n5108 & n5109;
  assign n5111 = n12310 & n5110;
  assign n5112 = n12310 | n5110;
  assign n5113 = ~n5111 & n5112;
  assign n5114 = x50 & x94;
  assign n5115 = n5113 & n5114;
  assign n5116 = n5113 | n5114;
  assign n5117 = ~n5115 & n5116;
  assign n5118 = n12308 & n5117;
  assign n5119 = n12308 | n5117;
  assign n5120 = ~n5118 & n5119;
  assign n5121 = x49 & x95;
  assign n5122 = n5120 & n5121;
  assign n5123 = n5120 | n5121;
  assign n5124 = ~n5122 & n5123;
  assign n5125 = n5005 & n5124;
  assign n5126 = n5005 | n5124;
  assign n5127 = ~n5125 & n5126;
  assign n5128 = x48 & x96;
  assign n5129 = n5127 & n5128;
  assign n5130 = n5127 | n5128;
  assign n5131 = ~n5129 & n5130;
  assign n17694 = n5004 | n5121;
  assign n17695 = (n5003 & n5121) | (n5003 & n17694) | (n5121 & n17694);
  assign n15808 = (n5005 & n5120) | (n5005 & n17695) | (n5120 & n17695);
  assign n12362 = (n5122 & n5124) | (n5122 & n15808) | (n5124 & n15808);
  assign n12363 = n5115 | n12308;
  assign n12364 = (n5115 & n5117) | (n5115 & n12363) | (n5117 & n12363);
  assign n12365 = n5108 | n12310;
  assign n12366 = (n5108 & n5110) | (n5108 & n12365) | (n5110 & n12365);
  assign n15809 = n5101 | n15780;
  assign n15810 = (n5101 & n5103) | (n5101 & n15809) | (n5103 & n15809);
  assign n12367 = n5094 | n5096;
  assign n12368 = (n5011 & n5094) | (n5011 & n12367) | (n5094 & n12367);
  assign n12369 = n5087 | n5089;
  assign n12370 = (n5087 & n12312) | (n5087 & n12369) | (n12312 & n12369);
  assign n12372 = n5052 | n5054;
  assign n15811 = n4935 | n5052;
  assign n15812 = (n5052 & n5054) | (n5052 & n15811) | (n5054 & n15811);
  assign n15813 = (n12285 & n12372) | (n12285 & n15812) | (n12372 & n15812);
  assign n15814 = (n4937 & n12372) | (n4937 & n15812) | (n12372 & n15812);
  assign n15815 = (n12249 & n15813) | (n12249 & n15814) | (n15813 & n15814);
  assign n5147 = x65 & x80;
  assign n5148 = x64 & x81;
  assign n5149 = n5147 & n5148;
  assign n5150 = n5147 | n5148;
  assign n5151 = ~n5149 & n5150;
  assign n12379 = n5024 & n5151;
  assign n12380 = (n5151 & n15794) | (n5151 & n12379) | (n15794 & n12379);
  assign n12381 = n5024 | n5151;
  assign n12382 = n15794 | n12381;
  assign n5154 = ~n12380 & n12382;
  assign n5155 = x63 & x82;
  assign n5156 = n5154 & n5155;
  assign n5157 = n5154 | n5155;
  assign n5158 = ~n5156 & n5157;
  assign n15816 = n5031 | n5033;
  assign n15817 = (n5031 & n12318) | (n5031 & n15816) | (n12318 & n15816);
  assign n12383 = n5158 & n15817;
  assign n15818 = n4914 | n5031;
  assign n15819 = (n5031 & n5033) | (n5031 & n15818) | (n5033 & n15818);
  assign n12384 = n5158 & n15819;
  assign n12385 = (n15760 & n12383) | (n15760 & n12384) | (n12383 & n12384);
  assign n12386 = n5158 | n15817;
  assign n12387 = n5158 | n15819;
  assign n12388 = (n15760 & n12386) | (n15760 & n12387) | (n12386 & n12387);
  assign n5161 = ~n12385 & n12388;
  assign n5162 = x62 & x83;
  assign n5163 = n5161 & n5162;
  assign n5164 = n5161 | n5162;
  assign n5165 = ~n5163 & n5164;
  assign n12374 = n5038 | n5040;
  assign n12389 = n5165 & n12374;
  assign n12390 = n5038 & n5165;
  assign n12391 = (n15785 & n12389) | (n15785 & n12390) | (n12389 & n12390);
  assign n12392 = n5165 | n12374;
  assign n12393 = n5038 | n5165;
  assign n12394 = (n15785 & n12392) | (n15785 & n12393) | (n12392 & n12393);
  assign n5168 = ~n12391 & n12394;
  assign n5169 = x61 & x84;
  assign n5170 = n5168 & n5169;
  assign n5171 = n5168 | n5169;
  assign n5172 = ~n5170 & n5171;
  assign n12395 = n5045 & n5172;
  assign n15820 = (n5172 & n12336) | (n5172 & n12395) | (n12336 & n12395);
  assign n15821 = (n5172 & n12335) | (n5172 & n12395) | (n12335 & n12395);
  assign n15822 = (n15753 & n15820) | (n15753 & n15821) | (n15820 & n15821);
  assign n12397 = n5045 | n5172;
  assign n15823 = n12336 | n12397;
  assign n15824 = n12335 | n12397;
  assign n15825 = (n15753 & n15823) | (n15753 & n15824) | (n15823 & n15824);
  assign n5175 = ~n15822 & n15825;
  assign n5176 = x60 & x85;
  assign n5177 = n5175 & n5176;
  assign n5178 = n5175 | n5176;
  assign n5179 = ~n5177 & n5178;
  assign n5180 = n15815 & n5179;
  assign n5181 = n15815 | n5179;
  assign n5182 = ~n5180 & n5181;
  assign n5183 = x59 & x86;
  assign n5184 = n5182 & n5183;
  assign n5185 = n5182 | n5183;
  assign n5186 = ~n5184 & n5185;
  assign n12399 = n5059 & n5186;
  assign n12400 = (n5186 & n12346) | (n5186 & n12399) | (n12346 & n12399);
  assign n12401 = n5059 | n5186;
  assign n12402 = n12346 | n12401;
  assign n5189 = ~n12400 & n12402;
  assign n5190 = x58 & x87;
  assign n5191 = n5189 & n5190;
  assign n5192 = n5189 | n5190;
  assign n5193 = ~n5191 & n5192;
  assign n12403 = n5066 & n5193;
  assign n12404 = (n5193 & n12350) | (n5193 & n12403) | (n12350 & n12403);
  assign n12405 = n5066 | n5193;
  assign n12406 = n12350 | n12405;
  assign n5196 = ~n12404 & n12406;
  assign n5197 = x57 & x88;
  assign n5198 = n5196 & n5197;
  assign n5199 = n5196 | n5197;
  assign n5200 = ~n5198 & n5199;
  assign n12407 = n5073 & n5200;
  assign n12408 = (n5200 & n12354) | (n5200 & n12407) | (n12354 & n12407);
  assign n12409 = n5073 | n5200;
  assign n12410 = n12354 | n12409;
  assign n5203 = ~n12408 & n12410;
  assign n5204 = x56 & x89;
  assign n5205 = n5203 & n5204;
  assign n5206 = n5203 | n5204;
  assign n5207 = ~n5205 & n5206;
  assign n12411 = n5080 & n5207;
  assign n12412 = (n5207 & n12358) | (n5207 & n12411) | (n12358 & n12411);
  assign n12413 = n5080 | n5207;
  assign n12414 = n12358 | n12413;
  assign n5210 = ~n12412 & n12414;
  assign n5211 = x55 & x90;
  assign n5212 = n5210 & n5211;
  assign n5213 = n5210 | n5211;
  assign n5214 = ~n5212 & n5213;
  assign n5215 = n12370 & n5214;
  assign n5216 = n12370 | n5214;
  assign n5217 = ~n5215 & n5216;
  assign n5218 = x54 & x91;
  assign n5219 = n5217 & n5218;
  assign n5220 = n5217 | n5218;
  assign n5221 = ~n5219 & n5220;
  assign n5222 = n12368 & n5221;
  assign n5223 = n12368 | n5221;
  assign n5224 = ~n5222 & n5223;
  assign n5225 = x53 & x92;
  assign n5226 = n5224 & n5225;
  assign n5227 = n5224 | n5225;
  assign n5228 = ~n5226 & n5227;
  assign n5229 = n15810 & n5228;
  assign n5230 = n15810 | n5228;
  assign n5231 = ~n5229 & n5230;
  assign n5232 = x52 & x93;
  assign n5233 = n5231 & n5232;
  assign n5234 = n5231 | n5232;
  assign n5235 = ~n5233 & n5234;
  assign n5236 = n12366 & n5235;
  assign n5237 = n12366 | n5235;
  assign n5238 = ~n5236 & n5237;
  assign n5239 = x51 & x94;
  assign n5240 = n5238 & n5239;
  assign n5241 = n5238 | n5239;
  assign n5242 = ~n5240 & n5241;
  assign n5243 = n12364 & n5242;
  assign n5244 = n12364 | n5242;
  assign n5245 = ~n5243 & n5244;
  assign n5246 = x50 & x95;
  assign n5247 = n5245 & n5246;
  assign n5248 = n5245 | n5246;
  assign n5249 = ~n5247 & n5248;
  assign n5250 = n12362 & n5249;
  assign n5251 = n12362 | n5249;
  assign n5252 = ~n5250 & n5251;
  assign n5253 = x49 & x96;
  assign n5254 = n5252 & n5253;
  assign n5255 = n5252 | n5253;
  assign n5256 = ~n5254 & n5255;
  assign n5257 = n5129 & n5256;
  assign n5258 = n5129 | n5256;
  assign n5259 = ~n5257 & n5258;
  assign n5260 = x48 & x97;
  assign n5261 = n5259 & n5260;
  assign n5262 = n5259 | n5260;
  assign n5263 = ~n5261 & n5262;
  assign n12415 = n5129 | n5254;
  assign n12416 = (n5254 & n5256) | (n5254 & n12415) | (n5256 & n12415);
  assign n12417 = n5247 | n12362;
  assign n12418 = (n5247 & n5249) | (n5247 & n12417) | (n5249 & n12417);
  assign n12419 = n5240 | n12364;
  assign n12420 = (n5240 & n5242) | (n5240 & n12419) | (n5242 & n12419);
  assign n12421 = n5233 | n12366;
  assign n12422 = (n5233 & n5235) | (n5233 & n12421) | (n5235 & n12421);
  assign n12423 = n5226 | n5228;
  assign n12424 = (n15810 & n5226) | (n15810 & n12423) | (n5226 & n12423);
  assign n12425 = n5219 | n5221;
  assign n12426 = (n5219 & n12368) | (n5219 & n12425) | (n12368 & n12425);
  assign n12427 = n5212 | n5214;
  assign n12428 = (n5212 & n12370) | (n5212 & n12427) | (n12370 & n12427);
  assign n12432 = n5170 | n5172;
  assign n15826 = n5045 | n5170;
  assign n15827 = (n5170 & n5172) | (n5170 & n15826) | (n5172 & n15826);
  assign n15828 = (n12336 & n12432) | (n12336 & n15827) | (n12432 & n15827);
  assign n15829 = (n12335 & n12432) | (n12335 & n15827) | (n12432 & n15827);
  assign n15830 = (n15753 & n15828) | (n15753 & n15829) | (n15828 & n15829);
  assign n5280 = x66 & x80;
  assign n5281 = x65 & x81;
  assign n5282 = n5280 & n5281;
  assign n5283 = n5280 | n5281;
  assign n5284 = ~n5282 & n5283;
  assign n15835 = n5024 | n5149;
  assign n15836 = (n5149 & n5151) | (n5149 & n15835) | (n5151 & n15835);
  assign n12440 = n5284 & n15836;
  assign n12438 = n5149 | n5151;
  assign n12441 = n5284 & n12438;
  assign n12442 = (n15794 & n12440) | (n15794 & n12441) | (n12440 & n12441);
  assign n12443 = n5284 | n15836;
  assign n12444 = n5284 | n12438;
  assign n12445 = (n15794 & n12443) | (n15794 & n12444) | (n12443 & n12444);
  assign n5287 = ~n12442 & n12445;
  assign n5288 = x64 & x82;
  assign n5289 = n5287 & n5288;
  assign n5290 = n5287 | n5288;
  assign n5291 = ~n5289 & n5290;
  assign n12446 = n5156 & n5291;
  assign n15837 = (n5291 & n12383) | (n5291 & n12446) | (n12383 & n12446);
  assign n15838 = (n5291 & n12384) | (n5291 & n12446) | (n12384 & n12446);
  assign n15839 = (n15760 & n15837) | (n15760 & n15838) | (n15837 & n15838);
  assign n12448 = n5156 | n5291;
  assign n15840 = n12383 | n12448;
  assign n15841 = n12384 | n12448;
  assign n15842 = (n15760 & n15840) | (n15760 & n15841) | (n15840 & n15841);
  assign n5294 = ~n15839 & n15842;
  assign n5295 = x63 & x83;
  assign n5296 = n5294 & n5295;
  assign n5297 = n5294 | n5295;
  assign n5298 = ~n5296 & n5297;
  assign n15831 = n5163 | n5165;
  assign n15832 = (n5163 & n12374) | (n5163 & n15831) | (n12374 & n15831);
  assign n15843 = n5298 & n15832;
  assign n15833 = n5038 | n5163;
  assign n15834 = (n5163 & n5165) | (n5163 & n15833) | (n5165 & n15833);
  assign n15844 = n5298 & n15834;
  assign n15845 = (n15785 & n15843) | (n15785 & n15844) | (n15843 & n15844);
  assign n15846 = n5298 | n15832;
  assign n15847 = n5298 | n15834;
  assign n15848 = (n15785 & n15846) | (n15785 & n15847) | (n15846 & n15847);
  assign n5301 = ~n15845 & n15848;
  assign n5302 = x62 & x84;
  assign n5303 = n5301 & n5302;
  assign n5304 = n5301 | n5302;
  assign n5305 = ~n5303 & n5304;
  assign n5306 = n15830 & n5305;
  assign n5307 = n15830 | n5305;
  assign n5308 = ~n5306 & n5307;
  assign n5309 = x61 & x85;
  assign n5310 = n5308 & n5309;
  assign n5311 = n5308 | n5309;
  assign n5312 = ~n5310 & n5311;
  assign n12429 = n5177 | n5179;
  assign n12450 = n5312 & n12429;
  assign n12451 = n5177 & n5312;
  assign n12452 = (n15815 & n12450) | (n15815 & n12451) | (n12450 & n12451);
  assign n12453 = n5312 | n12429;
  assign n12454 = n5177 | n5312;
  assign n12455 = (n15815 & n12453) | (n15815 & n12454) | (n12453 & n12454);
  assign n5315 = ~n12452 & n12455;
  assign n5316 = x60 & x86;
  assign n5317 = n5315 & n5316;
  assign n5318 = n5315 | n5316;
  assign n5319 = ~n5317 & n5318;
  assign n12456 = n5184 & n5319;
  assign n15849 = (n5319 & n12399) | (n5319 & n12456) | (n12399 & n12456);
  assign n15850 = (n5186 & n5319) | (n5186 & n12456) | (n5319 & n12456);
  assign n15851 = (n12346 & n15849) | (n12346 & n15850) | (n15849 & n15850);
  assign n12458 = n5184 | n5319;
  assign n15852 = n12399 | n12458;
  assign n15853 = n5186 | n12458;
  assign n15854 = (n12346 & n15852) | (n12346 & n15853) | (n15852 & n15853);
  assign n5322 = ~n15851 & n15854;
  assign n5323 = x59 & x87;
  assign n5324 = n5322 & n5323;
  assign n5325 = n5322 | n5323;
  assign n5326 = ~n5324 & n5325;
  assign n12460 = n5191 & n5326;
  assign n12461 = (n5326 & n12404) | (n5326 & n12460) | (n12404 & n12460);
  assign n12462 = n5191 | n5326;
  assign n12463 = n12404 | n12462;
  assign n5329 = ~n12461 & n12463;
  assign n5330 = x58 & x88;
  assign n5331 = n5329 & n5330;
  assign n5332 = n5329 | n5330;
  assign n5333 = ~n5331 & n5332;
  assign n12464 = n5198 & n5333;
  assign n12465 = (n5333 & n12408) | (n5333 & n12464) | (n12408 & n12464);
  assign n12466 = n5198 | n5333;
  assign n12467 = n12408 | n12466;
  assign n5336 = ~n12465 & n12467;
  assign n5337 = x57 & x89;
  assign n5338 = n5336 & n5337;
  assign n5339 = n5336 | n5337;
  assign n5340 = ~n5338 & n5339;
  assign n12468 = n5205 & n5340;
  assign n12469 = (n5340 & n12412) | (n5340 & n12468) | (n12412 & n12468);
  assign n12470 = n5205 | n5340;
  assign n12471 = n12412 | n12470;
  assign n5343 = ~n12469 & n12471;
  assign n5344 = x56 & x90;
  assign n5345 = n5343 & n5344;
  assign n5346 = n5343 | n5344;
  assign n5347 = ~n5345 & n5346;
  assign n5348 = n12428 & n5347;
  assign n5349 = n12428 | n5347;
  assign n5350 = ~n5348 & n5349;
  assign n5351 = x55 & x91;
  assign n5352 = n5350 & n5351;
  assign n5353 = n5350 | n5351;
  assign n5354 = ~n5352 & n5353;
  assign n5355 = n12426 & n5354;
  assign n5356 = n12426 | n5354;
  assign n5357 = ~n5355 & n5356;
  assign n5358 = x54 & x92;
  assign n5359 = n5357 & n5358;
  assign n5360 = n5357 | n5358;
  assign n5361 = ~n5359 & n5360;
  assign n5362 = n12424 & n5361;
  assign n5363 = n12424 | n5361;
  assign n5364 = ~n5362 & n5363;
  assign n5365 = x53 & x93;
  assign n5366 = n5364 & n5365;
  assign n5367 = n5364 | n5365;
  assign n5368 = ~n5366 & n5367;
  assign n5369 = n12422 & n5368;
  assign n5370 = n12422 | n5368;
  assign n5371 = ~n5369 & n5370;
  assign n5372 = x52 & x94;
  assign n5373 = n5371 & n5372;
  assign n5374 = n5371 | n5372;
  assign n5375 = ~n5373 & n5374;
  assign n5376 = n12420 & n5375;
  assign n5377 = n12420 | n5375;
  assign n5378 = ~n5376 & n5377;
  assign n5379 = x51 & x95;
  assign n5380 = n5378 & n5379;
  assign n5381 = n5378 | n5379;
  assign n5382 = ~n5380 & n5381;
  assign n5383 = n12418 & n5382;
  assign n5384 = n12418 | n5382;
  assign n5385 = ~n5383 & n5384;
  assign n5386 = x50 & x96;
  assign n5387 = n5385 & n5386;
  assign n5388 = n5385 | n5386;
  assign n5389 = ~n5387 & n5388;
  assign n5390 = n12416 & n5389;
  assign n5391 = n12416 | n5389;
  assign n5392 = ~n5390 & n5391;
  assign n5393 = x49 & x97;
  assign n5394 = n5392 & n5393;
  assign n5395 = n5392 | n5393;
  assign n5396 = ~n5394 & n5395;
  assign n5397 = n5261 & n5396;
  assign n5398 = n5261 | n5396;
  assign n5399 = ~n5397 & n5398;
  assign n5400 = x48 & x98;
  assign n5401 = n5399 & n5400;
  assign n5402 = n5399 | n5400;
  assign n5403 = ~n5401 & n5402;
  assign n17696 = n5260 | n5393;
  assign n17697 = (n5259 & n5393) | (n5259 & n17696) | (n5393 & n17696);
  assign n15856 = (n5261 & n5392) | (n5261 & n17697) | (n5392 & n17697);
  assign n12473 = (n5394 & n5396) | (n5394 & n15856) | (n5396 & n15856);
  assign n15857 = n5387 | n12416;
  assign n15858 = (n5387 & n5389) | (n5387 & n15857) | (n5389 & n15857);
  assign n5406 = n5380 | n5383;
  assign n5407 = n5373 | n5376;
  assign n5408 = n5366 | n5369;
  assign n12474 = n5359 | n5361;
  assign n12475 = (n5359 & n12424) | (n5359 & n12474) | (n12424 & n12474);
  assign n12476 = n5352 | n5354;
  assign n12477 = (n5352 & n12426) | (n5352 & n12476) | (n12426 & n12476);
  assign n12478 = n5345 | n5347;
  assign n12479 = (n5345 & n12428) | (n5345 & n12478) | (n12428 & n12478);
  assign n12481 = n5317 | n5319;
  assign n15859 = n5184 | n5317;
  assign n15860 = (n5317 & n5319) | (n5317 & n15859) | (n5319 & n15859);
  assign n15861 = (n12399 & n12481) | (n12399 & n15860) | (n12481 & n15860);
  assign n15862 = (n5186 & n12481) | (n5186 & n15860) | (n12481 & n15860);
  assign n15863 = (n12346 & n15861) | (n12346 & n15862) | (n15861 & n15862);
  assign n5421 = x67 & x80;
  assign n5422 = x66 & x81;
  assign n5423 = n5421 & n5422;
  assign n5424 = n5421 | n5422;
  assign n5425 = ~n5423 & n5424;
  assign n15864 = n5282 | n5284;
  assign n15865 = (n5282 & n15836) | (n5282 & n15864) | (n15836 & n15864);
  assign n12493 = n5425 & n15865;
  assign n15866 = (n5282 & n12438) | (n5282 & n15864) | (n12438 & n15864);
  assign n12494 = n5425 & n15866;
  assign n12495 = (n15794 & n12493) | (n15794 & n12494) | (n12493 & n12494);
  assign n12496 = n5425 | n15865;
  assign n12497 = n5425 | n15866;
  assign n12498 = (n15794 & n12496) | (n15794 & n12497) | (n12496 & n12497);
  assign n5428 = ~n12495 & n12498;
  assign n5429 = x65 & x82;
  assign n5430 = n5428 & n5429;
  assign n5431 = n5428 | n5429;
  assign n5432 = ~n5430 & n5431;
  assign n15867 = n5156 | n5289;
  assign n15868 = (n5289 & n5291) | (n5289 & n15867) | (n5291 & n15867);
  assign n12499 = n5432 & n15868;
  assign n12488 = n5289 | n5291;
  assign n12500 = n5432 & n12488;
  assign n15869 = (n12383 & n12499) | (n12383 & n12500) | (n12499 & n12500);
  assign n15870 = (n12384 & n12499) | (n12384 & n12500) | (n12499 & n12500);
  assign n15871 = (n15760 & n15869) | (n15760 & n15870) | (n15869 & n15870);
  assign n12502 = n5432 | n15868;
  assign n12503 = n5432 | n12488;
  assign n15872 = (n12383 & n12502) | (n12383 & n12503) | (n12502 & n12503);
  assign n15873 = (n12384 & n12502) | (n12384 & n12503) | (n12502 & n12503);
  assign n15874 = (n15760 & n15872) | (n15760 & n15873) | (n15872 & n15873);
  assign n5435 = ~n15871 & n15874;
  assign n5436 = x64 & x83;
  assign n5437 = n5435 & n5436;
  assign n5438 = n5435 | n5436;
  assign n5439 = ~n5437 & n5438;
  assign n12485 = n5296 | n5298;
  assign n12505 = n5439 & n12485;
  assign n12506 = n5296 & n5439;
  assign n15875 = (n12505 & n12506) | (n12505 & n15832) | (n12506 & n15832);
  assign n15876 = (n12505 & n12506) | (n12505 & n15834) | (n12506 & n15834);
  assign n15877 = (n15785 & n15875) | (n15785 & n15876) | (n15875 & n15876);
  assign n12508 = n5439 | n12485;
  assign n12509 = n5296 | n5439;
  assign n15878 = (n12508 & n12509) | (n12508 & n15832) | (n12509 & n15832);
  assign n15879 = (n12508 & n12509) | (n12508 & n15834) | (n12509 & n15834);
  assign n15880 = (n15785 & n15878) | (n15785 & n15879) | (n15878 & n15879);
  assign n5442 = ~n15877 & n15880;
  assign n5443 = x63 & x84;
  assign n5444 = n5442 & n5443;
  assign n5445 = n5442 | n5443;
  assign n5446 = ~n5444 & n5445;
  assign n12483 = n5303 | n5305;
  assign n12511 = n5446 & n12483;
  assign n12512 = n5303 & n5446;
  assign n12513 = (n15830 & n12511) | (n15830 & n12512) | (n12511 & n12512);
  assign n12514 = n5446 | n12483;
  assign n12515 = n5303 | n5446;
  assign n12516 = (n15830 & n12514) | (n15830 & n12515) | (n12514 & n12515);
  assign n5449 = ~n12513 & n12516;
  assign n5450 = x62 & x85;
  assign n5451 = n5449 & n5450;
  assign n5452 = n5449 | n5450;
  assign n5453 = ~n5451 & n5452;
  assign n12517 = n5310 & n5453;
  assign n15881 = (n5453 & n12451) | (n5453 & n12517) | (n12451 & n12517);
  assign n15882 = (n5453 & n12450) | (n5453 & n12517) | (n12450 & n12517);
  assign n15883 = (n15815 & n15881) | (n15815 & n15882) | (n15881 & n15882);
  assign n12519 = n5310 | n5453;
  assign n15884 = n12451 | n12519;
  assign n15885 = n12450 | n12519;
  assign n15886 = (n15815 & n15884) | (n15815 & n15885) | (n15884 & n15885);
  assign n5456 = ~n15883 & n15886;
  assign n5457 = x61 & x86;
  assign n5458 = n5456 & n5457;
  assign n5459 = n5456 | n5457;
  assign n5460 = ~n5458 & n5459;
  assign n5461 = n15863 & n5460;
  assign n5462 = n15863 | n5460;
  assign n5463 = ~n5461 & n5462;
  assign n5464 = x60 & x87;
  assign n5465 = n5463 & n5464;
  assign n5466 = n5463 | n5464;
  assign n5467 = ~n5465 & n5466;
  assign n12521 = n5324 & n5467;
  assign n12522 = (n5467 & n12461) | (n5467 & n12521) | (n12461 & n12521);
  assign n12523 = n5324 | n5467;
  assign n12524 = n12461 | n12523;
  assign n5470 = ~n12522 & n12524;
  assign n5471 = x59 & x88;
  assign n5472 = n5470 & n5471;
  assign n5473 = n5470 | n5471;
  assign n5474 = ~n5472 & n5473;
  assign n12525 = n5331 & n5474;
  assign n12526 = (n5474 & n12465) | (n5474 & n12525) | (n12465 & n12525);
  assign n12527 = n5331 | n5474;
  assign n12528 = n12465 | n12527;
  assign n5477 = ~n12526 & n12528;
  assign n5478 = x58 & x89;
  assign n5479 = n5477 & n5478;
  assign n5480 = n5477 | n5478;
  assign n5481 = ~n5479 & n5480;
  assign n12529 = n5338 & n5481;
  assign n12530 = (n5481 & n12469) | (n5481 & n12529) | (n12469 & n12529);
  assign n12531 = n5338 | n5481;
  assign n12532 = n12469 | n12531;
  assign n5484 = ~n12530 & n12532;
  assign n5485 = x57 & x90;
  assign n5486 = n5484 & n5485;
  assign n5487 = n5484 | n5485;
  assign n5488 = ~n5486 & n5487;
  assign n5489 = n12479 & n5488;
  assign n5490 = n12479 | n5488;
  assign n5491 = ~n5489 & n5490;
  assign n5492 = x56 & x91;
  assign n5493 = n5491 & n5492;
  assign n5494 = n5491 | n5492;
  assign n5495 = ~n5493 & n5494;
  assign n5496 = n12477 & n5495;
  assign n5497 = n12477 | n5495;
  assign n5498 = ~n5496 & n5497;
  assign n5499 = x55 & x92;
  assign n5500 = n5498 & n5499;
  assign n5501 = n5498 | n5499;
  assign n5502 = ~n5500 & n5501;
  assign n5503 = n12475 & n5502;
  assign n5504 = n12475 | n5502;
  assign n5505 = ~n5503 & n5504;
  assign n5506 = x54 & x93;
  assign n5507 = n5505 & n5506;
  assign n5508 = n5505 | n5506;
  assign n5509 = ~n5507 & n5508;
  assign n5510 = n5408 & n5509;
  assign n5511 = n5408 | n5509;
  assign n5512 = ~n5510 & n5511;
  assign n5513 = x53 & x94;
  assign n5514 = n5512 & n5513;
  assign n5515 = n5512 | n5513;
  assign n5516 = ~n5514 & n5515;
  assign n5517 = n5407 & n5516;
  assign n5518 = n5407 | n5516;
  assign n5519 = ~n5517 & n5518;
  assign n5520 = x52 & x95;
  assign n5521 = n5519 & n5520;
  assign n5522 = n5519 | n5520;
  assign n5523 = ~n5521 & n5522;
  assign n5524 = n5406 & n5523;
  assign n5525 = n5406 | n5523;
  assign n5526 = ~n5524 & n5525;
  assign n5527 = x51 & x96;
  assign n5528 = n5526 & n5527;
  assign n5529 = n5526 | n5527;
  assign n5530 = ~n5528 & n5529;
  assign n5531 = n15858 & n5530;
  assign n5532 = n15858 | n5530;
  assign n5533 = ~n5531 & n5532;
  assign n5534 = x50 & x97;
  assign n5535 = n5533 & n5534;
  assign n5536 = n5533 | n5534;
  assign n5537 = ~n5535 & n5536;
  assign n5538 = n12473 & n5537;
  assign n5539 = n12473 | n5537;
  assign n5540 = ~n5538 & n5539;
  assign n5541 = x49 & x98;
  assign n5542 = n5540 & n5541;
  assign n5543 = n5540 | n5541;
  assign n5544 = ~n5542 & n5543;
  assign n5545 = n5401 & n5544;
  assign n5546 = n5401 | n5544;
  assign n5547 = ~n5545 & n5546;
  assign n5548 = x48 & x99;
  assign n5549 = n5547 & n5548;
  assign n5550 = n5547 | n5548;
  assign n5551 = ~n5549 & n5550;
  assign n17698 = n5400 | n5541;
  assign n17699 = (n5399 & n5541) | (n5399 & n17698) | (n5541 & n17698);
  assign n15888 = (n5401 & n5540) | (n5401 & n17699) | (n5540 & n17699);
  assign n12534 = (n5542 & n5544) | (n5542 & n15888) | (n5544 & n15888);
  assign n12535 = n5535 | n12473;
  assign n12536 = (n5535 & n5537) | (n5535 & n12535) | (n5537 & n12535);
  assign n15889 = n5528 | n15858;
  assign n15890 = (n5528 & n5530) | (n5528 & n15889) | (n5530 & n15889);
  assign n5555 = n5521 | n5524;
  assign n5556 = n5514 | n5517;
  assign n12537 = n5507 | n5509;
  assign n12538 = (n5408 & n5507) | (n5408 & n12537) | (n5507 & n12537);
  assign n12539 = n5500 | n5502;
  assign n12540 = (n5500 & n12475) | (n5500 & n12539) | (n12475 & n12539);
  assign n12541 = n5493 | n5495;
  assign n12542 = (n5493 & n12477) | (n5493 & n12541) | (n12477 & n12541);
  assign n12543 = n5486 | n5488;
  assign n12544 = (n5486 & n12479) | (n5486 & n12543) | (n12479 & n12543);
  assign n12548 = n5451 | n5453;
  assign n15891 = n5310 | n5451;
  assign n15892 = (n5451 & n5453) | (n5451 & n15891) | (n5453 & n15891);
  assign n15893 = (n12451 & n12548) | (n12451 & n15892) | (n12548 & n15892);
  assign n15894 = (n12450 & n12548) | (n12450 & n15892) | (n12548 & n15892);
  assign n15895 = (n15815 & n15893) | (n15815 & n15894) | (n15893 & n15894);
  assign n15896 = n5437 | n5439;
  assign n15897 = (n5437 & n12485) | (n5437 & n15896) | (n12485 & n15896);
  assign n15898 = n5296 | n5437;
  assign n15899 = (n5437 & n5439) | (n5437 & n15898) | (n5439 & n15898);
  assign n15900 = (n15832 & n15897) | (n15832 & n15899) | (n15897 & n15899);
  assign n15901 = (n15834 & n15897) | (n15834 & n15899) | (n15897 & n15899);
  assign n15902 = (n15785 & n15900) | (n15785 & n15901) | (n15900 & n15901);
  assign n15903 = n5430 | n5432;
  assign n15904 = (n5430 & n15868) | (n5430 & n15903) | (n15868 & n15903);
  assign n15905 = (n5430 & n12488) | (n5430 & n15903) | (n12488 & n15903);
  assign n15906 = (n12383 & n15904) | (n12383 & n15905) | (n15904 & n15905);
  assign n15907 = (n12384 & n15904) | (n12384 & n15905) | (n15904 & n15905);
  assign n15908 = (n15760 & n15906) | (n15760 & n15907) | (n15906 & n15907);
  assign n5570 = x68 & x80;
  assign n5571 = x67 & x81;
  assign n5572 = n5570 & n5571;
  assign n5573 = n5570 | n5571;
  assign n5574 = ~n5572 & n5573;
  assign n15909 = n5423 | n5425;
  assign n15911 = n5574 & n15909;
  assign n15912 = n5423 & n5574;
  assign n15913 = (n15865 & n15911) | (n15865 & n15912) | (n15911 & n15912);
  assign n15915 = (n15866 & n15911) | (n15866 & n15912) | (n15911 & n15912);
  assign n12561 = (n15794 & n15913) | (n15794 & n15915) | (n15913 & n15915);
  assign n15916 = n5574 | n15909;
  assign n15917 = n5423 | n5574;
  assign n15918 = (n15865 & n15916) | (n15865 & n15917) | (n15916 & n15917);
  assign n15919 = (n15866 & n15916) | (n15866 & n15917) | (n15916 & n15917);
  assign n12564 = (n15794 & n15918) | (n15794 & n15919) | (n15918 & n15919);
  assign n5577 = ~n12561 & n12564;
  assign n5578 = x66 & x82;
  assign n5579 = n5577 & n5578;
  assign n5580 = n5577 | n5578;
  assign n5581 = ~n5579 & n5580;
  assign n5582 = n15908 & n5581;
  assign n5583 = n15908 | n5581;
  assign n5584 = ~n5582 & n5583;
  assign n5585 = x65 & x83;
  assign n5586 = n5584 & n5585;
  assign n5587 = n5584 | n5585;
  assign n5588 = ~n5586 & n5587;
  assign n5589 = n15902 & n5588;
  assign n5590 = n15902 | n5588;
  assign n5591 = ~n5589 & n5590;
  assign n5592 = x64 & x84;
  assign n5593 = n5591 & n5592;
  assign n5594 = n5591 | n5592;
  assign n5595 = ~n5593 & n5594;
  assign n12565 = n5444 & n5595;
  assign n15920 = (n5595 & n12511) | (n5595 & n12565) | (n12511 & n12565);
  assign n15921 = (n5595 & n12512) | (n5595 & n12565) | (n12512 & n12565);
  assign n15922 = (n15830 & n15920) | (n15830 & n15921) | (n15920 & n15921);
  assign n12567 = n5444 | n5595;
  assign n15923 = n12511 | n12567;
  assign n15924 = n12512 | n12567;
  assign n15925 = (n15830 & n15923) | (n15830 & n15924) | (n15923 & n15924);
  assign n5598 = ~n15922 & n15925;
  assign n5599 = x63 & x85;
  assign n5600 = n5598 & n5599;
  assign n5601 = n5598 | n5599;
  assign n5602 = ~n5600 & n5601;
  assign n5603 = n15895 & n5602;
  assign n5604 = n15895 | n5602;
  assign n5605 = ~n5603 & n5604;
  assign n5606 = x62 & x86;
  assign n5607 = n5605 & n5606;
  assign n5608 = n5605 | n5606;
  assign n5609 = ~n5607 & n5608;
  assign n12545 = n5458 | n5460;
  assign n12569 = n5609 & n12545;
  assign n12570 = n5458 & n5609;
  assign n12571 = (n15863 & n12569) | (n15863 & n12570) | (n12569 & n12570);
  assign n12572 = n5609 | n12545;
  assign n12573 = n5458 | n5609;
  assign n12574 = (n15863 & n12572) | (n15863 & n12573) | (n12572 & n12573);
  assign n5612 = ~n12571 & n12574;
  assign n5613 = x61 & x87;
  assign n5614 = n5612 & n5613;
  assign n5615 = n5612 | n5613;
  assign n5616 = ~n5614 & n5615;
  assign n12575 = n5465 & n5616;
  assign n15926 = (n5616 & n12521) | (n5616 & n12575) | (n12521 & n12575);
  assign n15927 = (n5467 & n5616) | (n5467 & n12575) | (n5616 & n12575);
  assign n15928 = (n12461 & n15926) | (n12461 & n15927) | (n15926 & n15927);
  assign n12577 = n5465 | n5616;
  assign n15929 = n12521 | n12577;
  assign n15930 = n5467 | n12577;
  assign n15931 = (n12461 & n15929) | (n12461 & n15930) | (n15929 & n15930);
  assign n5619 = ~n15928 & n15931;
  assign n5620 = x60 & x88;
  assign n5621 = n5619 & n5620;
  assign n5622 = n5619 | n5620;
  assign n5623 = ~n5621 & n5622;
  assign n12579 = n5472 & n5623;
  assign n12580 = (n5623 & n12526) | (n5623 & n12579) | (n12526 & n12579);
  assign n12581 = n5472 | n5623;
  assign n12582 = n12526 | n12581;
  assign n5626 = ~n12580 & n12582;
  assign n5627 = x59 & x89;
  assign n5628 = n5626 & n5627;
  assign n5629 = n5626 | n5627;
  assign n5630 = ~n5628 & n5629;
  assign n12583 = n5479 & n5630;
  assign n12584 = (n5630 & n12530) | (n5630 & n12583) | (n12530 & n12583);
  assign n12585 = n5479 | n5630;
  assign n12586 = n12530 | n12585;
  assign n5633 = ~n12584 & n12586;
  assign n5634 = x58 & x90;
  assign n5635 = n5633 & n5634;
  assign n5636 = n5633 | n5634;
  assign n5637 = ~n5635 & n5636;
  assign n5638 = n12544 & n5637;
  assign n5639 = n12544 | n5637;
  assign n5640 = ~n5638 & n5639;
  assign n5641 = x57 & x91;
  assign n5642 = n5640 & n5641;
  assign n5643 = n5640 | n5641;
  assign n5644 = ~n5642 & n5643;
  assign n5645 = n12542 & n5644;
  assign n5646 = n12542 | n5644;
  assign n5647 = ~n5645 & n5646;
  assign n5648 = x56 & x92;
  assign n5649 = n5647 & n5648;
  assign n5650 = n5647 | n5648;
  assign n5651 = ~n5649 & n5650;
  assign n5652 = n12540 & n5651;
  assign n5653 = n12540 | n5651;
  assign n5654 = ~n5652 & n5653;
  assign n5655 = x55 & x93;
  assign n5656 = n5654 & n5655;
  assign n5657 = n5654 | n5655;
  assign n5658 = ~n5656 & n5657;
  assign n5659 = n12538 & n5658;
  assign n5660 = n12538 | n5658;
  assign n5661 = ~n5659 & n5660;
  assign n5662 = x54 & x94;
  assign n5663 = n5661 & n5662;
  assign n5664 = n5661 | n5662;
  assign n5665 = ~n5663 & n5664;
  assign n5666 = n5556 & n5665;
  assign n5667 = n5556 | n5665;
  assign n5668 = ~n5666 & n5667;
  assign n5669 = x53 & x95;
  assign n5670 = n5668 & n5669;
  assign n5671 = n5668 | n5669;
  assign n5672 = ~n5670 & n5671;
  assign n5673 = n5555 & n5672;
  assign n5674 = n5555 | n5672;
  assign n5675 = ~n5673 & n5674;
  assign n5676 = x52 & x96;
  assign n5677 = n5675 & n5676;
  assign n5678 = n5675 | n5676;
  assign n5679 = ~n5677 & n5678;
  assign n5680 = n15890 & n5679;
  assign n5681 = n15890 | n5679;
  assign n5682 = ~n5680 & n5681;
  assign n5683 = x51 & x97;
  assign n5684 = n5682 & n5683;
  assign n5685 = n5682 | n5683;
  assign n5686 = ~n5684 & n5685;
  assign n5687 = n12536 & n5686;
  assign n5688 = n12536 | n5686;
  assign n5689 = ~n5687 & n5688;
  assign n5690 = x50 & x98;
  assign n5691 = n5689 & n5690;
  assign n5692 = n5689 | n5690;
  assign n5693 = ~n5691 & n5692;
  assign n5694 = n12534 & n5693;
  assign n5695 = n12534 | n5693;
  assign n5696 = ~n5694 & n5695;
  assign n5697 = x49 & x99;
  assign n5698 = n5696 & n5697;
  assign n5699 = n5696 | n5697;
  assign n5700 = ~n5698 & n5699;
  assign n5701 = n5549 & n5700;
  assign n5702 = n5549 | n5700;
  assign n5703 = ~n5701 & n5702;
  assign n5704 = x48 & x100;
  assign n5705 = n5703 & n5704;
  assign n5706 = n5703 | n5704;
  assign n5707 = ~n5705 & n5706;
  assign n17700 = n5548 | n5697;
  assign n17701 = (n5547 & n5697) | (n5547 & n17700) | (n5697 & n17700);
  assign n15933 = (n5549 & n5696) | (n5549 & n17701) | (n5696 & n17701);
  assign n12588 = (n5698 & n5700) | (n5698 & n15933) | (n5700 & n15933);
  assign n12589 = n5691 | n12534;
  assign n12590 = (n5691 & n5693) | (n5691 & n12589) | (n5693 & n12589);
  assign n12591 = n5684 | n12536;
  assign n12592 = (n5684 & n5686) | (n5684 & n12591) | (n5686 & n12591);
  assign n15934 = n5677 | n15890;
  assign n15935 = (n5677 & n5679) | (n5677 & n15934) | (n5679 & n15934);
  assign n5712 = n5670 | n5673;
  assign n12593 = n5663 | n5665;
  assign n12594 = (n5556 & n5663) | (n5556 & n12593) | (n5663 & n12593);
  assign n12595 = n5656 | n5658;
  assign n12596 = (n5656 & n12538) | (n5656 & n12595) | (n12538 & n12595);
  assign n12597 = n5649 | n5651;
  assign n12598 = (n5649 & n12540) | (n5649 & n12597) | (n12540 & n12597);
  assign n12599 = n5642 | n5644;
  assign n12600 = (n5642 & n12542) | (n5642 & n12599) | (n12542 & n12599);
  assign n12601 = n5635 | n5637;
  assign n12602 = (n5635 & n12544) | (n5635 & n12601) | (n12544 & n12601);
  assign n12604 = n5614 | n5616;
  assign n15936 = n5465 | n5614;
  assign n15937 = (n5614 & n5616) | (n5614 & n15936) | (n5616 & n15936);
  assign n15938 = (n12521 & n12604) | (n12521 & n15937) | (n12604 & n15937);
  assign n15939 = (n5467 & n12604) | (n5467 & n15937) | (n12604 & n15937);
  assign n15940 = (n12461 & n15938) | (n12461 & n15939) | (n15938 & n15939);
  assign n12609 = n5593 | n5595;
  assign n15941 = n5444 | n5593;
  assign n15942 = (n5593 & n5595) | (n5593 & n15941) | (n5595 & n15941);
  assign n15943 = (n12511 & n12609) | (n12511 & n15942) | (n12609 & n15942);
  assign n15944 = (n12512 & n12609) | (n12512 & n15942) | (n12609 & n15942);
  assign n15945 = (n15830 & n15943) | (n15830 & n15944) | (n15943 & n15944);
  assign n5727 = x69 & x80;
  assign n5728 = x68 & x81;
  assign n5729 = n5727 & n5728;
  assign n5730 = n5727 | n5728;
  assign n5731 = ~n5729 & n5730;
  assign n12615 = n5572 & n5731;
  assign n15946 = (n5731 & n12615) | (n5731 & n15915) | (n12615 & n15915);
  assign n15947 = (n5731 & n12615) | (n5731 & n15913) | (n12615 & n15913);
  assign n15948 = (n15794 & n15946) | (n15794 & n15947) | (n15946 & n15947);
  assign n12617 = n5572 | n5731;
  assign n15949 = n12617 | n15915;
  assign n15950 = n12617 | n15913;
  assign n15951 = (n15794 & n15949) | (n15794 & n15950) | (n15949 & n15950);
  assign n5734 = ~n15948 & n15951;
  assign n5735 = x67 & x82;
  assign n5736 = n5734 & n5735;
  assign n5737 = n5734 | n5735;
  assign n5738 = ~n5736 & n5737;
  assign n12613 = n5579 | n5581;
  assign n12619 = n5738 & n12613;
  assign n12620 = n5579 & n5738;
  assign n12621 = (n15908 & n12619) | (n15908 & n12620) | (n12619 & n12620);
  assign n12622 = n5738 | n12613;
  assign n12623 = n5579 | n5738;
  assign n12624 = (n15908 & n12622) | (n15908 & n12623) | (n12622 & n12623);
  assign n5741 = ~n12621 & n12624;
  assign n5742 = x66 & x83;
  assign n5743 = n5741 & n5742;
  assign n5744 = n5741 | n5742;
  assign n5745 = ~n5743 & n5744;
  assign n12611 = n5586 | n5588;
  assign n12625 = n5745 & n12611;
  assign n12626 = n5586 & n5745;
  assign n12627 = (n15902 & n12625) | (n15902 & n12626) | (n12625 & n12626);
  assign n12628 = n5745 | n12611;
  assign n12629 = n5586 | n5745;
  assign n12630 = (n15902 & n12628) | (n15902 & n12629) | (n12628 & n12629);
  assign n5748 = ~n12627 & n12630;
  assign n5749 = x65 & x84;
  assign n5750 = n5748 & n5749;
  assign n5751 = n5748 | n5749;
  assign n5752 = ~n5750 & n5751;
  assign n5753 = n15945 & n5752;
  assign n5754 = n15945 | n5752;
  assign n5755 = ~n5753 & n5754;
  assign n5756 = x64 & x85;
  assign n5757 = n5755 & n5756;
  assign n5758 = n5755 | n5756;
  assign n5759 = ~n5757 & n5758;
  assign n12606 = n5600 | n5602;
  assign n12631 = n5759 & n12606;
  assign n12632 = n5600 & n5759;
  assign n12633 = (n15895 & n12631) | (n15895 & n12632) | (n12631 & n12632);
  assign n12634 = n5759 | n12606;
  assign n12635 = n5600 | n5759;
  assign n12636 = (n15895 & n12634) | (n15895 & n12635) | (n12634 & n12635);
  assign n5762 = ~n12633 & n12636;
  assign n5763 = x63 & x86;
  assign n5764 = n5762 & n5763;
  assign n5765 = n5762 | n5763;
  assign n5766 = ~n5764 & n5765;
  assign n12637 = n5607 & n5766;
  assign n15952 = (n5766 & n12570) | (n5766 & n12637) | (n12570 & n12637);
  assign n15953 = (n5766 & n12569) | (n5766 & n12637) | (n12569 & n12637);
  assign n15954 = (n15863 & n15952) | (n15863 & n15953) | (n15952 & n15953);
  assign n12639 = n5607 | n5766;
  assign n15955 = n12570 | n12639;
  assign n15956 = n12569 | n12639;
  assign n15957 = (n15863 & n15955) | (n15863 & n15956) | (n15955 & n15956);
  assign n5769 = ~n15954 & n15957;
  assign n5770 = x62 & x87;
  assign n5771 = n5769 & n5770;
  assign n5772 = n5769 | n5770;
  assign n5773 = ~n5771 & n5772;
  assign n5774 = n15940 & n5773;
  assign n5775 = n15940 | n5773;
  assign n5776 = ~n5774 & n5775;
  assign n5777 = x61 & x88;
  assign n5778 = n5776 & n5777;
  assign n5779 = n5776 | n5777;
  assign n5780 = ~n5778 & n5779;
  assign n12641 = n5621 & n5780;
  assign n12642 = (n5780 & n12580) | (n5780 & n12641) | (n12580 & n12641);
  assign n12643 = n5621 | n5780;
  assign n12644 = n12580 | n12643;
  assign n5783 = ~n12642 & n12644;
  assign n5784 = x60 & x89;
  assign n5785 = n5783 & n5784;
  assign n5786 = n5783 | n5784;
  assign n5787 = ~n5785 & n5786;
  assign n12645 = n5628 & n5787;
  assign n12646 = (n5787 & n12584) | (n5787 & n12645) | (n12584 & n12645);
  assign n12647 = n5628 | n5787;
  assign n12648 = n12584 | n12647;
  assign n5790 = ~n12646 & n12648;
  assign n5791 = x59 & x90;
  assign n5792 = n5790 & n5791;
  assign n5793 = n5790 | n5791;
  assign n5794 = ~n5792 & n5793;
  assign n5795 = n12602 & n5794;
  assign n5796 = n12602 | n5794;
  assign n5797 = ~n5795 & n5796;
  assign n5798 = x58 & x91;
  assign n5799 = n5797 & n5798;
  assign n5800 = n5797 | n5798;
  assign n5801 = ~n5799 & n5800;
  assign n5802 = n12600 & n5801;
  assign n5803 = n12600 | n5801;
  assign n5804 = ~n5802 & n5803;
  assign n5805 = x57 & x92;
  assign n5806 = n5804 & n5805;
  assign n5807 = n5804 | n5805;
  assign n5808 = ~n5806 & n5807;
  assign n5809 = n12598 & n5808;
  assign n5810 = n12598 | n5808;
  assign n5811 = ~n5809 & n5810;
  assign n5812 = x56 & x93;
  assign n5813 = n5811 & n5812;
  assign n5814 = n5811 | n5812;
  assign n5815 = ~n5813 & n5814;
  assign n5816 = n12596 & n5815;
  assign n5817 = n12596 | n5815;
  assign n5818 = ~n5816 & n5817;
  assign n5819 = x55 & x94;
  assign n5820 = n5818 & n5819;
  assign n5821 = n5818 | n5819;
  assign n5822 = ~n5820 & n5821;
  assign n5823 = n12594 & n5822;
  assign n5824 = n12594 | n5822;
  assign n5825 = ~n5823 & n5824;
  assign n5826 = x54 & x95;
  assign n5827 = n5825 & n5826;
  assign n5828 = n5825 | n5826;
  assign n5829 = ~n5827 & n5828;
  assign n5830 = n5712 & n5829;
  assign n5831 = n5712 | n5829;
  assign n5832 = ~n5830 & n5831;
  assign n5833 = x53 & x96;
  assign n5834 = n5832 & n5833;
  assign n5835 = n5832 | n5833;
  assign n5836 = ~n5834 & n5835;
  assign n5837 = n15935 & n5836;
  assign n5838 = n15935 | n5836;
  assign n5839 = ~n5837 & n5838;
  assign n5840 = x52 & x97;
  assign n5841 = n5839 & n5840;
  assign n5842 = n5839 | n5840;
  assign n5843 = ~n5841 & n5842;
  assign n5844 = n12592 & n5843;
  assign n5845 = n12592 | n5843;
  assign n5846 = ~n5844 & n5845;
  assign n5847 = x51 & x98;
  assign n5848 = n5846 & n5847;
  assign n5849 = n5846 | n5847;
  assign n5850 = ~n5848 & n5849;
  assign n5851 = n12590 & n5850;
  assign n5852 = n12590 | n5850;
  assign n5853 = ~n5851 & n5852;
  assign n5854 = x50 & x99;
  assign n5855 = n5853 & n5854;
  assign n5856 = n5853 | n5854;
  assign n5857 = ~n5855 & n5856;
  assign n5858 = n12588 & n5857;
  assign n5859 = n12588 | n5857;
  assign n5860 = ~n5858 & n5859;
  assign n5861 = x49 & x100;
  assign n5862 = n5860 & n5861;
  assign n5863 = n5860 | n5861;
  assign n5864 = ~n5862 & n5863;
  assign n5865 = n5705 & n5864;
  assign n5866 = n5705 | n5864;
  assign n5867 = ~n5865 & n5866;
  assign n5868 = x48 & x101;
  assign n5869 = n5867 & n5868;
  assign n5870 = n5867 | n5868;
  assign n5871 = ~n5869 & n5870;
  assign n17702 = n5704 | n5861;
  assign n17703 = (n5703 & n5861) | (n5703 & n17702) | (n5861 & n17702);
  assign n15959 = (n5705 & n5860) | (n5705 & n17703) | (n5860 & n17703);
  assign n12650 = (n5862 & n5864) | (n5862 & n15959) | (n5864 & n15959);
  assign n12651 = n5855 | n12588;
  assign n12652 = (n5855 & n5857) | (n5855 & n12651) | (n5857 & n12651);
  assign n12653 = n5848 | n12590;
  assign n12654 = (n5848 & n5850) | (n5848 & n12653) | (n5850 & n12653);
  assign n12655 = n5841 | n12592;
  assign n12656 = (n5841 & n5843) | (n5841 & n12655) | (n5843 & n12655);
  assign n15960 = n5834 | n15935;
  assign n15961 = (n5834 & n5836) | (n5834 & n15960) | (n5836 & n15960);
  assign n12657 = n5827 | n5829;
  assign n12658 = (n5712 & n5827) | (n5712 & n12657) | (n5827 & n12657);
  assign n12659 = n5820 | n5822;
  assign n12660 = (n5820 & n12594) | (n5820 & n12659) | (n12594 & n12659);
  assign n12661 = n5813 | n5815;
  assign n12662 = (n5813 & n12596) | (n5813 & n12661) | (n12596 & n12661);
  assign n12663 = n5806 | n5808;
  assign n12664 = (n5806 & n12598) | (n5806 & n12663) | (n12598 & n12663);
  assign n12665 = n5799 | n5801;
  assign n12666 = (n5799 & n12600) | (n5799 & n12665) | (n12600 & n12665);
  assign n12667 = n5792 | n5794;
  assign n12668 = (n5792 & n12602) | (n5792 & n12667) | (n12602 & n12667);
  assign n12672 = n5764 | n5766;
  assign n15962 = n5607 | n5764;
  assign n15963 = (n5764 & n5766) | (n5764 & n15962) | (n5766 & n15962);
  assign n15964 = (n12570 & n12672) | (n12570 & n15963) | (n12672 & n15963);
  assign n15965 = (n12569 & n12672) | (n12569 & n15963) | (n12672 & n15963);
  assign n15966 = (n15863 & n15964) | (n15863 & n15965) | (n15964 & n15965);
  assign n5892 = x70 & x80;
  assign n5893 = x69 & x81;
  assign n5894 = n5892 & n5893;
  assign n5895 = n5892 | n5893;
  assign n5896 = ~n5894 & n5895;
  assign n15971 = n5572 | n5729;
  assign n15972 = (n5729 & n5731) | (n5729 & n15971) | (n5731 & n15971);
  assign n12685 = n5896 & n15972;
  assign n12683 = n5729 | n5731;
  assign n12686 = n5896 & n12683;
  assign n15973 = (n12685 & n12686) | (n12685 & n15915) | (n12686 & n15915);
  assign n15974 = (n12685 & n12686) | (n12685 & n15913) | (n12686 & n15913);
  assign n15975 = (n15794 & n15973) | (n15794 & n15974) | (n15973 & n15974);
  assign n12688 = n5896 | n15972;
  assign n12689 = n5896 | n12683;
  assign n15976 = (n12688 & n12689) | (n12688 & n15915) | (n12689 & n15915);
  assign n15977 = (n12688 & n12689) | (n12688 & n15913) | (n12689 & n15913);
  assign n15978 = (n15794 & n15976) | (n15794 & n15977) | (n15976 & n15977);
  assign n5899 = ~n15975 & n15978;
  assign n5900 = x68 & x82;
  assign n5901 = n5899 & n5900;
  assign n5902 = n5899 | n5900;
  assign n5903 = ~n5901 & n5902;
  assign n15979 = n5736 | n5738;
  assign n15980 = (n5736 & n12613) | (n5736 & n15979) | (n12613 & n15979);
  assign n12691 = n5903 & n15980;
  assign n15981 = n5579 | n5736;
  assign n15982 = (n5736 & n5738) | (n5736 & n15981) | (n5738 & n15981);
  assign n12692 = n5903 & n15982;
  assign n12693 = (n15908 & n12691) | (n15908 & n12692) | (n12691 & n12692);
  assign n12694 = n5903 | n15980;
  assign n12695 = n5903 | n15982;
  assign n12696 = (n15908 & n12694) | (n15908 & n12695) | (n12694 & n12695);
  assign n5906 = ~n12693 & n12696;
  assign n5907 = x67 & x83;
  assign n5908 = n5906 & n5907;
  assign n5909 = n5906 | n5907;
  assign n5910 = ~n5908 & n5909;
  assign n15967 = n5743 | n5745;
  assign n15968 = (n5743 & n12611) | (n5743 & n15967) | (n12611 & n15967);
  assign n15983 = n5910 & n15968;
  assign n15969 = n5586 | n5743;
  assign n15970 = (n5743 & n5745) | (n5743 & n15969) | (n5745 & n15969);
  assign n15984 = n5910 & n15970;
  assign n15985 = (n15902 & n15983) | (n15902 & n15984) | (n15983 & n15984);
  assign n15986 = n5910 | n15968;
  assign n15987 = n5910 | n15970;
  assign n15988 = (n15902 & n15986) | (n15902 & n15987) | (n15986 & n15987);
  assign n5913 = ~n15985 & n15988;
  assign n5914 = x66 & x84;
  assign n5915 = n5913 & n5914;
  assign n5916 = n5913 | n5914;
  assign n5917 = ~n5915 & n5916;
  assign n12674 = n5750 | n5752;
  assign n12697 = n5917 & n12674;
  assign n12698 = n5750 & n5917;
  assign n12699 = (n15945 & n12697) | (n15945 & n12698) | (n12697 & n12698);
  assign n12700 = n5917 | n12674;
  assign n12701 = n5750 | n5917;
  assign n12702 = (n15945 & n12700) | (n15945 & n12701) | (n12700 & n12701);
  assign n5920 = ~n12699 & n12702;
  assign n5921 = x65 & x85;
  assign n5922 = n5920 & n5921;
  assign n5923 = n5920 | n5921;
  assign n5924 = ~n5922 & n5923;
  assign n12703 = n5757 & n5924;
  assign n15989 = (n5924 & n12632) | (n5924 & n12703) | (n12632 & n12703);
  assign n15990 = (n5924 & n12631) | (n5924 & n12703) | (n12631 & n12703);
  assign n15991 = (n15895 & n15989) | (n15895 & n15990) | (n15989 & n15990);
  assign n12705 = n5757 | n5924;
  assign n15992 = n12632 | n12705;
  assign n15993 = n12631 | n12705;
  assign n15994 = (n15895 & n15992) | (n15895 & n15993) | (n15992 & n15993);
  assign n5927 = ~n15991 & n15994;
  assign n5928 = x64 & x86;
  assign n5929 = n5927 & n5928;
  assign n5930 = n5927 | n5928;
  assign n5931 = ~n5929 & n5930;
  assign n5932 = n15966 & n5931;
  assign n5933 = n15966 | n5931;
  assign n5934 = ~n5932 & n5933;
  assign n5935 = x63 & x87;
  assign n5936 = n5934 & n5935;
  assign n5937 = n5934 | n5935;
  assign n5938 = ~n5936 & n5937;
  assign n12669 = n5771 | n5773;
  assign n12707 = n5938 & n12669;
  assign n12708 = n5771 & n5938;
  assign n12709 = (n15940 & n12707) | (n15940 & n12708) | (n12707 & n12708);
  assign n12710 = n5938 | n12669;
  assign n12711 = n5771 | n5938;
  assign n12712 = (n15940 & n12710) | (n15940 & n12711) | (n12710 & n12711);
  assign n5941 = ~n12709 & n12712;
  assign n5942 = x62 & x88;
  assign n5943 = n5941 & n5942;
  assign n5944 = n5941 | n5942;
  assign n5945 = ~n5943 & n5944;
  assign n12713 = n5778 & n5945;
  assign n15995 = (n5945 & n12641) | (n5945 & n12713) | (n12641 & n12713);
  assign n15996 = (n5780 & n5945) | (n5780 & n12713) | (n5945 & n12713);
  assign n15997 = (n12580 & n15995) | (n12580 & n15996) | (n15995 & n15996);
  assign n12715 = n5778 | n5945;
  assign n15998 = n12641 | n12715;
  assign n15999 = n5780 | n12715;
  assign n16000 = (n12580 & n15998) | (n12580 & n15999) | (n15998 & n15999);
  assign n5948 = ~n15997 & n16000;
  assign n5949 = x61 & x89;
  assign n5950 = n5948 & n5949;
  assign n5951 = n5948 | n5949;
  assign n5952 = ~n5950 & n5951;
  assign n12717 = n5785 & n5952;
  assign n12718 = (n5952 & n12646) | (n5952 & n12717) | (n12646 & n12717);
  assign n12719 = n5785 | n5952;
  assign n12720 = n12646 | n12719;
  assign n5955 = ~n12718 & n12720;
  assign n5956 = x60 & x90;
  assign n5957 = n5955 & n5956;
  assign n5958 = n5955 | n5956;
  assign n5959 = ~n5957 & n5958;
  assign n5960 = n12668 & n5959;
  assign n5961 = n12668 | n5959;
  assign n5962 = ~n5960 & n5961;
  assign n5963 = x59 & x91;
  assign n5964 = n5962 & n5963;
  assign n5965 = n5962 | n5963;
  assign n5966 = ~n5964 & n5965;
  assign n5967 = n12666 & n5966;
  assign n5968 = n12666 | n5966;
  assign n5969 = ~n5967 & n5968;
  assign n5970 = x58 & x92;
  assign n5971 = n5969 & n5970;
  assign n5972 = n5969 | n5970;
  assign n5973 = ~n5971 & n5972;
  assign n5974 = n12664 & n5973;
  assign n5975 = n12664 | n5973;
  assign n5976 = ~n5974 & n5975;
  assign n5977 = x57 & x93;
  assign n5978 = n5976 & n5977;
  assign n5979 = n5976 | n5977;
  assign n5980 = ~n5978 & n5979;
  assign n5981 = n12662 & n5980;
  assign n5982 = n12662 | n5980;
  assign n5983 = ~n5981 & n5982;
  assign n5984 = x56 & x94;
  assign n5985 = n5983 & n5984;
  assign n5986 = n5983 | n5984;
  assign n5987 = ~n5985 & n5986;
  assign n5988 = n12660 & n5987;
  assign n5989 = n12660 | n5987;
  assign n5990 = ~n5988 & n5989;
  assign n5991 = x55 & x95;
  assign n5992 = n5990 & n5991;
  assign n5993 = n5990 | n5991;
  assign n5994 = ~n5992 & n5993;
  assign n5995 = n12658 & n5994;
  assign n5996 = n12658 | n5994;
  assign n5997 = ~n5995 & n5996;
  assign n5998 = x54 & x96;
  assign n5999 = n5997 & n5998;
  assign n6000 = n5997 | n5998;
  assign n6001 = ~n5999 & n6000;
  assign n6002 = n15961 & n6001;
  assign n6003 = n15961 | n6001;
  assign n6004 = ~n6002 & n6003;
  assign n6005 = x53 & x97;
  assign n6006 = n6004 & n6005;
  assign n6007 = n6004 | n6005;
  assign n6008 = ~n6006 & n6007;
  assign n6009 = n12656 & n6008;
  assign n6010 = n12656 | n6008;
  assign n6011 = ~n6009 & n6010;
  assign n6012 = x52 & x98;
  assign n6013 = n6011 & n6012;
  assign n6014 = n6011 | n6012;
  assign n6015 = ~n6013 & n6014;
  assign n6016 = n12654 & n6015;
  assign n6017 = n12654 | n6015;
  assign n6018 = ~n6016 & n6017;
  assign n6019 = x51 & x99;
  assign n6020 = n6018 & n6019;
  assign n6021 = n6018 | n6019;
  assign n6022 = ~n6020 & n6021;
  assign n6023 = n12652 & n6022;
  assign n6024 = n12652 | n6022;
  assign n6025 = ~n6023 & n6024;
  assign n6026 = x50 & x100;
  assign n6027 = n6025 & n6026;
  assign n6028 = n6025 | n6026;
  assign n6029 = ~n6027 & n6028;
  assign n6030 = n12650 & n6029;
  assign n6031 = n12650 | n6029;
  assign n6032 = ~n6030 & n6031;
  assign n6033 = x49 & x101;
  assign n6034 = n6032 & n6033;
  assign n6035 = n6032 | n6033;
  assign n6036 = ~n6034 & n6035;
  assign n6037 = n5869 & n6036;
  assign n6038 = n5869 | n6036;
  assign n6039 = ~n6037 & n6038;
  assign n6040 = x48 & x102;
  assign n6041 = n6039 & n6040;
  assign n6042 = n6039 | n6040;
  assign n6043 = ~n6041 & n6042;
  assign n12721 = n5869 | n6034;
  assign n12722 = (n6034 & n6036) | (n6034 & n12721) | (n6036 & n12721);
  assign n12723 = n6027 | n12650;
  assign n12724 = (n6027 & n6029) | (n6027 & n12723) | (n6029 & n12723);
  assign n12725 = n6020 | n12652;
  assign n12726 = (n6020 & n6022) | (n6020 & n12725) | (n6022 & n12725);
  assign n12727 = n6013 | n12654;
  assign n12728 = (n6013 & n6015) | (n6013 & n12727) | (n6015 & n12727);
  assign n12729 = n6006 | n12656;
  assign n12730 = (n6006 & n6008) | (n6006 & n12729) | (n6008 & n12729);
  assign n12731 = n5999 | n6001;
  assign n12732 = (n15961 & n5999) | (n15961 & n12731) | (n5999 & n12731);
  assign n12733 = n5992 | n5994;
  assign n12734 = (n5992 & n12658) | (n5992 & n12733) | (n12658 & n12733);
  assign n12735 = n5985 | n5987;
  assign n12736 = (n5985 & n12660) | (n5985 & n12735) | (n12660 & n12735);
  assign n12737 = n5978 | n5980;
  assign n12738 = (n5978 & n12662) | (n5978 & n12737) | (n12662 & n12737);
  assign n12739 = n5971 | n5973;
  assign n12740 = (n5971 & n12664) | (n5971 & n12739) | (n12664 & n12739);
  assign n12741 = n5964 | n5966;
  assign n12742 = (n5964 & n12666) | (n5964 & n12741) | (n12666 & n12741);
  assign n12743 = n5957 | n5959;
  assign n12744 = (n5957 & n12668) | (n5957 & n12743) | (n12668 & n12743);
  assign n12746 = n5943 | n5945;
  assign n16001 = n5778 | n5943;
  assign n16002 = (n5943 & n5945) | (n5943 & n16001) | (n5945 & n16001);
  assign n16003 = (n12641 & n12746) | (n12641 & n16002) | (n12746 & n16002);
  assign n16004 = (n5780 & n12746) | (n5780 & n16002) | (n12746 & n16002);
  assign n16005 = (n12580 & n16003) | (n12580 & n16004) | (n16003 & n16004);
  assign n12751 = n5922 | n5924;
  assign n16006 = n5757 | n5922;
  assign n16007 = (n5922 & n5924) | (n5922 & n16006) | (n5924 & n16006);
  assign n16008 = (n12632 & n12751) | (n12632 & n16007) | (n12751 & n16007);
  assign n16009 = (n12631 & n12751) | (n12631 & n16007) | (n12751 & n16007);
  assign n16010 = (n15895 & n16008) | (n15895 & n16009) | (n16008 & n16009);
  assign n6065 = x71 & x80;
  assign n6066 = x70 & x81;
  assign n6067 = n6065 & n6066;
  assign n6068 = n6065 | n6066;
  assign n6069 = ~n6067 & n6068;
  assign n16018 = n5894 | n5896;
  assign n16019 = (n5894 & n15972) | (n5894 & n16018) | (n15972 & n16018);
  assign n12764 = n6069 & n16019;
  assign n16020 = (n5894 & n12683) | (n5894 & n16018) | (n12683 & n16018);
  assign n12765 = n6069 & n16020;
  assign n16021 = (n12764 & n12765) | (n12764 & n15915) | (n12765 & n15915);
  assign n16022 = (n12764 & n12765) | (n12764 & n15913) | (n12765 & n15913);
  assign n16023 = (n15794 & n16021) | (n15794 & n16022) | (n16021 & n16022);
  assign n12767 = n6069 | n16019;
  assign n12768 = n6069 | n16020;
  assign n16024 = (n12767 & n12768) | (n12767 & n15915) | (n12768 & n15915);
  assign n16025 = (n12767 & n12768) | (n12767 & n15913) | (n12768 & n15913);
  assign n16026 = (n15794 & n16024) | (n15794 & n16025) | (n16024 & n16025);
  assign n6072 = ~n16023 & n16026;
  assign n6073 = x69 & x82;
  assign n6074 = n6072 & n6073;
  assign n6075 = n6072 | n6073;
  assign n6076 = ~n6074 & n6075;
  assign n16015 = n5901 | n5903;
  assign n17704 = n6076 & n16015;
  assign n17705 = n5901 & n6076;
  assign n17706 = (n15980 & n17704) | (n15980 & n17705) | (n17704 & n17705);
  assign n16016 = (n5901 & n15982) | (n5901 & n16015) | (n15982 & n16015);
  assign n16028 = n6076 & n16016;
  assign n16029 = (n15908 & n17706) | (n15908 & n16028) | (n17706 & n16028);
  assign n17707 = n6076 | n16015;
  assign n17708 = n5901 | n6076;
  assign n17709 = (n15980 & n17707) | (n15980 & n17708) | (n17707 & n17708);
  assign n16031 = n6076 | n16016;
  assign n16032 = (n15908 & n17709) | (n15908 & n16031) | (n17709 & n16031);
  assign n6079 = ~n16029 & n16032;
  assign n6080 = x68 & x83;
  assign n6081 = n6079 & n6080;
  assign n6082 = n6079 | n6080;
  assign n6083 = ~n6081 & n6082;
  assign n12756 = n5908 | n5910;
  assign n12770 = n6083 & n12756;
  assign n12771 = n5908 & n6083;
  assign n16033 = (n12770 & n12771) | (n12770 & n15968) | (n12771 & n15968);
  assign n16034 = (n12770 & n12771) | (n12770 & n15970) | (n12771 & n15970);
  assign n16035 = (n15902 & n16033) | (n15902 & n16034) | (n16033 & n16034);
  assign n12773 = n6083 | n12756;
  assign n12774 = n5908 | n6083;
  assign n16036 = (n12773 & n12774) | (n12773 & n15968) | (n12774 & n15968);
  assign n16037 = (n12773 & n12774) | (n12773 & n15970) | (n12774 & n15970);
  assign n16038 = (n15902 & n16036) | (n15902 & n16037) | (n16036 & n16037);
  assign n6086 = ~n16035 & n16038;
  assign n6087 = x67 & x84;
  assign n6088 = n6086 & n6087;
  assign n6089 = n6086 | n6087;
  assign n6090 = ~n6088 & n6089;
  assign n16013 = n5915 | n5917;
  assign n16014 = (n5915 & n12674) | (n5915 & n16013) | (n12674 & n16013);
  assign n16039 = n6090 & n16014;
  assign n16011 = n5750 | n5915;
  assign n16012 = (n5915 & n5917) | (n5915 & n16011) | (n5917 & n16011);
  assign n16040 = n6090 & n16012;
  assign n16041 = (n15945 & n16039) | (n15945 & n16040) | (n16039 & n16040);
  assign n16042 = n6090 | n16014;
  assign n16043 = n6090 | n16012;
  assign n16044 = (n15945 & n16042) | (n15945 & n16043) | (n16042 & n16043);
  assign n6093 = ~n16041 & n16044;
  assign n6094 = x66 & x85;
  assign n6095 = n6093 & n6094;
  assign n6096 = n6093 | n6094;
  assign n6097 = ~n6095 & n6096;
  assign n6098 = n16010 & n6097;
  assign n6099 = n16010 | n6097;
  assign n6100 = ~n6098 & n6099;
  assign n6101 = x65 & x86;
  assign n6102 = n6100 & n6101;
  assign n6103 = n6100 | n6101;
  assign n6104 = ~n6102 & n6103;
  assign n12748 = n5929 | n5931;
  assign n12776 = n6104 & n12748;
  assign n12777 = n5929 & n6104;
  assign n12778 = (n15966 & n12776) | (n15966 & n12777) | (n12776 & n12777);
  assign n12779 = n6104 | n12748;
  assign n12780 = n5929 | n6104;
  assign n12781 = (n15966 & n12779) | (n15966 & n12780) | (n12779 & n12780);
  assign n6107 = ~n12778 & n12781;
  assign n6108 = x64 & x87;
  assign n6109 = n6107 & n6108;
  assign n6110 = n6107 | n6108;
  assign n6111 = ~n6109 & n6110;
  assign n12782 = n5936 & n6111;
  assign n16045 = (n6111 & n12708) | (n6111 & n12782) | (n12708 & n12782);
  assign n16046 = (n6111 & n12707) | (n6111 & n12782) | (n12707 & n12782);
  assign n16047 = (n15940 & n16045) | (n15940 & n16046) | (n16045 & n16046);
  assign n12784 = n5936 | n6111;
  assign n16048 = n12708 | n12784;
  assign n16049 = n12707 | n12784;
  assign n16050 = (n15940 & n16048) | (n15940 & n16049) | (n16048 & n16049);
  assign n6114 = ~n16047 & n16050;
  assign n6115 = x63 & x88;
  assign n6116 = n6114 & n6115;
  assign n6117 = n6114 | n6115;
  assign n6118 = ~n6116 & n6117;
  assign n6119 = n16005 & n6118;
  assign n6120 = n16005 | n6118;
  assign n6121 = ~n6119 & n6120;
  assign n6122 = x62 & x89;
  assign n6123 = n6121 & n6122;
  assign n6124 = n6121 | n6122;
  assign n6125 = ~n6123 & n6124;
  assign n12786 = n5950 & n6125;
  assign n12787 = (n6125 & n12718) | (n6125 & n12786) | (n12718 & n12786);
  assign n12788 = n5950 | n6125;
  assign n12789 = n12718 | n12788;
  assign n6128 = ~n12787 & n12789;
  assign n6129 = x61 & x90;
  assign n6130 = n6128 & n6129;
  assign n6131 = n6128 | n6129;
  assign n6132 = ~n6130 & n6131;
  assign n6133 = n12744 & n6132;
  assign n6134 = n12744 | n6132;
  assign n6135 = ~n6133 & n6134;
  assign n6136 = x60 & x91;
  assign n6137 = n6135 & n6136;
  assign n6138 = n6135 | n6136;
  assign n6139 = ~n6137 & n6138;
  assign n6140 = n12742 & n6139;
  assign n6141 = n12742 | n6139;
  assign n6142 = ~n6140 & n6141;
  assign n6143 = x59 & x92;
  assign n6144 = n6142 & n6143;
  assign n6145 = n6142 | n6143;
  assign n6146 = ~n6144 & n6145;
  assign n6147 = n12740 & n6146;
  assign n6148 = n12740 | n6146;
  assign n6149 = ~n6147 & n6148;
  assign n6150 = x58 & x93;
  assign n6151 = n6149 & n6150;
  assign n6152 = n6149 | n6150;
  assign n6153 = ~n6151 & n6152;
  assign n6154 = n12738 & n6153;
  assign n6155 = n12738 | n6153;
  assign n6156 = ~n6154 & n6155;
  assign n6157 = x57 & x94;
  assign n6158 = n6156 & n6157;
  assign n6159 = n6156 | n6157;
  assign n6160 = ~n6158 & n6159;
  assign n6161 = n12736 & n6160;
  assign n6162 = n12736 | n6160;
  assign n6163 = ~n6161 & n6162;
  assign n6164 = x56 & x95;
  assign n6165 = n6163 & n6164;
  assign n6166 = n6163 | n6164;
  assign n6167 = ~n6165 & n6166;
  assign n6168 = n12734 & n6167;
  assign n6169 = n12734 | n6167;
  assign n6170 = ~n6168 & n6169;
  assign n6171 = x55 & x96;
  assign n6172 = n6170 & n6171;
  assign n6173 = n6170 | n6171;
  assign n6174 = ~n6172 & n6173;
  assign n6175 = n12732 & n6174;
  assign n6176 = n12732 | n6174;
  assign n6177 = ~n6175 & n6176;
  assign n6178 = x54 & x97;
  assign n6179 = n6177 & n6178;
  assign n6180 = n6177 | n6178;
  assign n6181 = ~n6179 & n6180;
  assign n6182 = n12730 & n6181;
  assign n6183 = n12730 | n6181;
  assign n6184 = ~n6182 & n6183;
  assign n6185 = x53 & x98;
  assign n6186 = n6184 & n6185;
  assign n6187 = n6184 | n6185;
  assign n6188 = ~n6186 & n6187;
  assign n6189 = n12728 & n6188;
  assign n6190 = n12728 | n6188;
  assign n6191 = ~n6189 & n6190;
  assign n6192 = x52 & x99;
  assign n6193 = n6191 & n6192;
  assign n6194 = n6191 | n6192;
  assign n6195 = ~n6193 & n6194;
  assign n6196 = n12726 & n6195;
  assign n6197 = n12726 | n6195;
  assign n6198 = ~n6196 & n6197;
  assign n6199 = x51 & x100;
  assign n6200 = n6198 & n6199;
  assign n6201 = n6198 | n6199;
  assign n6202 = ~n6200 & n6201;
  assign n6203 = n12724 & n6202;
  assign n6204 = n12724 | n6202;
  assign n6205 = ~n6203 & n6204;
  assign n6206 = x50 & x101;
  assign n6207 = n6205 & n6206;
  assign n6208 = n6205 | n6206;
  assign n6209 = ~n6207 & n6208;
  assign n6210 = n12722 & n6209;
  assign n6211 = n12722 | n6209;
  assign n6212 = ~n6210 & n6211;
  assign n6213 = x49 & x102;
  assign n6214 = n6212 & n6213;
  assign n6215 = n6212 | n6213;
  assign n6216 = ~n6214 & n6215;
  assign n6217 = n6041 & n6216;
  assign n6218 = n6041 | n6216;
  assign n6219 = ~n6217 & n6218;
  assign n6220 = x48 & x103;
  assign n6221 = n6219 & n6220;
  assign n6222 = n6219 | n6220;
  assign n6223 = ~n6221 & n6222;
  assign n17710 = n6040 | n6213;
  assign n17711 = (n6039 & n6213) | (n6039 & n17710) | (n6213 & n17710);
  assign n16052 = (n6041 & n6212) | (n6041 & n17711) | (n6212 & n17711);
  assign n12791 = (n6214 & n6216) | (n6214 & n16052) | (n6216 & n16052);
  assign n16053 = n6207 | n12722;
  assign n16054 = (n6207 & n6209) | (n6207 & n16053) | (n6209 & n16053);
  assign n6226 = n6200 | n6203;
  assign n6227 = n6193 | n6196;
  assign n6228 = n6186 | n6189;
  assign n6229 = n6179 | n6182;
  assign n12792 = n6172 | n6174;
  assign n12793 = (n6172 & n12732) | (n6172 & n12792) | (n12732 & n12792);
  assign n12794 = n6165 | n6167;
  assign n12795 = (n6165 & n12734) | (n6165 & n12794) | (n12734 & n12794);
  assign n12796 = n6158 | n6160;
  assign n12797 = (n6158 & n12736) | (n6158 & n12796) | (n12736 & n12796);
  assign n12798 = n6151 | n6153;
  assign n12799 = (n6151 & n12738) | (n6151 & n12798) | (n12738 & n12798);
  assign n12800 = n6144 | n6146;
  assign n12801 = (n6144 & n12740) | (n6144 & n12800) | (n12740 & n12800);
  assign n12802 = n6137 | n6139;
  assign n12803 = (n6137 & n12742) | (n6137 & n12802) | (n12742 & n12802);
  assign n12804 = n6130 | n6132;
  assign n12805 = (n6130 & n12744) | (n6130 & n12804) | (n12744 & n12804);
  assign n12809 = n6109 | n6111;
  assign n16055 = n5936 | n6109;
  assign n16056 = (n6109 & n6111) | (n6109 & n16055) | (n6111 & n16055);
  assign n16057 = (n12708 & n12809) | (n12708 & n16056) | (n12809 & n16056);
  assign n16058 = (n12707 & n12809) | (n12707 & n16056) | (n12809 & n16056);
  assign n16059 = (n15940 & n16057) | (n15940 & n16058) | (n16057 & n16058);
  assign n12678 = (n15902 & n15968) | (n15902 & n15970) | (n15968 & n15970);
  assign n6246 = x72 & x80;
  assign n6247 = x71 & x81;
  assign n6248 = n6246 & n6247;
  assign n6249 = n6246 | n6247;
  assign n6250 = ~n6248 & n6249;
  assign n16060 = n6067 | n6069;
  assign n16062 = n6250 & n16060;
  assign n16063 = n6067 & n6250;
  assign n16064 = (n16019 & n16062) | (n16019 & n16063) | (n16062 & n16063);
  assign n16066 = (n16020 & n16062) | (n16020 & n16063) | (n16062 & n16063);
  assign n16067 = (n15915 & n16064) | (n15915 & n16066) | (n16064 & n16066);
  assign n16068 = (n15913 & n16064) | (n15913 & n16066) | (n16064 & n16066);
  assign n16069 = (n15794 & n16067) | (n15794 & n16068) | (n16067 & n16068);
  assign n16070 = n6250 | n16060;
  assign n16071 = n6067 | n6250;
  assign n16072 = (n16019 & n16070) | (n16019 & n16071) | (n16070 & n16071);
  assign n16073 = (n16020 & n16070) | (n16020 & n16071) | (n16070 & n16071);
  assign n16074 = (n15915 & n16072) | (n15915 & n16073) | (n16072 & n16073);
  assign n16075 = (n15913 & n16072) | (n15913 & n16073) | (n16072 & n16073);
  assign n16076 = (n15794 & n16074) | (n15794 & n16075) | (n16074 & n16075);
  assign n6253 = ~n16069 & n16076;
  assign n6254 = x70 & x82;
  assign n6255 = n6253 & n6254;
  assign n6256 = n6253 | n6254;
  assign n6257 = ~n6255 & n6256;
  assign n12818 = n6074 | n6076;
  assign n12829 = n6257 & n12818;
  assign n12830 = n6074 & n6257;
  assign n16017 = (n5901 & n15980) | (n5901 & n16015) | (n15980 & n16015);
  assign n16077 = (n12829 & n12830) | (n12829 & n16017) | (n12830 & n16017);
  assign n16078 = (n12829 & n12830) | (n12829 & n16016) | (n12830 & n16016);
  assign n16079 = (n15908 & n16077) | (n15908 & n16078) | (n16077 & n16078);
  assign n12832 = n6257 | n12818;
  assign n12833 = n6074 | n6257;
  assign n16080 = (n12832 & n12833) | (n12832 & n16017) | (n12833 & n16017);
  assign n16081 = (n12832 & n12833) | (n12832 & n16016) | (n12833 & n16016);
  assign n16082 = (n15908 & n16080) | (n15908 & n16081) | (n16080 & n16081);
  assign n6260 = ~n16079 & n16082;
  assign n6261 = x69 & x83;
  assign n6262 = n6260 & n6261;
  assign n6263 = n6260 | n6261;
  assign n6264 = ~n6262 & n6263;
  assign n16083 = n6081 | n6083;
  assign n16084 = (n6081 & n12756) | (n6081 & n16083) | (n12756 & n16083);
  assign n12835 = n6264 & n16084;
  assign n16085 = n5908 | n6081;
  assign n16086 = (n6081 & n6083) | (n6081 & n16085) | (n6083 & n16085);
  assign n12836 = n6264 & n16086;
  assign n12837 = (n12678 & n12835) | (n12678 & n12836) | (n12835 & n12836);
  assign n12838 = n6264 | n16084;
  assign n12839 = n6264 | n16086;
  assign n12840 = (n12678 & n12838) | (n12678 & n12839) | (n12838 & n12839);
  assign n6267 = ~n12837 & n12840;
  assign n6268 = x68 & x84;
  assign n6269 = n6267 & n6268;
  assign n6270 = n6267 | n6268;
  assign n6271 = ~n6269 & n6270;
  assign n12813 = n6088 | n6090;
  assign n12841 = n6271 & n12813;
  assign n12842 = n6088 & n6271;
  assign n16087 = (n12841 & n12842) | (n12841 & n16014) | (n12842 & n16014);
  assign n16088 = (n12841 & n12842) | (n12841 & n16012) | (n12842 & n16012);
  assign n16089 = (n15945 & n16087) | (n15945 & n16088) | (n16087 & n16088);
  assign n12844 = n6271 | n12813;
  assign n12845 = n6088 | n6271;
  assign n16090 = (n12844 & n12845) | (n12844 & n16014) | (n12845 & n16014);
  assign n16091 = (n12844 & n12845) | (n12844 & n16012) | (n12845 & n16012);
  assign n16092 = (n15945 & n16090) | (n15945 & n16091) | (n16090 & n16091);
  assign n6274 = ~n16089 & n16092;
  assign n6275 = x67 & x85;
  assign n6276 = n6274 & n6275;
  assign n6277 = n6274 | n6275;
  assign n6278 = ~n6276 & n6277;
  assign n12811 = n6095 | n6097;
  assign n12847 = n6278 & n12811;
  assign n12848 = n6095 & n6278;
  assign n12849 = (n16010 & n12847) | (n16010 & n12848) | (n12847 & n12848);
  assign n12850 = n6278 | n12811;
  assign n12851 = n6095 | n6278;
  assign n12852 = (n16010 & n12850) | (n16010 & n12851) | (n12850 & n12851);
  assign n6281 = ~n12849 & n12852;
  assign n6282 = x66 & x86;
  assign n6283 = n6281 & n6282;
  assign n6284 = n6281 | n6282;
  assign n6285 = ~n6283 & n6284;
  assign n12853 = n6102 & n6285;
  assign n16093 = (n6285 & n12777) | (n6285 & n12853) | (n12777 & n12853);
  assign n16094 = (n6285 & n12776) | (n6285 & n12853) | (n12776 & n12853);
  assign n16095 = (n15966 & n16093) | (n15966 & n16094) | (n16093 & n16094);
  assign n12855 = n6102 | n6285;
  assign n16096 = n12777 | n12855;
  assign n16097 = n12776 | n12855;
  assign n16098 = (n15966 & n16096) | (n15966 & n16097) | (n16096 & n16097);
  assign n6288 = ~n16095 & n16098;
  assign n6289 = x65 & x87;
  assign n6290 = n6288 & n6289;
  assign n6291 = n6288 | n6289;
  assign n6292 = ~n6290 & n6291;
  assign n6293 = n16059 & n6292;
  assign n6294 = n16059 | n6292;
  assign n6295 = ~n6293 & n6294;
  assign n6296 = x64 & x88;
  assign n6297 = n6295 & n6296;
  assign n6298 = n6295 | n6296;
  assign n6299 = ~n6297 & n6298;
  assign n12806 = n6116 | n6118;
  assign n12857 = n6299 & n12806;
  assign n12858 = n6116 & n6299;
  assign n12859 = (n16005 & n12857) | (n16005 & n12858) | (n12857 & n12858);
  assign n12860 = n6299 | n12806;
  assign n12861 = n6116 | n6299;
  assign n12862 = (n16005 & n12860) | (n16005 & n12861) | (n12860 & n12861);
  assign n6302 = ~n12859 & n12862;
  assign n6303 = x63 & x89;
  assign n6304 = n6302 & n6303;
  assign n6305 = n6302 | n6303;
  assign n6306 = ~n6304 & n6305;
  assign n12863 = n6123 & n6306;
  assign n16099 = (n6306 & n12786) | (n6306 & n12863) | (n12786 & n12863);
  assign n16100 = (n6125 & n6306) | (n6125 & n12863) | (n6306 & n12863);
  assign n16101 = (n12718 & n16099) | (n12718 & n16100) | (n16099 & n16100);
  assign n12865 = n6123 | n6306;
  assign n16102 = n12786 | n12865;
  assign n16103 = n6125 | n12865;
  assign n16104 = (n12718 & n16102) | (n12718 & n16103) | (n16102 & n16103);
  assign n6309 = ~n16101 & n16104;
  assign n6310 = x62 & x90;
  assign n6311 = n6309 & n6310;
  assign n6312 = n6309 | n6310;
  assign n6313 = ~n6311 & n6312;
  assign n6314 = n12805 & n6313;
  assign n6315 = n12805 | n6313;
  assign n6316 = ~n6314 & n6315;
  assign n6317 = x61 & x91;
  assign n6318 = n6316 & n6317;
  assign n6319 = n6316 | n6317;
  assign n6320 = ~n6318 & n6319;
  assign n6321 = n12803 & n6320;
  assign n6322 = n12803 | n6320;
  assign n6323 = ~n6321 & n6322;
  assign n6324 = x60 & x92;
  assign n6325 = n6323 & n6324;
  assign n6326 = n6323 | n6324;
  assign n6327 = ~n6325 & n6326;
  assign n6328 = n12801 & n6327;
  assign n6329 = n12801 | n6327;
  assign n6330 = ~n6328 & n6329;
  assign n6331 = x59 & x93;
  assign n6332 = n6330 & n6331;
  assign n6333 = n6330 | n6331;
  assign n6334 = ~n6332 & n6333;
  assign n6335 = n12799 & n6334;
  assign n6336 = n12799 | n6334;
  assign n6337 = ~n6335 & n6336;
  assign n6338 = x58 & x94;
  assign n6339 = n6337 & n6338;
  assign n6340 = n6337 | n6338;
  assign n6341 = ~n6339 & n6340;
  assign n6342 = n12797 & n6341;
  assign n6343 = n12797 | n6341;
  assign n6344 = ~n6342 & n6343;
  assign n6345 = x57 & x95;
  assign n6346 = n6344 & n6345;
  assign n6347 = n6344 | n6345;
  assign n6348 = ~n6346 & n6347;
  assign n6349 = n12795 & n6348;
  assign n6350 = n12795 | n6348;
  assign n6351 = ~n6349 & n6350;
  assign n6352 = x56 & x96;
  assign n6353 = n6351 & n6352;
  assign n6354 = n6351 | n6352;
  assign n6355 = ~n6353 & n6354;
  assign n6356 = n12793 & n6355;
  assign n6357 = n12793 | n6355;
  assign n6358 = ~n6356 & n6357;
  assign n6359 = x55 & x97;
  assign n6360 = n6358 & n6359;
  assign n6361 = n6358 | n6359;
  assign n6362 = ~n6360 & n6361;
  assign n6363 = n6229 & n6362;
  assign n6364 = n6229 | n6362;
  assign n6365 = ~n6363 & n6364;
  assign n6366 = x54 & x98;
  assign n6367 = n6365 & n6366;
  assign n6368 = n6365 | n6366;
  assign n6369 = ~n6367 & n6368;
  assign n6370 = n6228 & n6369;
  assign n6371 = n6228 | n6369;
  assign n6372 = ~n6370 & n6371;
  assign n6373 = x53 & x99;
  assign n6374 = n6372 & n6373;
  assign n6375 = n6372 | n6373;
  assign n6376 = ~n6374 & n6375;
  assign n6377 = n6227 & n6376;
  assign n6378 = n6227 | n6376;
  assign n6379 = ~n6377 & n6378;
  assign n6380 = x52 & x100;
  assign n6381 = n6379 & n6380;
  assign n6382 = n6379 | n6380;
  assign n6383 = ~n6381 & n6382;
  assign n6384 = n6226 & n6383;
  assign n6385 = n6226 | n6383;
  assign n6386 = ~n6384 & n6385;
  assign n6387 = x51 & x101;
  assign n6388 = n6386 & n6387;
  assign n6389 = n6386 | n6387;
  assign n6390 = ~n6388 & n6389;
  assign n6391 = n16054 & n6390;
  assign n6392 = n16054 | n6390;
  assign n6393 = ~n6391 & n6392;
  assign n6394 = x50 & x102;
  assign n6395 = n6393 & n6394;
  assign n6396 = n6393 | n6394;
  assign n6397 = ~n6395 & n6396;
  assign n6398 = n12791 & n6397;
  assign n6399 = n12791 | n6397;
  assign n6400 = ~n6398 & n6399;
  assign n6401 = x49 & x103;
  assign n6402 = n6400 & n6401;
  assign n6403 = n6400 | n6401;
  assign n6404 = ~n6402 & n6403;
  assign n6405 = n6221 & n6404;
  assign n6406 = n6221 | n6404;
  assign n6407 = ~n6405 & n6406;
  assign n6408 = x48 & x104;
  assign n6409 = n6407 & n6408;
  assign n6410 = n6407 | n6408;
  assign n6411 = ~n6409 & n6410;
  assign n17712 = n6220 | n6401;
  assign n17713 = (n6219 & n6401) | (n6219 & n17712) | (n6401 & n17712);
  assign n16106 = (n6221 & n6400) | (n6221 & n17713) | (n6400 & n17713);
  assign n12868 = (n6402 & n6404) | (n6402 & n16106) | (n6404 & n16106);
  assign n12869 = n6395 | n12791;
  assign n12870 = (n6395 & n6397) | (n6395 & n12869) | (n6397 & n12869);
  assign n16107 = n6388 | n16054;
  assign n16108 = (n6388 & n6390) | (n6388 & n16107) | (n6390 & n16107);
  assign n6415 = n6381 | n6384;
  assign n6416 = n6374 | n6377;
  assign n6417 = n6367 | n6370;
  assign n12871 = n6360 | n6362;
  assign n12872 = (n6229 & n6360) | (n6229 & n12871) | (n6360 & n12871);
  assign n12873 = n6353 | n6355;
  assign n12874 = (n6353 & n12793) | (n6353 & n12873) | (n12793 & n12873);
  assign n12875 = n6346 | n6348;
  assign n12876 = (n6346 & n12795) | (n6346 & n12875) | (n12795 & n12875);
  assign n12877 = n6339 | n6341;
  assign n12878 = (n6339 & n12797) | (n6339 & n12877) | (n12797 & n12877);
  assign n12879 = n6332 | n6334;
  assign n12880 = (n6332 & n12799) | (n6332 & n12879) | (n12799 & n12879);
  assign n12881 = n6325 | n6327;
  assign n12882 = (n6325 & n12801) | (n6325 & n12881) | (n12801 & n12881);
  assign n12883 = n6318 | n6320;
  assign n12884 = (n6318 & n12803) | (n6318 & n12883) | (n12803 & n12883);
  assign n12888 = n6304 | n6306;
  assign n16109 = n6123 | n6304;
  assign n16110 = (n6304 & n6306) | (n6304 & n16109) | (n6306 & n16109);
  assign n16111 = (n12786 & n12888) | (n12786 & n16110) | (n12888 & n16110);
  assign n16112 = (n6125 & n12888) | (n6125 & n16110) | (n12888 & n16110);
  assign n16113 = (n12718 & n16111) | (n12718 & n16112) | (n16111 & n16112);
  assign n12893 = n6283 | n6285;
  assign n16114 = n6102 | n6283;
  assign n16115 = (n6283 & n6285) | (n6283 & n16114) | (n6285 & n16114);
  assign n16116 = (n12777 & n12893) | (n12777 & n16115) | (n12893 & n16115);
  assign n16117 = (n12776 & n12893) | (n12776 & n16115) | (n12893 & n16115);
  assign n16118 = (n15966 & n16116) | (n15966 & n16117) | (n16116 & n16117);
  assign n12755 = (n15945 & n16012) | (n15945 & n16014) | (n16012 & n16014);
  assign n12901 = n6248 | n16064;
  assign n12902 = n6248 | n16066;
  assign n16121 = (n12901 & n12902) | (n12901 & n15915) | (n12902 & n15915);
  assign n16122 = (n12901 & n12902) | (n12901 & n15913) | (n12902 & n15913);
  assign n16123 = (n15794 & n16121) | (n15794 & n16122) | (n16121 & n16122);
  assign n6435 = x73 & x80;
  assign n6436 = x72 & x81;
  assign n6437 = n6435 & n6436;
  assign n6438 = n6435 | n6436;
  assign n6439 = ~n6437 & n6438;
  assign n6440 = n16123 & n6439;
  assign n6441 = n16123 | n6439;
  assign n6442 = ~n6440 & n6441;
  assign n6443 = x71 & x82;
  assign n6444 = n6442 & n6443;
  assign n6445 = n6442 | n6443;
  assign n6446 = ~n6444 & n6445;
  assign n16124 = n6255 | n6257;
  assign n16125 = (n6255 & n12818) | (n6255 & n16124) | (n12818 & n16124);
  assign n12904 = n6446 & n16125;
  assign n16126 = n6074 | n6255;
  assign n16127 = (n6255 & n6257) | (n6255 & n16126) | (n6257 & n16126);
  assign n12905 = n6446 & n16127;
  assign n16128 = (n12904 & n12905) | (n12904 & n16017) | (n12905 & n16017);
  assign n16129 = (n12904 & n12905) | (n12904 & n16016) | (n12905 & n16016);
  assign n16130 = (n15908 & n16128) | (n15908 & n16129) | (n16128 & n16129);
  assign n12907 = n6446 | n16125;
  assign n12908 = n6446 | n16127;
  assign n16131 = (n12907 & n12908) | (n12907 & n16017) | (n12908 & n16017);
  assign n16132 = (n12907 & n12908) | (n12907 & n16016) | (n12908 & n16016);
  assign n16133 = (n15908 & n16131) | (n15908 & n16132) | (n16131 & n16132);
  assign n6449 = ~n16130 & n16133;
  assign n6450 = x70 & x83;
  assign n6451 = n6449 & n6450;
  assign n6452 = n6449 | n6450;
  assign n6453 = ~n6451 & n6452;
  assign n12910 = n6262 & n6453;
  assign n17714 = (n6264 & n6453) | (n6264 & n12910) | (n6453 & n12910);
  assign n17715 = n6453 & n12910;
  assign n17716 = (n16084 & n17714) | (n16084 & n17715) | (n17714 & n17715);
  assign n16135 = (n6453 & n12836) | (n6453 & n12910) | (n12836 & n12910);
  assign n16136 = (n12678 & n17716) | (n12678 & n16135) | (n17716 & n16135);
  assign n12912 = n6262 | n6453;
  assign n17717 = n6264 | n12912;
  assign n17718 = (n12912 & n16084) | (n12912 & n17717) | (n16084 & n17717);
  assign n16138 = n12836 | n12912;
  assign n16139 = (n12678 & n17718) | (n12678 & n16138) | (n17718 & n16138);
  assign n6456 = ~n16136 & n16139;
  assign n6457 = x69 & x84;
  assign n6458 = n6456 & n6457;
  assign n6459 = n6456 | n6457;
  assign n6460 = ~n6458 & n6459;
  assign n17719 = n6269 & n6460;
  assign n17720 = (n6460 & n12841) | (n6460 & n17719) | (n12841 & n17719);
  assign n16119 = n6088 | n6269;
  assign n16120 = (n6269 & n6271) | (n6269 & n16119) | (n6271 & n16119);
  assign n16141 = n6460 & n16120;
  assign n16142 = (n12755 & n17720) | (n12755 & n16141) | (n17720 & n16141);
  assign n17721 = n6269 | n6460;
  assign n17722 = n12841 | n17721;
  assign n16144 = n6460 | n16120;
  assign n16145 = (n12755 & n17722) | (n12755 & n16144) | (n17722 & n16144);
  assign n6463 = ~n16142 & n16145;
  assign n6464 = x68 & x85;
  assign n6465 = n6463 & n6464;
  assign n6466 = n6463 | n6464;
  assign n6467 = ~n6465 & n6466;
  assign n12914 = n6276 & n6467;
  assign n16146 = (n6467 & n12847) | (n6467 & n12914) | (n12847 & n12914);
  assign n16147 = (n6467 & n12848) | (n6467 & n12914) | (n12848 & n12914);
  assign n16148 = (n16010 & n16146) | (n16010 & n16147) | (n16146 & n16147);
  assign n12916 = n6276 | n6467;
  assign n16149 = n12847 | n12916;
  assign n16150 = n12848 | n12916;
  assign n16151 = (n16010 & n16149) | (n16010 & n16150) | (n16149 & n16150);
  assign n6470 = ~n16148 & n16151;
  assign n6471 = x67 & x86;
  assign n6472 = n6470 & n6471;
  assign n6473 = n6470 | n6471;
  assign n6474 = ~n6472 & n6473;
  assign n6475 = n16118 & n6474;
  assign n6476 = n16118 | n6474;
  assign n6477 = ~n6475 & n6476;
  assign n6478 = x66 & x87;
  assign n6479 = n6477 & n6478;
  assign n6480 = n6477 | n6478;
  assign n6481 = ~n6479 & n6480;
  assign n12890 = n6290 | n6292;
  assign n12918 = n6481 & n12890;
  assign n12919 = n6290 & n6481;
  assign n12920 = (n16059 & n12918) | (n16059 & n12919) | (n12918 & n12919);
  assign n12921 = n6481 | n12890;
  assign n12922 = n6290 | n6481;
  assign n12923 = (n16059 & n12921) | (n16059 & n12922) | (n12921 & n12922);
  assign n6484 = ~n12920 & n12923;
  assign n6485 = x65 & x88;
  assign n6486 = n6484 & n6485;
  assign n6487 = n6484 | n6485;
  assign n6488 = ~n6486 & n6487;
  assign n12924 = n6297 & n6488;
  assign n16152 = (n6488 & n12858) | (n6488 & n12924) | (n12858 & n12924);
  assign n16153 = (n6488 & n12857) | (n6488 & n12924) | (n12857 & n12924);
  assign n16154 = (n16005 & n16152) | (n16005 & n16153) | (n16152 & n16153);
  assign n12926 = n6297 | n6488;
  assign n16155 = n12858 | n12926;
  assign n16156 = n12857 | n12926;
  assign n16157 = (n16005 & n16155) | (n16005 & n16156) | (n16155 & n16156);
  assign n6491 = ~n16154 & n16157;
  assign n6492 = x64 & x89;
  assign n6493 = n6491 & n6492;
  assign n6494 = n6491 | n6492;
  assign n6495 = ~n6493 & n6494;
  assign n6496 = n16113 & n6495;
  assign n6497 = n16113 | n6495;
  assign n6498 = ~n6496 & n6497;
  assign n6499 = x63 & x90;
  assign n6500 = n6498 & n6499;
  assign n6501 = n6498 | n6499;
  assign n6502 = ~n6500 & n6501;
  assign n12885 = n6311 | n6313;
  assign n16158 = n6502 & n12885;
  assign n16159 = n6311 & n6502;
  assign n16160 = (n12805 & n16158) | (n12805 & n16159) | (n16158 & n16159);
  assign n16161 = n6502 | n12885;
  assign n16162 = n6311 | n6502;
  assign n16163 = (n12805 & n16161) | (n12805 & n16162) | (n16161 & n16162);
  assign n6505 = ~n16160 & n16163;
  assign n6506 = x62 & x91;
  assign n6507 = n6505 & n6506;
  assign n6508 = n6505 | n6506;
  assign n6509 = ~n6507 & n6508;
  assign n6510 = n12884 & n6509;
  assign n6511 = n12884 | n6509;
  assign n6512 = ~n6510 & n6511;
  assign n6513 = x61 & x92;
  assign n6514 = n6512 & n6513;
  assign n6515 = n6512 | n6513;
  assign n6516 = ~n6514 & n6515;
  assign n6517 = n12882 & n6516;
  assign n6518 = n12882 | n6516;
  assign n6519 = ~n6517 & n6518;
  assign n6520 = x60 & x93;
  assign n6521 = n6519 & n6520;
  assign n6522 = n6519 | n6520;
  assign n6523 = ~n6521 & n6522;
  assign n6524 = n12880 & n6523;
  assign n6525 = n12880 | n6523;
  assign n6526 = ~n6524 & n6525;
  assign n6527 = x59 & x94;
  assign n6528 = n6526 & n6527;
  assign n6529 = n6526 | n6527;
  assign n6530 = ~n6528 & n6529;
  assign n6531 = n12878 & n6530;
  assign n6532 = n12878 | n6530;
  assign n6533 = ~n6531 & n6532;
  assign n6534 = x58 & x95;
  assign n6535 = n6533 & n6534;
  assign n6536 = n6533 | n6534;
  assign n6537 = ~n6535 & n6536;
  assign n6538 = n12876 & n6537;
  assign n6539 = n12876 | n6537;
  assign n6540 = ~n6538 & n6539;
  assign n6541 = x57 & x96;
  assign n6542 = n6540 & n6541;
  assign n6543 = n6540 | n6541;
  assign n6544 = ~n6542 & n6543;
  assign n6545 = n12874 & n6544;
  assign n6546 = n12874 | n6544;
  assign n6547 = ~n6545 & n6546;
  assign n6548 = x56 & x97;
  assign n6549 = n6547 & n6548;
  assign n6550 = n6547 | n6548;
  assign n6551 = ~n6549 & n6550;
  assign n6552 = n12872 & n6551;
  assign n6553 = n12872 | n6551;
  assign n6554 = ~n6552 & n6553;
  assign n6555 = x55 & x98;
  assign n6556 = n6554 & n6555;
  assign n6557 = n6554 | n6555;
  assign n6558 = ~n6556 & n6557;
  assign n6559 = n6417 & n6558;
  assign n6560 = n6417 | n6558;
  assign n6561 = ~n6559 & n6560;
  assign n6562 = x54 & x99;
  assign n6563 = n6561 & n6562;
  assign n6564 = n6561 | n6562;
  assign n6565 = ~n6563 & n6564;
  assign n6566 = n6416 & n6565;
  assign n6567 = n6416 | n6565;
  assign n6568 = ~n6566 & n6567;
  assign n6569 = x53 & x100;
  assign n6570 = n6568 & n6569;
  assign n6571 = n6568 | n6569;
  assign n6572 = ~n6570 & n6571;
  assign n6573 = n6415 & n6572;
  assign n6574 = n6415 | n6572;
  assign n6575 = ~n6573 & n6574;
  assign n6576 = x52 & x101;
  assign n6577 = n6575 & n6576;
  assign n6578 = n6575 | n6576;
  assign n6579 = ~n6577 & n6578;
  assign n6580 = n16108 & n6579;
  assign n6581 = n16108 | n6579;
  assign n6582 = ~n6580 & n6581;
  assign n6583 = x51 & x102;
  assign n6584 = n6582 & n6583;
  assign n6585 = n6582 | n6583;
  assign n6586 = ~n6584 & n6585;
  assign n6587 = n12870 & n6586;
  assign n6588 = n12870 | n6586;
  assign n6589 = ~n6587 & n6588;
  assign n6590 = x50 & x103;
  assign n6591 = n6589 & n6590;
  assign n6592 = n6589 | n6590;
  assign n6593 = ~n6591 & n6592;
  assign n6594 = n12868 & n6593;
  assign n6595 = n12868 | n6593;
  assign n6596 = ~n6594 & n6595;
  assign n6597 = x49 & x104;
  assign n6598 = n6596 & n6597;
  assign n6599 = n6596 | n6597;
  assign n6600 = ~n6598 & n6599;
  assign n6601 = n6409 & n6600;
  assign n6602 = n6409 | n6600;
  assign n6603 = ~n6601 & n6602;
  assign n6604 = x48 & x105;
  assign n6605 = n6603 & n6604;
  assign n6606 = n6603 | n6604;
  assign n6607 = ~n6605 & n6606;
  assign n17723 = n6408 | n6597;
  assign n17724 = (n6407 & n6597) | (n6407 & n17723) | (n6597 & n17723);
  assign n16165 = (n6409 & n6596) | (n6409 & n17724) | (n6596 & n17724);
  assign n12929 = (n6598 & n6600) | (n6598 & n16165) | (n6600 & n16165);
  assign n12930 = n6591 | n12868;
  assign n12931 = (n6591 & n6593) | (n6591 & n12930) | (n6593 & n12930);
  assign n12932 = n6584 | n12870;
  assign n12933 = (n6584 & n6586) | (n6584 & n12932) | (n6586 & n12932);
  assign n16166 = n6577 | n16108;
  assign n16167 = (n6577 & n6579) | (n6577 & n16166) | (n6579 & n16166);
  assign n6612 = n6570 | n6573;
  assign n6613 = n6563 | n6566;
  assign n12934 = n6556 | n6558;
  assign n12935 = (n6417 & n6556) | (n6417 & n12934) | (n6556 & n12934);
  assign n12936 = n6549 | n6551;
  assign n12937 = (n6549 & n12872) | (n6549 & n12936) | (n12872 & n12936);
  assign n12938 = n6542 | n6544;
  assign n12939 = (n6542 & n12874) | (n6542 & n12938) | (n12874 & n12938);
  assign n12940 = n6535 | n6537;
  assign n12941 = (n6535 & n12876) | (n6535 & n12940) | (n12876 & n12940);
  assign n12942 = n6528 | n6530;
  assign n12943 = (n6528 & n12878) | (n6528 & n12942) | (n12878 & n12942);
  assign n12944 = n6521 | n6523;
  assign n12945 = (n6521 & n12880) | (n6521 & n12944) | (n12880 & n12944);
  assign n12946 = n6514 | n6516;
  assign n12947 = (n6514 & n12882) | (n6514 & n12946) | (n12882 & n12946);
  assign n12886 = (n6311 & n12805) | (n6311 & n12885) | (n12805 & n12885);
  assign n12955 = n6486 | n6488;
  assign n16168 = n6297 | n6486;
  assign n16169 = (n6486 & n6488) | (n6486 & n16168) | (n6488 & n16168);
  assign n16170 = (n12858 & n12955) | (n12858 & n16169) | (n12955 & n16169);
  assign n16171 = (n12857 & n12955) | (n12857 & n16169) | (n12955 & n16169);
  assign n16172 = (n16005 & n16170) | (n16005 & n16171) | (n16170 & n16171);
  assign n12960 = n6465 | n6467;
  assign n16173 = n6276 | n6465;
  assign n16174 = (n6465 & n6467) | (n6465 & n16173) | (n6467 & n16173);
  assign n16175 = (n12847 & n12960) | (n12847 & n16174) | (n12960 & n16174);
  assign n16176 = (n12848 & n12960) | (n12848 & n16174) | (n12960 & n16174);
  assign n16177 = (n16010 & n16175) | (n16010 & n16176) | (n16175 & n16176);
  assign n12895 = n6269 | n12841;
  assign n12968 = n6444 | n12905;
  assign n16178 = n6444 | n6446;
  assign n16179 = (n6444 & n16125) | (n6444 & n16178) | (n16125 & n16178);
  assign n16180 = (n12968 & n16017) | (n12968 & n16179) | (n16017 & n16179);
  assign n16181 = (n12968 & n16016) | (n12968 & n16179) | (n16016 & n16179);
  assign n16182 = (n15908 & n16180) | (n15908 & n16181) | (n16180 & n16181);
  assign n6632 = x74 & x80;
  assign n6633 = x73 & x81;
  assign n6634 = n6632 & n6633;
  assign n6635 = n6632 | n6633;
  assign n6636 = ~n6634 & n6635;
  assign n12970 = n6437 | n6439;
  assign n12972 = n6636 & n12970;
  assign n12973 = n6437 & n6636;
  assign n12974 = (n16123 & n12972) | (n16123 & n12973) | (n12972 & n12973);
  assign n12975 = n6636 | n12970;
  assign n12976 = n6437 | n6636;
  assign n12977 = (n16123 & n12975) | (n16123 & n12976) | (n12975 & n12976);
  assign n6639 = ~n12974 & n12977;
  assign n6640 = x72 & x82;
  assign n6641 = n6639 & n6640;
  assign n6642 = n6639 | n6640;
  assign n6643 = ~n6641 & n6642;
  assign n6644 = n16182 & n6643;
  assign n6645 = n16182 | n6643;
  assign n6646 = ~n6644 & n6645;
  assign n6647 = x71 & x83;
  assign n6648 = n6646 & n6647;
  assign n6649 = n6646 | n6647;
  assign n6650 = ~n6648 & n6649;
  assign n16183 = n6262 | n6451;
  assign n16184 = (n6451 & n6453) | (n6451 & n16183) | (n6453 & n16183);
  assign n12978 = n6650 & n16184;
  assign n12965 = n6451 | n6453;
  assign n12979 = n6650 & n12965;
  assign n16185 = (n12835 & n12978) | (n12835 & n12979) | (n12978 & n12979);
  assign n16186 = (n12836 & n12978) | (n12836 & n12979) | (n12978 & n12979);
  assign n16187 = (n12678 & n16185) | (n12678 & n16186) | (n16185 & n16186);
  assign n12981 = n6650 | n16184;
  assign n12982 = n6650 | n12965;
  assign n16188 = (n12835 & n12981) | (n12835 & n12982) | (n12981 & n12982);
  assign n16189 = (n12836 & n12981) | (n12836 & n12982) | (n12981 & n12982);
  assign n16190 = (n12678 & n16188) | (n12678 & n16189) | (n16188 & n16189);
  assign n6653 = ~n16187 & n16190;
  assign n6654 = x70 & x84;
  assign n6655 = n6653 & n6654;
  assign n6656 = n6653 | n6654;
  assign n6657 = ~n6655 & n6656;
  assign n12962 = n6458 | n6460;
  assign n12984 = n6657 & n12962;
  assign n12985 = n6458 & n6657;
  assign n16191 = (n12895 & n12984) | (n12895 & n12985) | (n12984 & n12985);
  assign n16192 = (n12984 & n12985) | (n12984 & n16120) | (n12985 & n16120);
  assign n16193 = (n12755 & n16191) | (n12755 & n16192) | (n16191 & n16192);
  assign n12987 = n6657 | n12962;
  assign n12988 = n6458 | n6657;
  assign n16194 = (n12895 & n12987) | (n12895 & n12988) | (n12987 & n12988);
  assign n16195 = (n12987 & n12988) | (n12987 & n16120) | (n12988 & n16120);
  assign n16196 = (n12755 & n16194) | (n12755 & n16195) | (n16194 & n16195);
  assign n6660 = ~n16193 & n16196;
  assign n6661 = x69 & x85;
  assign n6662 = n6660 & n6661;
  assign n6663 = n6660 | n6661;
  assign n6664 = ~n6662 & n6663;
  assign n6665 = n16177 & n6664;
  assign n6666 = n16177 | n6664;
  assign n6667 = ~n6665 & n6666;
  assign n6668 = x68 & x86;
  assign n6669 = n6667 & n6668;
  assign n6670 = n6667 | n6668;
  assign n6671 = ~n6669 & n6670;
  assign n12957 = n6472 | n6474;
  assign n12990 = n6671 & n12957;
  assign n12991 = n6472 & n6671;
  assign n12992 = (n16118 & n12990) | (n16118 & n12991) | (n12990 & n12991);
  assign n12993 = n6671 | n12957;
  assign n12994 = n6472 | n6671;
  assign n12995 = (n16118 & n12993) | (n16118 & n12994) | (n12993 & n12994);
  assign n6674 = ~n12992 & n12995;
  assign n6675 = x67 & x87;
  assign n6676 = n6674 & n6675;
  assign n6677 = n6674 | n6675;
  assign n6678 = ~n6676 & n6677;
  assign n12996 = n6479 & n6678;
  assign n16197 = (n6678 & n12919) | (n6678 & n12996) | (n12919 & n12996);
  assign n16198 = (n6678 & n12918) | (n6678 & n12996) | (n12918 & n12996);
  assign n16199 = (n16059 & n16197) | (n16059 & n16198) | (n16197 & n16198);
  assign n12998 = n6479 | n6678;
  assign n16200 = n12919 | n12998;
  assign n16201 = n12918 | n12998;
  assign n16202 = (n16059 & n16200) | (n16059 & n16201) | (n16200 & n16201);
  assign n6681 = ~n16199 & n16202;
  assign n6682 = x66 & x88;
  assign n6683 = n6681 & n6682;
  assign n6684 = n6681 | n6682;
  assign n6685 = ~n6683 & n6684;
  assign n6686 = n16172 & n6685;
  assign n6687 = n16172 | n6685;
  assign n6688 = ~n6686 & n6687;
  assign n6689 = x65 & x89;
  assign n6690 = n6688 & n6689;
  assign n6691 = n6688 | n6689;
  assign n6692 = ~n6690 & n6691;
  assign n12952 = n6493 | n6495;
  assign n13000 = n6692 & n12952;
  assign n13001 = n6493 & n6692;
  assign n13002 = (n16113 & n13000) | (n16113 & n13001) | (n13000 & n13001);
  assign n13003 = n6692 | n12952;
  assign n13004 = n6493 | n6692;
  assign n13005 = (n16113 & n13003) | (n16113 & n13004) | (n13003 & n13004);
  assign n6695 = ~n13002 & n13005;
  assign n6696 = x64 & x90;
  assign n6697 = n6695 & n6696;
  assign n6698 = n6695 | n6696;
  assign n6699 = ~n6697 & n6698;
  assign n12950 = n6500 | n6502;
  assign n16203 = n6699 & n12950;
  assign n16204 = n6500 & n6699;
  assign n16205 = (n12886 & n16203) | (n12886 & n16204) | (n16203 & n16204);
  assign n16206 = n6699 | n12950;
  assign n16207 = n6500 | n6699;
  assign n16208 = (n12886 & n16206) | (n12886 & n16207) | (n16206 & n16207);
  assign n6702 = ~n16205 & n16208;
  assign n6703 = x63 & x91;
  assign n6704 = n6702 & n6703;
  assign n6705 = n6702 | n6703;
  assign n6706 = ~n6704 & n6705;
  assign n12948 = n6507 | n6509;
  assign n16209 = n6706 & n12948;
  assign n16210 = n6507 & n6706;
  assign n16211 = (n12884 & n16209) | (n12884 & n16210) | (n16209 & n16210);
  assign n16212 = n6706 | n12948;
  assign n16213 = n6507 | n6706;
  assign n16214 = (n12884 & n16212) | (n12884 & n16213) | (n16212 & n16213);
  assign n6709 = ~n16211 & n16214;
  assign n6710 = x62 & x92;
  assign n6711 = n6709 & n6710;
  assign n6712 = n6709 | n6710;
  assign n6713 = ~n6711 & n6712;
  assign n6714 = n12947 & n6713;
  assign n6715 = n12947 | n6713;
  assign n6716 = ~n6714 & n6715;
  assign n6717 = x61 & x93;
  assign n6718 = n6716 & n6717;
  assign n6719 = n6716 | n6717;
  assign n6720 = ~n6718 & n6719;
  assign n6721 = n12945 & n6720;
  assign n6722 = n12945 | n6720;
  assign n6723 = ~n6721 & n6722;
  assign n6724 = x60 & x94;
  assign n6725 = n6723 & n6724;
  assign n6726 = n6723 | n6724;
  assign n6727 = ~n6725 & n6726;
  assign n6728 = n12943 & n6727;
  assign n6729 = n12943 | n6727;
  assign n6730 = ~n6728 & n6729;
  assign n6731 = x59 & x95;
  assign n6732 = n6730 & n6731;
  assign n6733 = n6730 | n6731;
  assign n6734 = ~n6732 & n6733;
  assign n6735 = n12941 & n6734;
  assign n6736 = n12941 | n6734;
  assign n6737 = ~n6735 & n6736;
  assign n6738 = x58 & x96;
  assign n6739 = n6737 & n6738;
  assign n6740 = n6737 | n6738;
  assign n6741 = ~n6739 & n6740;
  assign n6742 = n12939 & n6741;
  assign n6743 = n12939 | n6741;
  assign n6744 = ~n6742 & n6743;
  assign n6745 = x57 & x97;
  assign n6746 = n6744 & n6745;
  assign n6747 = n6744 | n6745;
  assign n6748 = ~n6746 & n6747;
  assign n6749 = n12937 & n6748;
  assign n6750 = n12937 | n6748;
  assign n6751 = ~n6749 & n6750;
  assign n6752 = x56 & x98;
  assign n6753 = n6751 & n6752;
  assign n6754 = n6751 | n6752;
  assign n6755 = ~n6753 & n6754;
  assign n6756 = n12935 & n6755;
  assign n6757 = n12935 | n6755;
  assign n6758 = ~n6756 & n6757;
  assign n6759 = x55 & x99;
  assign n6760 = n6758 & n6759;
  assign n6761 = n6758 | n6759;
  assign n6762 = ~n6760 & n6761;
  assign n6763 = n6613 & n6762;
  assign n6764 = n6613 | n6762;
  assign n6765 = ~n6763 & n6764;
  assign n6766 = x54 & x100;
  assign n6767 = n6765 & n6766;
  assign n6768 = n6765 | n6766;
  assign n6769 = ~n6767 & n6768;
  assign n6770 = n6612 & n6769;
  assign n6771 = n6612 | n6769;
  assign n6772 = ~n6770 & n6771;
  assign n6773 = x53 & x101;
  assign n6774 = n6772 & n6773;
  assign n6775 = n6772 | n6773;
  assign n6776 = ~n6774 & n6775;
  assign n6777 = n16167 & n6776;
  assign n6778 = n16167 | n6776;
  assign n6779 = ~n6777 & n6778;
  assign n6780 = x52 & x102;
  assign n6781 = n6779 & n6780;
  assign n6782 = n6779 | n6780;
  assign n6783 = ~n6781 & n6782;
  assign n6784 = n12933 & n6783;
  assign n6785 = n12933 | n6783;
  assign n6786 = ~n6784 & n6785;
  assign n6787 = x51 & x103;
  assign n6788 = n6786 & n6787;
  assign n6789 = n6786 | n6787;
  assign n6790 = ~n6788 & n6789;
  assign n6791 = n12931 & n6790;
  assign n6792 = n12931 | n6790;
  assign n6793 = ~n6791 & n6792;
  assign n6794 = x50 & x104;
  assign n6795 = n6793 & n6794;
  assign n6796 = n6793 | n6794;
  assign n6797 = ~n6795 & n6796;
  assign n6798 = n12929 & n6797;
  assign n6799 = n12929 | n6797;
  assign n6800 = ~n6798 & n6799;
  assign n6801 = x49 & x105;
  assign n6802 = n6800 & n6801;
  assign n6803 = n6800 | n6801;
  assign n6804 = ~n6802 & n6803;
  assign n6805 = n6605 & n6804;
  assign n6806 = n6605 | n6804;
  assign n6807 = ~n6805 & n6806;
  assign n6808 = x48 & x106;
  assign n6809 = n6807 & n6808;
  assign n6810 = n6807 | n6808;
  assign n6811 = ~n6809 & n6810;
  assign n17725 = n6604 | n6801;
  assign n17726 = (n6603 & n6801) | (n6603 & n17725) | (n6801 & n17725);
  assign n16216 = (n6605 & n6800) | (n6605 & n17726) | (n6800 & n17726);
  assign n13007 = (n6802 & n6804) | (n6802 & n16216) | (n6804 & n16216);
  assign n13008 = n6795 | n12929;
  assign n13009 = (n6795 & n6797) | (n6795 & n13008) | (n6797 & n13008);
  assign n13010 = n6788 | n12931;
  assign n13011 = (n6788 & n6790) | (n6788 & n13010) | (n6790 & n13010);
  assign n13012 = n6781 | n12933;
  assign n13013 = (n6781 & n6783) | (n6781 & n13012) | (n6783 & n13012);
  assign n16217 = n6774 | n16167;
  assign n16218 = (n6774 & n6776) | (n6774 & n16217) | (n6776 & n16217);
  assign n6817 = n6767 | n6770;
  assign n13014 = n6760 | n6762;
  assign n13015 = (n6613 & n6760) | (n6613 & n13014) | (n6760 & n13014);
  assign n13016 = n6753 | n6755;
  assign n13017 = (n6753 & n12935) | (n6753 & n13016) | (n12935 & n13016);
  assign n13018 = n6746 | n6748;
  assign n13019 = (n6746 & n12937) | (n6746 & n13018) | (n12937 & n13018);
  assign n13020 = n6739 | n6741;
  assign n13021 = (n6739 & n12939) | (n6739 & n13020) | (n12939 & n13020);
  assign n13022 = n6732 | n6734;
  assign n13023 = (n6732 & n12941) | (n6732 & n13022) | (n12941 & n13022);
  assign n13024 = n6725 | n6727;
  assign n13025 = (n6725 & n12943) | (n6725 & n13024) | (n12943 & n13024);
  assign n13026 = n6718 | n6720;
  assign n13027 = (n6718 & n12945) | (n6718 & n13026) | (n12945 & n13026);
  assign n12949 = (n6507 & n12884) | (n6507 & n12948) | (n12884 & n12948);
  assign n12951 = (n6500 & n12886) | (n6500 & n12950) | (n12886 & n12950);
  assign n13037 = n6676 | n6678;
  assign n16219 = n6479 | n6676;
  assign n16220 = (n6676 & n6678) | (n6676 & n16219) | (n6678 & n16219);
  assign n16221 = (n12919 & n13037) | (n12919 & n16220) | (n13037 & n16220);
  assign n16222 = (n12918 & n13037) | (n12918 & n16220) | (n13037 & n16220);
  assign n16223 = (n16059 & n16221) | (n16059 & n16222) | (n16221 & n16222);
  assign n16224 = n6655 | n6657;
  assign n16225 = (n6655 & n12962) | (n6655 & n16224) | (n12962 & n16224);
  assign n16226 = n6458 | n6655;
  assign n16227 = (n6655 & n6657) | (n6655 & n16226) | (n6657 & n16226);
  assign n16228 = (n12895 & n16225) | (n12895 & n16227) | (n16225 & n16227);
  assign n16229 = (n16120 & n16225) | (n16120 & n16227) | (n16225 & n16227);
  assign n16230 = (n12755 & n16228) | (n12755 & n16229) | (n16228 & n16229);
  assign n13044 = n6648 | n12978;
  assign n13045 = n6648 | n12979;
  assign n16231 = (n12835 & n13044) | (n12835 & n13045) | (n13044 & n13045);
  assign n16232 = (n12836 & n13044) | (n12836 & n13045) | (n13044 & n13045);
  assign n16233 = (n12678 & n16231) | (n12678 & n16232) | (n16231 & n16232);
  assign n6837 = x75 & x80;
  assign n6838 = x74 & x81;
  assign n6839 = n6837 & n6838;
  assign n6840 = n6837 | n6838;
  assign n6841 = ~n6839 & n6840;
  assign n16234 = n6634 | n6636;
  assign n16235 = (n6634 & n12970) | (n6634 & n16234) | (n12970 & n16234);
  assign n13052 = n6841 & n16235;
  assign n16236 = n6437 | n6634;
  assign n16237 = (n6634 & n6636) | (n6634 & n16236) | (n6636 & n16236);
  assign n13053 = n6841 & n16237;
  assign n13054 = (n16123 & n13052) | (n16123 & n13053) | (n13052 & n13053);
  assign n13055 = n6841 | n16235;
  assign n13056 = n6841 | n16237;
  assign n13057 = (n16123 & n13055) | (n16123 & n13056) | (n13055 & n13056);
  assign n6844 = ~n13054 & n13057;
  assign n6845 = x73 & x82;
  assign n6846 = n6844 & n6845;
  assign n6847 = n6844 | n6845;
  assign n6848 = ~n6846 & n6847;
  assign n13047 = n6641 | n6643;
  assign n13058 = n6848 & n13047;
  assign n13059 = n6641 & n6848;
  assign n13060 = (n16182 & n13058) | (n16182 & n13059) | (n13058 & n13059);
  assign n13061 = n6848 | n13047;
  assign n13062 = n6641 | n6848;
  assign n13063 = (n16182 & n13061) | (n16182 & n13062) | (n13061 & n13062);
  assign n6851 = ~n13060 & n13063;
  assign n6852 = x72 & x83;
  assign n6853 = n6851 & n6852;
  assign n6854 = n6851 | n6852;
  assign n6855 = ~n6853 & n6854;
  assign n6856 = n16233 & n6855;
  assign n6857 = n16233 | n6855;
  assign n6858 = ~n6856 & n6857;
  assign n6859 = x71 & x84;
  assign n6860 = n6858 & n6859;
  assign n6861 = n6858 | n6859;
  assign n6862 = ~n6860 & n6861;
  assign n6863 = n16230 & n6862;
  assign n6864 = n16230 | n6862;
  assign n6865 = ~n6863 & n6864;
  assign n6866 = x70 & x85;
  assign n6867 = n6865 & n6866;
  assign n6868 = n6865 | n6866;
  assign n6869 = ~n6867 & n6868;
  assign n13039 = n6662 | n6664;
  assign n13064 = n6869 & n13039;
  assign n13065 = n6662 & n6869;
  assign n13066 = (n16177 & n13064) | (n16177 & n13065) | (n13064 & n13065);
  assign n13067 = n6869 | n13039;
  assign n13068 = n6662 | n6869;
  assign n13069 = (n16177 & n13067) | (n16177 & n13068) | (n13067 & n13068);
  assign n6872 = ~n13066 & n13069;
  assign n6873 = x69 & x86;
  assign n6874 = n6872 & n6873;
  assign n6875 = n6872 | n6873;
  assign n6876 = ~n6874 & n6875;
  assign n13070 = n6669 & n6876;
  assign n16238 = (n6876 & n12991) | (n6876 & n13070) | (n12991 & n13070);
  assign n16239 = (n6876 & n12990) | (n6876 & n13070) | (n12990 & n13070);
  assign n16240 = (n16118 & n16238) | (n16118 & n16239) | (n16238 & n16239);
  assign n13072 = n6669 | n6876;
  assign n16241 = n12991 | n13072;
  assign n16242 = n12990 | n13072;
  assign n16243 = (n16118 & n16241) | (n16118 & n16242) | (n16241 & n16242);
  assign n6879 = ~n16240 & n16243;
  assign n6880 = x68 & x87;
  assign n6881 = n6879 & n6880;
  assign n6882 = n6879 | n6880;
  assign n6883 = ~n6881 & n6882;
  assign n6884 = n16223 & n6883;
  assign n6885 = n16223 | n6883;
  assign n6886 = ~n6884 & n6885;
  assign n6887 = x67 & x88;
  assign n6888 = n6886 & n6887;
  assign n6889 = n6886 | n6887;
  assign n6890 = ~n6888 & n6889;
  assign n13034 = n6683 | n6685;
  assign n13074 = n6890 & n13034;
  assign n13075 = n6683 & n6890;
  assign n13076 = (n16172 & n13074) | (n16172 & n13075) | (n13074 & n13075);
  assign n13077 = n6890 | n13034;
  assign n13078 = n6683 | n6890;
  assign n13079 = (n16172 & n13077) | (n16172 & n13078) | (n13077 & n13078);
  assign n6893 = ~n13076 & n13079;
  assign n6894 = x66 & x89;
  assign n6895 = n6893 & n6894;
  assign n6896 = n6893 | n6894;
  assign n6897 = ~n6895 & n6896;
  assign n13080 = n6690 & n6897;
  assign n16244 = (n6897 & n13001) | (n6897 & n13080) | (n13001 & n13080);
  assign n16245 = (n6897 & n13000) | (n6897 & n13080) | (n13000 & n13080);
  assign n16246 = (n16113 & n16244) | (n16113 & n16245) | (n16244 & n16245);
  assign n13082 = n6690 | n6897;
  assign n16247 = n13001 | n13082;
  assign n16248 = n13000 | n13082;
  assign n16249 = (n16113 & n16247) | (n16113 & n16248) | (n16247 & n16248);
  assign n6900 = ~n16246 & n16249;
  assign n6901 = x65 & x90;
  assign n6902 = n6900 & n6901;
  assign n6903 = n6900 | n6901;
  assign n6904 = ~n6902 & n6903;
  assign n13032 = n6697 | n6699;
  assign n13084 = n6904 & n13032;
  assign n13085 = n6697 & n6904;
  assign n13086 = (n12951 & n13084) | (n12951 & n13085) | (n13084 & n13085);
  assign n13087 = n6904 | n13032;
  assign n13088 = n6697 | n6904;
  assign n13089 = (n12951 & n13087) | (n12951 & n13088) | (n13087 & n13088);
  assign n6907 = ~n13086 & n13089;
  assign n6908 = x64 & x91;
  assign n6909 = n6907 & n6908;
  assign n6910 = n6907 | n6908;
  assign n6911 = ~n6909 & n6910;
  assign n13030 = n6704 | n6706;
  assign n16250 = n6911 & n13030;
  assign n16251 = n6704 & n6911;
  assign n16252 = (n12949 & n16250) | (n12949 & n16251) | (n16250 & n16251);
  assign n16253 = n6911 | n13030;
  assign n16254 = n6704 | n6911;
  assign n16255 = (n12949 & n16253) | (n12949 & n16254) | (n16253 & n16254);
  assign n6914 = ~n16252 & n16255;
  assign n6915 = x63 & x92;
  assign n6916 = n6914 & n6915;
  assign n6917 = n6914 | n6915;
  assign n6918 = ~n6916 & n6917;
  assign n13028 = n6711 | n6713;
  assign n16256 = n6918 & n13028;
  assign n16257 = n6711 & n6918;
  assign n16258 = (n12947 & n16256) | (n12947 & n16257) | (n16256 & n16257);
  assign n16259 = n6918 | n13028;
  assign n16260 = n6711 | n6918;
  assign n16261 = (n12947 & n16259) | (n12947 & n16260) | (n16259 & n16260);
  assign n6921 = ~n16258 & n16261;
  assign n6922 = x62 & x93;
  assign n6923 = n6921 & n6922;
  assign n6924 = n6921 | n6922;
  assign n6925 = ~n6923 & n6924;
  assign n6926 = n13027 & n6925;
  assign n6927 = n13027 | n6925;
  assign n6928 = ~n6926 & n6927;
  assign n6929 = x61 & x94;
  assign n6930 = n6928 & n6929;
  assign n6931 = n6928 | n6929;
  assign n6932 = ~n6930 & n6931;
  assign n6933 = n13025 & n6932;
  assign n6934 = n13025 | n6932;
  assign n6935 = ~n6933 & n6934;
  assign n6936 = x60 & x95;
  assign n6937 = n6935 & n6936;
  assign n6938 = n6935 | n6936;
  assign n6939 = ~n6937 & n6938;
  assign n6940 = n13023 & n6939;
  assign n6941 = n13023 | n6939;
  assign n6942 = ~n6940 & n6941;
  assign n6943 = x59 & x96;
  assign n6944 = n6942 & n6943;
  assign n6945 = n6942 | n6943;
  assign n6946 = ~n6944 & n6945;
  assign n6947 = n13021 & n6946;
  assign n6948 = n13021 | n6946;
  assign n6949 = ~n6947 & n6948;
  assign n6950 = x58 & x97;
  assign n6951 = n6949 & n6950;
  assign n6952 = n6949 | n6950;
  assign n6953 = ~n6951 & n6952;
  assign n6954 = n13019 & n6953;
  assign n6955 = n13019 | n6953;
  assign n6956 = ~n6954 & n6955;
  assign n6957 = x57 & x98;
  assign n6958 = n6956 & n6957;
  assign n6959 = n6956 | n6957;
  assign n6960 = ~n6958 & n6959;
  assign n6961 = n13017 & n6960;
  assign n6962 = n13017 | n6960;
  assign n6963 = ~n6961 & n6962;
  assign n6964 = x56 & x99;
  assign n6965 = n6963 & n6964;
  assign n6966 = n6963 | n6964;
  assign n6967 = ~n6965 & n6966;
  assign n6968 = n13015 & n6967;
  assign n6969 = n13015 | n6967;
  assign n6970 = ~n6968 & n6969;
  assign n6971 = x55 & x100;
  assign n6972 = n6970 & n6971;
  assign n6973 = n6970 | n6971;
  assign n6974 = ~n6972 & n6973;
  assign n6975 = n6817 & n6974;
  assign n6976 = n6817 | n6974;
  assign n6977 = ~n6975 & n6976;
  assign n6978 = x54 & x101;
  assign n6979 = n6977 & n6978;
  assign n6980 = n6977 | n6978;
  assign n6981 = ~n6979 & n6980;
  assign n6982 = n16218 & n6981;
  assign n6983 = n16218 | n6981;
  assign n6984 = ~n6982 & n6983;
  assign n6985 = x53 & x102;
  assign n6986 = n6984 & n6985;
  assign n6987 = n6984 | n6985;
  assign n6988 = ~n6986 & n6987;
  assign n6989 = n13013 & n6988;
  assign n6990 = n13013 | n6988;
  assign n6991 = ~n6989 & n6990;
  assign n6992 = x52 & x103;
  assign n6993 = n6991 & n6992;
  assign n6994 = n6991 | n6992;
  assign n6995 = ~n6993 & n6994;
  assign n6996 = n13011 & n6995;
  assign n6997 = n13011 | n6995;
  assign n6998 = ~n6996 & n6997;
  assign n6999 = x51 & x104;
  assign n7000 = n6998 & n6999;
  assign n7001 = n6998 | n6999;
  assign n7002 = ~n7000 & n7001;
  assign n7003 = n13009 & n7002;
  assign n7004 = n13009 | n7002;
  assign n7005 = ~n7003 & n7004;
  assign n7006 = x50 & x105;
  assign n7007 = n7005 & n7006;
  assign n7008 = n7005 | n7006;
  assign n7009 = ~n7007 & n7008;
  assign n7010 = n13007 & n7009;
  assign n7011 = n13007 | n7009;
  assign n7012 = ~n7010 & n7011;
  assign n7013 = x49 & x106;
  assign n7014 = n7012 & n7013;
  assign n7015 = n7012 | n7013;
  assign n7016 = ~n7014 & n7015;
  assign n7017 = n6809 & n7016;
  assign n7018 = n6809 | n7016;
  assign n7019 = ~n7017 & n7018;
  assign n7020 = x48 & x107;
  assign n7021 = n7019 & n7020;
  assign n7022 = n7019 | n7020;
  assign n7023 = ~n7021 & n7022;
  assign n17727 = n6808 | n7013;
  assign n17728 = (n6807 & n7013) | (n6807 & n17727) | (n7013 & n17727);
  assign n16263 = (n6809 & n7012) | (n6809 & n17728) | (n7012 & n17728);
  assign n13091 = (n7014 & n7016) | (n7014 & n16263) | (n7016 & n16263);
  assign n13092 = n7007 | n13007;
  assign n13093 = (n7007 & n7009) | (n7007 & n13092) | (n7009 & n13092);
  assign n13094 = n7000 | n13009;
  assign n13095 = (n7000 & n7002) | (n7000 & n13094) | (n7002 & n13094);
  assign n13096 = n6993 | n13011;
  assign n13097 = (n6993 & n6995) | (n6993 & n13096) | (n6995 & n13096);
  assign n13098 = n6986 | n13013;
  assign n13099 = (n6986 & n6988) | (n6986 & n13098) | (n6988 & n13098);
  assign n16264 = n6979 | n16218;
  assign n16265 = (n6979 & n6981) | (n6979 & n16264) | (n6981 & n16264);
  assign n13100 = n6972 | n6974;
  assign n13101 = (n6817 & n6972) | (n6817 & n13100) | (n6972 & n13100);
  assign n13102 = n6965 | n6967;
  assign n13103 = (n6965 & n13015) | (n6965 & n13102) | (n13015 & n13102);
  assign n13104 = n6958 | n6960;
  assign n13105 = (n6958 & n13017) | (n6958 & n13104) | (n13017 & n13104);
  assign n13106 = n6951 | n6953;
  assign n13107 = (n6951 & n13019) | (n6951 & n13106) | (n13019 & n13106);
  assign n13108 = n6944 | n6946;
  assign n13109 = (n6944 & n13021) | (n6944 & n13108) | (n13021 & n13108);
  assign n13110 = n6937 | n6939;
  assign n13111 = (n6937 & n13023) | (n6937 & n13110) | (n13023 & n13110);
  assign n13112 = n6930 | n6932;
  assign n13113 = (n6930 & n13025) | (n6930 & n13112) | (n13025 & n13112);
  assign n13029 = (n6711 & n12947) | (n6711 & n13028) | (n12947 & n13028);
  assign n13031 = (n6704 & n12949) | (n6704 & n13030) | (n12949 & n13030);
  assign n13121 = n6895 | n6897;
  assign n16266 = n6690 | n6895;
  assign n16267 = (n6895 & n6897) | (n6895 & n16266) | (n6897 & n16266);
  assign n16268 = (n13001 & n13121) | (n13001 & n16267) | (n13121 & n16267);
  assign n16269 = (n13000 & n13121) | (n13000 & n16267) | (n13121 & n16267);
  assign n16270 = (n16113 & n16268) | (n16113 & n16269) | (n16268 & n16269);
  assign n13126 = n6874 | n6876;
  assign n16271 = n6669 | n6874;
  assign n16272 = (n6874 & n6876) | (n6874 & n16271) | (n6876 & n16271);
  assign n16273 = (n12991 & n13126) | (n12991 & n16272) | (n13126 & n16272);
  assign n16274 = (n12990 & n13126) | (n12990 & n16272) | (n13126 & n16272);
  assign n16275 = (n16118 & n16273) | (n16118 & n16274) | (n16273 & n16274);
  assign n16276 = n6662 | n6867;
  assign n16277 = (n6867 & n6869) | (n6867 & n16276) | (n6869 & n16276);
  assign n13129 = n6867 | n13064;
  assign n13130 = (n16177 & n16277) | (n16177 & n13129) | (n16277 & n13129);
  assign n7050 = x76 & x80;
  assign n7051 = x75 & x81;
  assign n7052 = n7050 & n7051;
  assign n7053 = n7050 | n7051;
  assign n7054 = ~n7052 & n7053;
  assign n16278 = n6839 | n6841;
  assign n16280 = n7054 & n16278;
  assign n16281 = n6839 & n7054;
  assign n16282 = (n16235 & n16280) | (n16235 & n16281) | (n16280 & n16281);
  assign n16283 = (n6839 & n16237) | (n6839 & n16278) | (n16237 & n16278);
  assign n13142 = n7054 & n16283;
  assign n13143 = (n16123 & n16282) | (n16123 & n13142) | (n16282 & n13142);
  assign n16284 = n7054 | n16278;
  assign n16285 = n6839 | n7054;
  assign n16286 = (n16235 & n16284) | (n16235 & n16285) | (n16284 & n16285);
  assign n13145 = n7054 | n16283;
  assign n13146 = (n16123 & n16286) | (n16123 & n13145) | (n16286 & n13145);
  assign n7057 = ~n13143 & n13146;
  assign n7058 = x74 & x82;
  assign n7059 = n7057 & n7058;
  assign n7060 = n7057 | n7058;
  assign n7061 = ~n7059 & n7060;
  assign n16287 = n6846 | n6848;
  assign n16288 = (n6846 & n13047) | (n6846 & n16287) | (n13047 & n16287);
  assign n13147 = n7061 & n16288;
  assign n16289 = n6641 | n6846;
  assign n16290 = (n6846 & n6848) | (n6846 & n16289) | (n6848 & n16289);
  assign n13148 = n7061 & n16290;
  assign n13149 = (n16182 & n13147) | (n16182 & n13148) | (n13147 & n13148);
  assign n13150 = n7061 | n16288;
  assign n13151 = n7061 | n16290;
  assign n13152 = (n16182 & n13150) | (n16182 & n13151) | (n13150 & n13151);
  assign n7064 = ~n13149 & n13152;
  assign n7065 = x73 & x83;
  assign n7066 = n7064 & n7065;
  assign n7067 = n7064 | n7065;
  assign n7068 = ~n7066 & n7067;
  assign n13133 = n6853 | n6855;
  assign n13153 = n7068 & n13133;
  assign n13154 = n6853 & n7068;
  assign n13155 = (n16233 & n13153) | (n16233 & n13154) | (n13153 & n13154);
  assign n13156 = n7068 | n13133;
  assign n13157 = n6853 | n7068;
  assign n13158 = (n16233 & n13156) | (n16233 & n13157) | (n13156 & n13157);
  assign n7071 = ~n13155 & n13158;
  assign n7072 = x72 & x84;
  assign n7073 = n7071 & n7072;
  assign n7074 = n7071 | n7072;
  assign n7075 = ~n7073 & n7074;
  assign n13131 = n6860 | n6862;
  assign n13159 = n7075 & n13131;
  assign n13160 = n6860 & n7075;
  assign n13161 = (n16230 & n13159) | (n16230 & n13160) | (n13159 & n13160);
  assign n13162 = n7075 | n13131;
  assign n13163 = n6860 | n7075;
  assign n13164 = (n16230 & n13162) | (n16230 & n13163) | (n13162 & n13163);
  assign n7078 = ~n13161 & n13164;
  assign n7079 = x71 & x85;
  assign n7080 = n7078 & n7079;
  assign n7081 = n7078 | n7079;
  assign n7082 = ~n7080 & n7081;
  assign n7083 = n13130 & n7082;
  assign n7084 = n13130 | n7082;
  assign n7085 = ~n7083 & n7084;
  assign n7086 = x70 & x86;
  assign n7087 = n7085 & n7086;
  assign n7088 = n7085 | n7086;
  assign n7089 = ~n7087 & n7088;
  assign n7090 = n16275 & n7089;
  assign n7091 = n16275 | n7089;
  assign n7092 = ~n7090 & n7091;
  assign n7093 = x69 & x87;
  assign n7094 = n7092 & n7093;
  assign n7095 = n7092 | n7093;
  assign n7096 = ~n7094 & n7095;
  assign n13123 = n6881 | n6883;
  assign n13165 = n7096 & n13123;
  assign n13166 = n6881 & n7096;
  assign n13167 = (n16223 & n13165) | (n16223 & n13166) | (n13165 & n13166);
  assign n13168 = n7096 | n13123;
  assign n13169 = n6881 | n7096;
  assign n13170 = (n16223 & n13168) | (n16223 & n13169) | (n13168 & n13169);
  assign n7099 = ~n13167 & n13170;
  assign n7100 = x68 & x88;
  assign n7101 = n7099 & n7100;
  assign n7102 = n7099 | n7100;
  assign n7103 = ~n7101 & n7102;
  assign n13171 = n6888 & n7103;
  assign n16291 = (n7103 & n13075) | (n7103 & n13171) | (n13075 & n13171);
  assign n16292 = (n7103 & n13074) | (n7103 & n13171) | (n13074 & n13171);
  assign n16293 = (n16172 & n16291) | (n16172 & n16292) | (n16291 & n16292);
  assign n13173 = n6888 | n7103;
  assign n16294 = n13075 | n13173;
  assign n16295 = n13074 | n13173;
  assign n16296 = (n16172 & n16294) | (n16172 & n16295) | (n16294 & n16295);
  assign n7106 = ~n16293 & n16296;
  assign n7107 = x67 & x89;
  assign n7108 = n7106 & n7107;
  assign n7109 = n7106 | n7107;
  assign n7110 = ~n7108 & n7109;
  assign n7111 = n16270 & n7110;
  assign n7112 = n16270 | n7110;
  assign n7113 = ~n7111 & n7112;
  assign n7114 = x66 & x90;
  assign n7115 = n7113 & n7114;
  assign n7116 = n7113 | n7114;
  assign n7117 = ~n7115 & n7116;
  assign n13175 = n6902 & n7117;
  assign n16297 = (n7117 & n13084) | (n7117 & n13175) | (n13084 & n13175);
  assign n16298 = (n7117 & n13085) | (n7117 & n13175) | (n13085 & n13175);
  assign n16299 = (n12951 & n16297) | (n12951 & n16298) | (n16297 & n16298);
  assign n13177 = n6902 | n7117;
  assign n16300 = n13084 | n13177;
  assign n16301 = n13085 | n13177;
  assign n16302 = (n12951 & n16300) | (n12951 & n16301) | (n16300 & n16301);
  assign n7120 = ~n16299 & n16302;
  assign n7121 = x65 & x91;
  assign n7122 = n7120 & n7121;
  assign n7123 = n7120 | n7121;
  assign n7124 = ~n7122 & n7123;
  assign n13118 = n6909 | n6911;
  assign n13179 = n7124 & n13118;
  assign n13180 = n6909 & n7124;
  assign n13181 = (n13031 & n13179) | (n13031 & n13180) | (n13179 & n13180);
  assign n13182 = n7124 | n13118;
  assign n13183 = n6909 | n7124;
  assign n13184 = (n13031 & n13182) | (n13031 & n13183) | (n13182 & n13183);
  assign n7127 = ~n13181 & n13184;
  assign n7128 = x64 & x92;
  assign n7129 = n7127 & n7128;
  assign n7130 = n7127 | n7128;
  assign n7131 = ~n7129 & n7130;
  assign n13116 = n6916 | n6918;
  assign n16303 = n7131 & n13116;
  assign n16304 = n6916 & n7131;
  assign n16305 = (n13029 & n16303) | (n13029 & n16304) | (n16303 & n16304);
  assign n16306 = n7131 | n13116;
  assign n16307 = n6916 | n7131;
  assign n16308 = (n13029 & n16306) | (n13029 & n16307) | (n16306 & n16307);
  assign n7134 = ~n16305 & n16308;
  assign n7135 = x63 & x93;
  assign n7136 = n7134 & n7135;
  assign n7137 = n7134 | n7135;
  assign n7138 = ~n7136 & n7137;
  assign n13114 = n6923 | n6925;
  assign n16309 = n7138 & n13114;
  assign n16310 = n6923 & n7138;
  assign n16311 = (n13027 & n16309) | (n13027 & n16310) | (n16309 & n16310);
  assign n16312 = n7138 | n13114;
  assign n16313 = n6923 | n7138;
  assign n16314 = (n13027 & n16312) | (n13027 & n16313) | (n16312 & n16313);
  assign n7141 = ~n16311 & n16314;
  assign n7142 = x62 & x94;
  assign n7143 = n7141 & n7142;
  assign n7144 = n7141 | n7142;
  assign n7145 = ~n7143 & n7144;
  assign n7146 = n13113 & n7145;
  assign n7147 = n13113 | n7145;
  assign n7148 = ~n7146 & n7147;
  assign n7149 = x61 & x95;
  assign n7150 = n7148 & n7149;
  assign n7151 = n7148 | n7149;
  assign n7152 = ~n7150 & n7151;
  assign n7153 = n13111 & n7152;
  assign n7154 = n13111 | n7152;
  assign n7155 = ~n7153 & n7154;
  assign n7156 = x60 & x96;
  assign n7157 = n7155 & n7156;
  assign n7158 = n7155 | n7156;
  assign n7159 = ~n7157 & n7158;
  assign n7160 = n13109 & n7159;
  assign n7161 = n13109 | n7159;
  assign n7162 = ~n7160 & n7161;
  assign n7163 = x59 & x97;
  assign n7164 = n7162 & n7163;
  assign n7165 = n7162 | n7163;
  assign n7166 = ~n7164 & n7165;
  assign n7167 = n13107 & n7166;
  assign n7168 = n13107 | n7166;
  assign n7169 = ~n7167 & n7168;
  assign n7170 = x58 & x98;
  assign n7171 = n7169 & n7170;
  assign n7172 = n7169 | n7170;
  assign n7173 = ~n7171 & n7172;
  assign n7174 = n13105 & n7173;
  assign n7175 = n13105 | n7173;
  assign n7176 = ~n7174 & n7175;
  assign n7177 = x57 & x99;
  assign n7178 = n7176 & n7177;
  assign n7179 = n7176 | n7177;
  assign n7180 = ~n7178 & n7179;
  assign n7181 = n13103 & n7180;
  assign n7182 = n13103 | n7180;
  assign n7183 = ~n7181 & n7182;
  assign n7184 = x56 & x100;
  assign n7185 = n7183 & n7184;
  assign n7186 = n7183 | n7184;
  assign n7187 = ~n7185 & n7186;
  assign n7188 = n13101 & n7187;
  assign n7189 = n13101 | n7187;
  assign n7190 = ~n7188 & n7189;
  assign n7191 = x55 & x101;
  assign n7192 = n7190 & n7191;
  assign n7193 = n7190 | n7191;
  assign n7194 = ~n7192 & n7193;
  assign n7195 = n16265 & n7194;
  assign n7196 = n16265 | n7194;
  assign n7197 = ~n7195 & n7196;
  assign n7198 = x54 & x102;
  assign n7199 = n7197 & n7198;
  assign n7200 = n7197 | n7198;
  assign n7201 = ~n7199 & n7200;
  assign n7202 = n13099 & n7201;
  assign n7203 = n13099 | n7201;
  assign n7204 = ~n7202 & n7203;
  assign n7205 = x53 & x103;
  assign n7206 = n7204 & n7205;
  assign n7207 = n7204 | n7205;
  assign n7208 = ~n7206 & n7207;
  assign n7209 = n13097 & n7208;
  assign n7210 = n13097 | n7208;
  assign n7211 = ~n7209 & n7210;
  assign n7212 = x52 & x104;
  assign n7213 = n7211 & n7212;
  assign n7214 = n7211 | n7212;
  assign n7215 = ~n7213 & n7214;
  assign n7216 = n13095 & n7215;
  assign n7217 = n13095 | n7215;
  assign n7218 = ~n7216 & n7217;
  assign n7219 = x51 & x105;
  assign n7220 = n7218 & n7219;
  assign n7221 = n7218 | n7219;
  assign n7222 = ~n7220 & n7221;
  assign n7223 = n13093 & n7222;
  assign n7224 = n13093 | n7222;
  assign n7225 = ~n7223 & n7224;
  assign n7226 = x50 & x106;
  assign n7227 = n7225 & n7226;
  assign n7228 = n7225 | n7226;
  assign n7229 = ~n7227 & n7228;
  assign n7230 = n13091 & n7229;
  assign n7231 = n13091 | n7229;
  assign n7232 = ~n7230 & n7231;
  assign n7233 = x49 & x107;
  assign n7234 = n7232 & n7233;
  assign n7235 = n7232 | n7233;
  assign n7236 = ~n7234 & n7235;
  assign n7237 = n7021 & n7236;
  assign n7238 = n7021 | n7236;
  assign n7239 = ~n7237 & n7238;
  assign n7240 = x48 & x108;
  assign n7241 = n7239 & n7240;
  assign n7242 = n7239 | n7240;
  assign n7243 = ~n7241 & n7242;
  assign n13185 = n7021 | n7234;
  assign n13186 = (n7234 & n7236) | (n7234 & n13185) | (n7236 & n13185);
  assign n13187 = n7227 | n13091;
  assign n13188 = (n7227 & n7229) | (n7227 & n13187) | (n7229 & n13187);
  assign n13189 = n7220 | n13093;
  assign n13190 = (n7220 & n7222) | (n7220 & n13189) | (n7222 & n13189);
  assign n13191 = n7213 | n13095;
  assign n13192 = (n7213 & n7215) | (n7213 & n13191) | (n7215 & n13191);
  assign n13193 = n7206 | n13097;
  assign n13194 = (n7206 & n7208) | (n7206 & n13193) | (n7208 & n13193);
  assign n13195 = n7199 | n13099;
  assign n13196 = (n7199 & n7201) | (n7199 & n13195) | (n7201 & n13195);
  assign n13197 = n7192 | n7194;
  assign n13198 = (n16265 & n7192) | (n16265 & n13197) | (n7192 & n13197);
  assign n13199 = n7185 | n7187;
  assign n13200 = (n7185 & n13101) | (n7185 & n13199) | (n13101 & n13199);
  assign n13201 = n7178 | n7180;
  assign n13202 = (n7178 & n13103) | (n7178 & n13201) | (n13103 & n13201);
  assign n13203 = n7171 | n7173;
  assign n13204 = (n7171 & n13105) | (n7171 & n13203) | (n13105 & n13203);
  assign n13205 = n7164 | n7166;
  assign n13206 = (n7164 & n13107) | (n7164 & n13205) | (n13107 & n13205);
  assign n13207 = n7157 | n7159;
  assign n13208 = (n7157 & n13109) | (n7157 & n13207) | (n13109 & n13207);
  assign n13209 = n7150 | n7152;
  assign n13210 = (n7150 & n13111) | (n7150 & n13209) | (n13111 & n13209);
  assign n13115 = (n6923 & n13027) | (n6923 & n13114) | (n13027 & n13114);
  assign n13117 = (n6916 & n13029) | (n6916 & n13116) | (n13029 & n13116);
  assign n13220 = n7101 | n7103;
  assign n16315 = n6888 | n7101;
  assign n16316 = (n7101 & n7103) | (n7101 & n16315) | (n7103 & n16315);
  assign n16317 = (n13075 & n13220) | (n13075 & n16316) | (n13220 & n16316);
  assign n16318 = (n13074 & n13220) | (n13074 & n16316) | (n13220 & n16316);
  assign n16319 = (n16172 & n16317) | (n16172 & n16318) | (n16317 & n16318);
  assign n7271 = x77 & x80;
  assign n7272 = x76 & x81;
  assign n7273 = n7271 & n7272;
  assign n7274 = n7271 | n7272;
  assign n7275 = ~n7273 & n7274;
  assign n16327 = n7052 & n7275;
  assign n16328 = (n7275 & n16282) | (n7275 & n16327) | (n16282 & n16327);
  assign n16329 = n7052 | n7054;
  assign n16331 = n7275 & n16329;
  assign n16332 = (n16283 & n16327) | (n16283 & n16331) | (n16327 & n16331);
  assign n13240 = (n16123 & n16328) | (n16123 & n16332) | (n16328 & n16332);
  assign n16333 = n7052 | n7275;
  assign n16334 = n16282 | n16333;
  assign n16335 = n7275 | n16329;
  assign n16336 = (n16283 & n16333) | (n16283 & n16335) | (n16333 & n16335);
  assign n13243 = (n16123 & n16334) | (n16123 & n16336) | (n16334 & n16336);
  assign n7278 = ~n13240 & n13243;
  assign n7279 = x75 & x82;
  assign n7280 = n7278 & n7279;
  assign n7281 = n7278 | n7279;
  assign n7282 = ~n7280 & n7281;
  assign n16324 = n7059 | n7061;
  assign n17729 = n7282 & n16324;
  assign n17730 = n7059 & n7282;
  assign n17731 = (n16288 & n17729) | (n16288 & n17730) | (n17729 & n17730);
  assign n16326 = (n7059 & n16290) | (n7059 & n16324) | (n16290 & n16324);
  assign n16338 = n7282 & n16326;
  assign n16339 = (n16182 & n17731) | (n16182 & n16338) | (n17731 & n16338);
  assign n17732 = n7282 | n16324;
  assign n17733 = n7059 | n7282;
  assign n17734 = (n16288 & n17732) | (n16288 & n17733) | (n17732 & n17733);
  assign n16341 = n7282 | n16326;
  assign n16342 = (n16182 & n17734) | (n16182 & n16341) | (n17734 & n16341);
  assign n7285 = ~n16339 & n16342;
  assign n7286 = x74 & x83;
  assign n7287 = n7285 & n7286;
  assign n7288 = n7285 | n7286;
  assign n7289 = ~n7287 & n7288;
  assign n16343 = n7066 | n7068;
  assign n16344 = (n7066 & n13133) | (n7066 & n16343) | (n13133 & n16343);
  assign n13244 = n7289 & n16344;
  assign n16345 = n6853 | n7066;
  assign n16346 = (n7066 & n7068) | (n7066 & n16345) | (n7068 & n16345);
  assign n13245 = n7289 & n16346;
  assign n13246 = (n16233 & n13244) | (n16233 & n13245) | (n13244 & n13245);
  assign n13247 = n7289 | n16344;
  assign n13248 = n7289 | n16346;
  assign n13249 = (n16233 & n13247) | (n16233 & n13248) | (n13247 & n13248);
  assign n7292 = ~n13246 & n13249;
  assign n7293 = x73 & x84;
  assign n7294 = n7292 & n7293;
  assign n7295 = n7292 | n7293;
  assign n7296 = ~n7294 & n7295;
  assign n16320 = n7073 | n7075;
  assign n16321 = (n7073 & n13131) | (n7073 & n16320) | (n13131 & n16320);
  assign n16347 = n7296 & n16321;
  assign n16322 = n6860 | n7073;
  assign n16323 = (n7073 & n7075) | (n7073 & n16322) | (n7075 & n16322);
  assign n16348 = n7296 & n16323;
  assign n16349 = (n16230 & n16347) | (n16230 & n16348) | (n16347 & n16348);
  assign n16350 = n7296 | n16321;
  assign n16351 = n7296 | n16323;
  assign n16352 = (n16230 & n16350) | (n16230 & n16351) | (n16350 & n16351);
  assign n7299 = ~n16349 & n16352;
  assign n7300 = x72 & x85;
  assign n7301 = n7299 & n7300;
  assign n7302 = n7299 | n7300;
  assign n7303 = ~n7301 & n7302;
  assign n13224 = n7080 | n7082;
  assign n13250 = n7303 & n13224;
  assign n13251 = n7080 & n7303;
  assign n13252 = (n13130 & n13250) | (n13130 & n13251) | (n13250 & n13251);
  assign n13253 = n7303 | n13224;
  assign n13254 = n7080 | n7303;
  assign n13255 = (n13130 & n13253) | (n13130 & n13254) | (n13253 & n13254);
  assign n7306 = ~n13252 & n13255;
  assign n7307 = x71 & x86;
  assign n7308 = n7306 & n7307;
  assign n7309 = n7306 | n7307;
  assign n7310 = ~n7308 & n7309;
  assign n13222 = n7087 | n7089;
  assign n13256 = n7310 & n13222;
  assign n13257 = n7087 & n7310;
  assign n13258 = (n16275 & n13256) | (n16275 & n13257) | (n13256 & n13257);
  assign n13259 = n7310 | n13222;
  assign n13260 = n7087 | n7310;
  assign n13261 = (n16275 & n13259) | (n16275 & n13260) | (n13259 & n13260);
  assign n7313 = ~n13258 & n13261;
  assign n7314 = x70 & x87;
  assign n7315 = n7313 & n7314;
  assign n7316 = n7313 | n7314;
  assign n7317 = ~n7315 & n7316;
  assign n13262 = n7094 & n7317;
  assign n16353 = (n7317 & n13166) | (n7317 & n13262) | (n13166 & n13262);
  assign n16354 = (n7317 & n13165) | (n7317 & n13262) | (n13165 & n13262);
  assign n16355 = (n16223 & n16353) | (n16223 & n16354) | (n16353 & n16354);
  assign n13264 = n7094 | n7317;
  assign n16356 = n13166 | n13264;
  assign n16357 = n13165 | n13264;
  assign n16358 = (n16223 & n16356) | (n16223 & n16357) | (n16356 & n16357);
  assign n7320 = ~n16355 & n16358;
  assign n7321 = x69 & x88;
  assign n7322 = n7320 & n7321;
  assign n7323 = n7320 | n7321;
  assign n7324 = ~n7322 & n7323;
  assign n7325 = n16319 & n7324;
  assign n7326 = n16319 | n7324;
  assign n7327 = ~n7325 & n7326;
  assign n7328 = x68 & x89;
  assign n7329 = n7327 & n7328;
  assign n7330 = n7327 | n7328;
  assign n7331 = ~n7329 & n7330;
  assign n13217 = n7108 | n7110;
  assign n13266 = n7331 & n13217;
  assign n13267 = n7108 & n7331;
  assign n13268 = (n16270 & n13266) | (n16270 & n13267) | (n13266 & n13267);
  assign n13269 = n7331 | n13217;
  assign n13270 = n7108 | n7331;
  assign n13271 = (n16270 & n13269) | (n16270 & n13270) | (n13269 & n13270);
  assign n7334 = ~n13268 & n13271;
  assign n7335 = x67 & x90;
  assign n7336 = n7334 & n7335;
  assign n7337 = n7334 | n7335;
  assign n7338 = ~n7336 & n7337;
  assign n13272 = n7115 & n7338;
  assign n13273 = (n7338 & n16299) | (n7338 & n13272) | (n16299 & n13272);
  assign n13274 = n7115 | n7338;
  assign n13275 = n16299 | n13274;
  assign n7341 = ~n13273 & n13275;
  assign n7342 = x66 & x91;
  assign n7343 = n7341 & n7342;
  assign n7344 = n7341 | n7342;
  assign n7345 = ~n7343 & n7344;
  assign n13276 = n7122 & n7345;
  assign n13277 = (n7345 & n13181) | (n7345 & n13276) | (n13181 & n13276);
  assign n13278 = n7122 | n7345;
  assign n13279 = n13181 | n13278;
  assign n7348 = ~n13277 & n13279;
  assign n7349 = x65 & x92;
  assign n7350 = n7348 & n7349;
  assign n7351 = n7348 | n7349;
  assign n7352 = ~n7350 & n7351;
  assign n13215 = n7129 | n7131;
  assign n13280 = n7352 & n13215;
  assign n13281 = n7129 & n7352;
  assign n13282 = (n13117 & n13280) | (n13117 & n13281) | (n13280 & n13281);
  assign n13283 = n7352 | n13215;
  assign n13284 = n7129 | n7352;
  assign n13285 = (n13117 & n13283) | (n13117 & n13284) | (n13283 & n13284);
  assign n7355 = ~n13282 & n13285;
  assign n7356 = x64 & x93;
  assign n7357 = n7355 & n7356;
  assign n7358 = n7355 | n7356;
  assign n7359 = ~n7357 & n7358;
  assign n13213 = n7136 | n7138;
  assign n16359 = n7359 & n13213;
  assign n16360 = n7136 & n7359;
  assign n16361 = (n13115 & n16359) | (n13115 & n16360) | (n16359 & n16360);
  assign n16362 = n7359 | n13213;
  assign n16363 = n7136 | n7359;
  assign n16364 = (n13115 & n16362) | (n13115 & n16363) | (n16362 & n16363);
  assign n7362 = ~n16361 & n16364;
  assign n7363 = x63 & x94;
  assign n7364 = n7362 & n7363;
  assign n7365 = n7362 | n7363;
  assign n7366 = ~n7364 & n7365;
  assign n13211 = n7143 | n7145;
  assign n16365 = n7366 & n13211;
  assign n16366 = n7143 & n7366;
  assign n16367 = (n13113 & n16365) | (n13113 & n16366) | (n16365 & n16366);
  assign n16368 = n7366 | n13211;
  assign n16369 = n7143 | n7366;
  assign n16370 = (n13113 & n16368) | (n13113 & n16369) | (n16368 & n16369);
  assign n7369 = ~n16367 & n16370;
  assign n7370 = x62 & x95;
  assign n7371 = n7369 & n7370;
  assign n7372 = n7369 | n7370;
  assign n7373 = ~n7371 & n7372;
  assign n7374 = n13210 & n7373;
  assign n7375 = n13210 | n7373;
  assign n7376 = ~n7374 & n7375;
  assign n7377 = x61 & x96;
  assign n7378 = n7376 & n7377;
  assign n7379 = n7376 | n7377;
  assign n7380 = ~n7378 & n7379;
  assign n7381 = n13208 & n7380;
  assign n7382 = n13208 | n7380;
  assign n7383 = ~n7381 & n7382;
  assign n7384 = x60 & x97;
  assign n7385 = n7383 & n7384;
  assign n7386 = n7383 | n7384;
  assign n7387 = ~n7385 & n7386;
  assign n7388 = n13206 & n7387;
  assign n7389 = n13206 | n7387;
  assign n7390 = ~n7388 & n7389;
  assign n7391 = x59 & x98;
  assign n7392 = n7390 & n7391;
  assign n7393 = n7390 | n7391;
  assign n7394 = ~n7392 & n7393;
  assign n7395 = n13204 & n7394;
  assign n7396 = n13204 | n7394;
  assign n7397 = ~n7395 & n7396;
  assign n7398 = x58 & x99;
  assign n7399 = n7397 & n7398;
  assign n7400 = n7397 | n7398;
  assign n7401 = ~n7399 & n7400;
  assign n7402 = n13202 & n7401;
  assign n7403 = n13202 | n7401;
  assign n7404 = ~n7402 & n7403;
  assign n7405 = x57 & x100;
  assign n7406 = n7404 & n7405;
  assign n7407 = n7404 | n7405;
  assign n7408 = ~n7406 & n7407;
  assign n7409 = n13200 & n7408;
  assign n7410 = n13200 | n7408;
  assign n7411 = ~n7409 & n7410;
  assign n7412 = x56 & x101;
  assign n7413 = n7411 & n7412;
  assign n7414 = n7411 | n7412;
  assign n7415 = ~n7413 & n7414;
  assign n7416 = n13198 & n7415;
  assign n7417 = n13198 | n7415;
  assign n7418 = ~n7416 & n7417;
  assign n7419 = x55 & x102;
  assign n7420 = n7418 & n7419;
  assign n7421 = n7418 | n7419;
  assign n7422 = ~n7420 & n7421;
  assign n7423 = n13196 & n7422;
  assign n7424 = n13196 | n7422;
  assign n7425 = ~n7423 & n7424;
  assign n7426 = x54 & x103;
  assign n7427 = n7425 & n7426;
  assign n7428 = n7425 | n7426;
  assign n7429 = ~n7427 & n7428;
  assign n7430 = n13194 & n7429;
  assign n7431 = n13194 | n7429;
  assign n7432 = ~n7430 & n7431;
  assign n7433 = x53 & x104;
  assign n7434 = n7432 & n7433;
  assign n7435 = n7432 | n7433;
  assign n7436 = ~n7434 & n7435;
  assign n7437 = n13192 & n7436;
  assign n7438 = n13192 | n7436;
  assign n7439 = ~n7437 & n7438;
  assign n7440 = x52 & x105;
  assign n7441 = n7439 & n7440;
  assign n7442 = n7439 | n7440;
  assign n7443 = ~n7441 & n7442;
  assign n7444 = n13190 & n7443;
  assign n7445 = n13190 | n7443;
  assign n7446 = ~n7444 & n7445;
  assign n7447 = x51 & x106;
  assign n7448 = n7446 & n7447;
  assign n7449 = n7446 | n7447;
  assign n7450 = ~n7448 & n7449;
  assign n7451 = n13188 & n7450;
  assign n7452 = n13188 | n7450;
  assign n7453 = ~n7451 & n7452;
  assign n7454 = x50 & x107;
  assign n7455 = n7453 & n7454;
  assign n7456 = n7453 | n7454;
  assign n7457 = ~n7455 & n7456;
  assign n7458 = n13186 & n7457;
  assign n7459 = n13186 | n7457;
  assign n7460 = ~n7458 & n7459;
  assign n7461 = x49 & x108;
  assign n7462 = n7460 & n7461;
  assign n7463 = n7460 | n7461;
  assign n7464 = ~n7462 & n7463;
  assign n7465 = n7241 & n7464;
  assign n7466 = n7241 | n7464;
  assign n7467 = ~n7465 & n7466;
  assign n7468 = x48 & x109;
  assign n7469 = n7467 & n7468;
  assign n7470 = n7467 | n7468;
  assign n7471 = ~n7469 & n7470;
  assign n17735 = n7240 | n7461;
  assign n17736 = (n7239 & n7461) | (n7239 & n17735) | (n7461 & n17735);
  assign n16372 = (n7241 & n7460) | (n7241 & n17736) | (n7460 & n17736);
  assign n13287 = (n7462 & n7464) | (n7462 & n16372) | (n7464 & n16372);
  assign n16373 = n7455 | n13186;
  assign n16374 = (n7455 & n7457) | (n7455 & n16373) | (n7457 & n16373);
  assign n7474 = n7448 | n7451;
  assign n7475 = n7441 | n7444;
  assign n7476 = n7434 | n7437;
  assign n7477 = n7427 | n7430;
  assign n7478 = n7420 | n7423;
  assign n13288 = n7413 | n7415;
  assign n13289 = (n7413 & n13198) | (n7413 & n13288) | (n13198 & n13288);
  assign n13290 = n7406 | n7408;
  assign n13291 = (n7406 & n13200) | (n7406 & n13290) | (n13200 & n13290);
  assign n13292 = n7399 | n7401;
  assign n13293 = (n7399 & n13202) | (n7399 & n13292) | (n13202 & n13292);
  assign n13294 = n7392 | n7394;
  assign n13295 = (n7392 & n13204) | (n7392 & n13294) | (n13204 & n13294);
  assign n13296 = n7385 | n7387;
  assign n13297 = (n7385 & n13206) | (n7385 & n13296) | (n13206 & n13296);
  assign n13298 = n7378 | n7380;
  assign n13299 = (n7378 & n13208) | (n7378 & n13298) | (n13208 & n13298);
  assign n13212 = (n7143 & n13113) | (n7143 & n13211) | (n13113 & n13211);
  assign n13214 = (n7136 & n13115) | (n7136 & n13213) | (n13115 & n13213);
  assign n13312 = n7315 | n7317;
  assign n16377 = n7094 | n7315;
  assign n16378 = (n7315 & n7317) | (n7315 & n16377) | (n7317 & n16377);
  assign n16379 = (n13166 & n13312) | (n13166 & n16378) | (n13312 & n16378);
  assign n16380 = (n13165 & n13312) | (n13165 & n16378) | (n13312 & n16378);
  assign n16381 = (n16223 & n16379) | (n16223 & n16380) | (n16379 & n16380);
  assign n7500 = x78 & x80;
  assign n7501 = x77 & x81;
  assign n7502 = n7500 & n7501;
  assign n7503 = n7500 | n7501;
  assign n7504 = ~n7502 & n7503;
  assign n17737 = n7273 & n7504;
  assign n17738 = (n7504 & n16332) | (n7504 & n17737) | (n16332 & n17737);
  assign n16387 = n7273 | n7275;
  assign n17741 = n7504 & n16387;
  assign n17739 = n7052 | n7273;
  assign n17740 = (n7273 & n7275) | (n7273 & n17739) | (n7275 & n17739);
  assign n17742 = n7504 & n17740;
  assign n17743 = (n16282 & n17741) | (n16282 & n17742) | (n17741 & n17742);
  assign n16391 = (n16123 & n17738) | (n16123 & n17743) | (n17738 & n17743);
  assign n17744 = n7273 | n7504;
  assign n17745 = n16332 | n17744;
  assign n17746 = n7504 | n16387;
  assign n17747 = n7504 | n17740;
  assign n17748 = (n16282 & n17746) | (n16282 & n17747) | (n17746 & n17747);
  assign n16394 = (n16123 & n17745) | (n16123 & n17748) | (n17745 & n17748);
  assign n7507 = ~n16391 & n16394;
  assign n7508 = x76 & x82;
  assign n7509 = n7507 & n7508;
  assign n7510 = n7507 | n7508;
  assign n7511 = ~n7509 & n7510;
  assign n13319 = n7280 | n7282;
  assign n13324 = n7511 & n13319;
  assign n13325 = n7280 & n7511;
  assign n16325 = (n7059 & n16288) | (n7059 & n16324) | (n16288 & n16324);
  assign n16395 = (n13324 & n13325) | (n13324 & n16325) | (n13325 & n16325);
  assign n16396 = (n13324 & n13325) | (n13324 & n16326) | (n13325 & n16326);
  assign n16397 = (n16182 & n16395) | (n16182 & n16396) | (n16395 & n16396);
  assign n13327 = n7511 | n13319;
  assign n13328 = n7280 | n7511;
  assign n16398 = (n13327 & n13328) | (n13327 & n16325) | (n13328 & n16325);
  assign n16399 = (n13327 & n13328) | (n13327 & n16326) | (n13328 & n16326);
  assign n16400 = (n16182 & n16398) | (n16182 & n16399) | (n16398 & n16399);
  assign n7514 = ~n16397 & n16400;
  assign n7515 = x75 & x83;
  assign n7516 = n7514 & n7515;
  assign n7517 = n7514 | n7515;
  assign n7518 = ~n7516 & n7517;
  assign n13330 = n7287 & n7518;
  assign n17749 = (n7289 & n7518) | (n7289 & n13330) | (n7518 & n13330);
  assign n17750 = n7518 & n13330;
  assign n17751 = (n16344 & n17749) | (n16344 & n17750) | (n17749 & n17750);
  assign n16402 = (n7518 & n13245) | (n7518 & n13330) | (n13245 & n13330);
  assign n16403 = (n16233 & n17751) | (n16233 & n16402) | (n17751 & n16402);
  assign n13332 = n7287 | n7518;
  assign n17752 = n7289 | n13332;
  assign n17753 = (n13332 & n16344) | (n13332 & n17752) | (n16344 & n17752);
  assign n16405 = n13245 | n13332;
  assign n16406 = (n16233 & n17753) | (n16233 & n16405) | (n17753 & n16405);
  assign n7521 = ~n16403 & n16406;
  assign n7522 = x74 & x84;
  assign n7523 = n7521 & n7522;
  assign n7524 = n7521 | n7522;
  assign n7525 = ~n7523 & n7524;
  assign n13317 = n7294 | n7296;
  assign n13334 = n7525 & n13317;
  assign n13335 = n7294 & n7525;
  assign n16407 = (n13334 & n13335) | (n13334 & n16321) | (n13335 & n16321);
  assign n16408 = (n13334 & n13335) | (n13334 & n16323) | (n13335 & n16323);
  assign n16409 = (n16230 & n16407) | (n16230 & n16408) | (n16407 & n16408);
  assign n13337 = n7525 | n13317;
  assign n13338 = n7294 | n7525;
  assign n16410 = (n13337 & n13338) | (n13337 & n16321) | (n13338 & n16321);
  assign n16411 = (n13337 & n13338) | (n13337 & n16323) | (n13338 & n16323);
  assign n16412 = (n16230 & n16410) | (n16230 & n16411) | (n16410 & n16411);
  assign n7528 = ~n16409 & n16412;
  assign n7529 = x73 & x85;
  assign n7530 = n7528 & n7529;
  assign n7531 = n7528 | n7529;
  assign n7532 = ~n7530 & n7531;
  assign n16384 = n7301 | n7303;
  assign n16385 = (n7301 & n13224) | (n7301 & n16384) | (n13224 & n16384);
  assign n16413 = n7532 & n16385;
  assign n16382 = n7080 | n7301;
  assign n16383 = (n7301 & n7303) | (n7301 & n16382) | (n7303 & n16382);
  assign n16414 = n7532 & n16383;
  assign n16415 = (n13130 & n16413) | (n13130 & n16414) | (n16413 & n16414);
  assign n16416 = n7532 | n16385;
  assign n16417 = n7532 | n16383;
  assign n16418 = (n13130 & n16416) | (n13130 & n16417) | (n16416 & n16417);
  assign n7535 = ~n16415 & n16418;
  assign n7536 = x72 & x86;
  assign n7537 = n7535 & n7536;
  assign n7538 = n7535 | n7536;
  assign n7539 = ~n7537 & n7538;
  assign n13340 = n7308 & n7539;
  assign n13341 = (n7539 & n13258) | (n7539 & n13340) | (n13258 & n13340);
  assign n13342 = n7308 | n7539;
  assign n13343 = n13258 | n13342;
  assign n7542 = ~n13341 & n13343;
  assign n7543 = x71 & x87;
  assign n7544 = n7542 & n7543;
  assign n7545 = n7542 | n7543;
  assign n7546 = ~n7544 & n7545;
  assign n7547 = n16381 & n7546;
  assign n7548 = n16381 | n7546;
  assign n7549 = ~n7547 & n7548;
  assign n7550 = x70 & x88;
  assign n7551 = n7549 & n7550;
  assign n7552 = n7549 | n7550;
  assign n7553 = ~n7551 & n7552;
  assign n13309 = n7322 | n7324;
  assign n13344 = n7553 & n13309;
  assign n13345 = n7322 & n7553;
  assign n13346 = (n16319 & n13344) | (n16319 & n13345) | (n13344 & n13345);
  assign n13347 = n7553 | n13309;
  assign n13348 = n7322 | n7553;
  assign n13349 = (n16319 & n13347) | (n16319 & n13348) | (n13347 & n13348);
  assign n7556 = ~n13346 & n13349;
  assign n7557 = x69 & x89;
  assign n7558 = n7556 & n7557;
  assign n7559 = n7556 | n7557;
  assign n7560 = ~n7558 & n7559;
  assign n13350 = n7329 & n7560;
  assign n16419 = (n7560 & n13267) | (n7560 & n13350) | (n13267 & n13350);
  assign n16420 = (n7560 & n13266) | (n7560 & n13350) | (n13266 & n13350);
  assign n16421 = (n16270 & n16419) | (n16270 & n16420) | (n16419 & n16420);
  assign n13352 = n7329 | n7560;
  assign n16422 = n13267 | n13352;
  assign n16423 = n13266 | n13352;
  assign n16424 = (n16270 & n16422) | (n16270 & n16423) | (n16422 & n16423);
  assign n7563 = ~n16421 & n16424;
  assign n7564 = x68 & x90;
  assign n7565 = n7563 & n7564;
  assign n7566 = n7563 | n7564;
  assign n7567 = ~n7565 & n7566;
  assign n13307 = n7336 | n7338;
  assign n16425 = n7567 & n13307;
  assign n16375 = n7115 | n7336;
  assign n16376 = (n7336 & n7338) | (n7336 & n16375) | (n7338 & n16375);
  assign n16426 = n7567 & n16376;
  assign n16427 = (n16299 & n16425) | (n16299 & n16426) | (n16425 & n16426);
  assign n16428 = n7567 | n13307;
  assign n16429 = n7567 | n16376;
  assign n16430 = (n16299 & n16428) | (n16299 & n16429) | (n16428 & n16429);
  assign n7570 = ~n16427 & n16430;
  assign n7571 = x67 & x91;
  assign n7572 = n7570 & n7571;
  assign n7573 = n7570 | n7571;
  assign n7574 = ~n7572 & n7573;
  assign n13354 = n7343 & n7574;
  assign n16431 = (n7574 & n13276) | (n7574 & n13354) | (n13276 & n13354);
  assign n16432 = (n7345 & n7574) | (n7345 & n13354) | (n7574 & n13354);
  assign n16433 = (n13181 & n16431) | (n13181 & n16432) | (n16431 & n16432);
  assign n13356 = n7343 | n7574;
  assign n16434 = n13276 | n13356;
  assign n16435 = n7345 | n13356;
  assign n16436 = (n13181 & n16434) | (n13181 & n16435) | (n16434 & n16435);
  assign n7577 = ~n16433 & n16436;
  assign n7578 = x66 & x92;
  assign n7579 = n7577 & n7578;
  assign n7580 = n7577 | n7578;
  assign n7581 = ~n7579 & n7580;
  assign n13358 = n7350 & n7581;
  assign n13359 = (n7581 & n13282) | (n7581 & n13358) | (n13282 & n13358);
  assign n13360 = n7350 | n7581;
  assign n13361 = n13282 | n13360;
  assign n7584 = ~n13359 & n13361;
  assign n7585 = x65 & x93;
  assign n7586 = n7584 & n7585;
  assign n7587 = n7584 | n7585;
  assign n7588 = ~n7586 & n7587;
  assign n13304 = n7357 | n7359;
  assign n13362 = n7588 & n13304;
  assign n13363 = n7357 & n7588;
  assign n13364 = (n13214 & n13362) | (n13214 & n13363) | (n13362 & n13363);
  assign n13365 = n7588 | n13304;
  assign n13366 = n7357 | n7588;
  assign n13367 = (n13214 & n13365) | (n13214 & n13366) | (n13365 & n13366);
  assign n7591 = ~n13364 & n13367;
  assign n7592 = x64 & x94;
  assign n7593 = n7591 & n7592;
  assign n7594 = n7591 | n7592;
  assign n7595 = ~n7593 & n7594;
  assign n13302 = n7364 | n7366;
  assign n16437 = n7595 & n13302;
  assign n16438 = n7364 & n7595;
  assign n16439 = (n13212 & n16437) | (n13212 & n16438) | (n16437 & n16438);
  assign n16440 = n7595 | n13302;
  assign n16441 = n7364 | n7595;
  assign n16442 = (n13212 & n16440) | (n13212 & n16441) | (n16440 & n16441);
  assign n7598 = ~n16439 & n16442;
  assign n7599 = x63 & x95;
  assign n7600 = n7598 & n7599;
  assign n7601 = n7598 | n7599;
  assign n7602 = ~n7600 & n7601;
  assign n13300 = n7371 | n7373;
  assign n16443 = n7602 & n13300;
  assign n16444 = n7371 & n7602;
  assign n16445 = (n13210 & n16443) | (n13210 & n16444) | (n16443 & n16444);
  assign n16446 = n7602 | n13300;
  assign n16447 = n7371 | n7602;
  assign n16448 = (n13210 & n16446) | (n13210 & n16447) | (n16446 & n16447);
  assign n7605 = ~n16445 & n16448;
  assign n7606 = x62 & x96;
  assign n7607 = n7605 & n7606;
  assign n7608 = n7605 | n7606;
  assign n7609 = ~n7607 & n7608;
  assign n7610 = n13299 & n7609;
  assign n7611 = n13299 | n7609;
  assign n7612 = ~n7610 & n7611;
  assign n7613 = x61 & x97;
  assign n7614 = n7612 & n7613;
  assign n7615 = n7612 | n7613;
  assign n7616 = ~n7614 & n7615;
  assign n7617 = n13297 & n7616;
  assign n7618 = n13297 | n7616;
  assign n7619 = ~n7617 & n7618;
  assign n7620 = x60 & x98;
  assign n7621 = n7619 & n7620;
  assign n7622 = n7619 | n7620;
  assign n7623 = ~n7621 & n7622;
  assign n7624 = n13295 & n7623;
  assign n7625 = n13295 | n7623;
  assign n7626 = ~n7624 & n7625;
  assign n7627 = x59 & x99;
  assign n7628 = n7626 & n7627;
  assign n7629 = n7626 | n7627;
  assign n7630 = ~n7628 & n7629;
  assign n7631 = n13293 & n7630;
  assign n7632 = n13293 | n7630;
  assign n7633 = ~n7631 & n7632;
  assign n7634 = x58 & x100;
  assign n7635 = n7633 & n7634;
  assign n7636 = n7633 | n7634;
  assign n7637 = ~n7635 & n7636;
  assign n7638 = n13291 & n7637;
  assign n7639 = n13291 | n7637;
  assign n7640 = ~n7638 & n7639;
  assign n7641 = x57 & x101;
  assign n7642 = n7640 & n7641;
  assign n7643 = n7640 | n7641;
  assign n7644 = ~n7642 & n7643;
  assign n7645 = n13289 & n7644;
  assign n7646 = n13289 | n7644;
  assign n7647 = ~n7645 & n7646;
  assign n7648 = x56 & x102;
  assign n7649 = n7647 & n7648;
  assign n7650 = n7647 | n7648;
  assign n7651 = ~n7649 & n7650;
  assign n7652 = n7478 & n7651;
  assign n7653 = n7478 | n7651;
  assign n7654 = ~n7652 & n7653;
  assign n7655 = x55 & x103;
  assign n7656 = n7654 & n7655;
  assign n7657 = n7654 | n7655;
  assign n7658 = ~n7656 & n7657;
  assign n7659 = n7477 & n7658;
  assign n7660 = n7477 | n7658;
  assign n7661 = ~n7659 & n7660;
  assign n7662 = x54 & x104;
  assign n7663 = n7661 & n7662;
  assign n7664 = n7661 | n7662;
  assign n7665 = ~n7663 & n7664;
  assign n7666 = n7476 & n7665;
  assign n7667 = n7476 | n7665;
  assign n7668 = ~n7666 & n7667;
  assign n7669 = x53 & x105;
  assign n7670 = n7668 & n7669;
  assign n7671 = n7668 | n7669;
  assign n7672 = ~n7670 & n7671;
  assign n7673 = n7475 & n7672;
  assign n7674 = n7475 | n7672;
  assign n7675 = ~n7673 & n7674;
  assign n7676 = x52 & x106;
  assign n7677 = n7675 & n7676;
  assign n7678 = n7675 | n7676;
  assign n7679 = ~n7677 & n7678;
  assign n7680 = n7474 & n7679;
  assign n7681 = n7474 | n7679;
  assign n7682 = ~n7680 & n7681;
  assign n7683 = x51 & x107;
  assign n7684 = n7682 & n7683;
  assign n7685 = n7682 | n7683;
  assign n7686 = ~n7684 & n7685;
  assign n7687 = n16374 & n7686;
  assign n7688 = n16374 | n7686;
  assign n7689 = ~n7687 & n7688;
  assign n7690 = x50 & x108;
  assign n7691 = n7689 & n7690;
  assign n7692 = n7689 | n7690;
  assign n7693 = ~n7691 & n7692;
  assign n7694 = n13287 & n7693;
  assign n7695 = n13287 | n7693;
  assign n7696 = ~n7694 & n7695;
  assign n7697 = x49 & x109;
  assign n7698 = n7696 & n7697;
  assign n7699 = n7696 | n7697;
  assign n7700 = ~n7698 & n7699;
  assign n7701 = n7469 & n7700;
  assign n7702 = n7469 | n7700;
  assign n7703 = ~n7701 & n7702;
  assign n7704 = x48 & x110;
  assign n7705 = n7703 & n7704;
  assign n7706 = n7703 | n7704;
  assign n7707 = ~n7705 & n7706;
  assign n17754 = n7468 | n7697;
  assign n17755 = (n7467 & n7697) | (n7467 & n17754) | (n7697 & n17754);
  assign n16450 = (n7469 & n7696) | (n7469 & n17755) | (n7696 & n17755);
  assign n13369 = (n7698 & n7700) | (n7698 & n16450) | (n7700 & n16450);
  assign n13370 = n7691 | n13287;
  assign n13371 = (n7691 & n7693) | (n7691 & n13370) | (n7693 & n13370);
  assign n16451 = n7684 | n16374;
  assign n16452 = (n7684 & n7686) | (n7684 & n16451) | (n7686 & n16451);
  assign n7711 = n7677 | n7680;
  assign n7712 = n7670 | n7673;
  assign n7713 = n7663 | n7666;
  assign n7714 = n7656 | n7659;
  assign n13372 = n7649 | n7651;
  assign n13373 = (n7478 & n7649) | (n7478 & n13372) | (n7649 & n13372);
  assign n13374 = n7642 | n7644;
  assign n13375 = (n7642 & n13289) | (n7642 & n13374) | (n13289 & n13374);
  assign n13376 = n7635 | n7637;
  assign n13377 = (n7635 & n13291) | (n7635 & n13376) | (n13291 & n13376);
  assign n13378 = n7628 | n7630;
  assign n13379 = (n7628 & n13293) | (n7628 & n13378) | (n13293 & n13378);
  assign n13380 = n7621 | n7623;
  assign n13381 = (n7621 & n13295) | (n7621 & n13380) | (n13295 & n13380);
  assign n13382 = n7614 | n7616;
  assign n13383 = (n7614 & n13297) | (n7614 & n13382) | (n13297 & n13382);
  assign n13301 = (n7371 & n13210) | (n7371 & n13300) | (n13210 & n13300);
  assign n13303 = (n7364 & n13212) | (n7364 & n13302) | (n13212 & n13302);
  assign n13393 = n7558 | n7560;
  assign n16453 = n7329 | n7558;
  assign n16454 = (n7558 & n7560) | (n7558 & n16453) | (n7560 & n16453);
  assign n16455 = (n13267 & n13393) | (n13267 & n16454) | (n13393 & n16454);
  assign n16456 = (n13266 & n13393) | (n13266 & n16454) | (n13393 & n16454);
  assign n16457 = (n16270 & n16455) | (n16270 & n16456) | (n16455 & n16456);
  assign n13228 = (n16230 & n16321) | (n16230 & n16323) | (n16321 & n16323);
  assign n7737 = x79 & x80;
  assign n7738 = x78 & x81;
  assign n7739 = n7737 & n7738;
  assign n7740 = n7737 | n7738;
  assign n7741 = ~n7739 & n7740;
  assign n13411 = n7502 | n7504;
  assign n13413 = n7741 & n13411;
  assign n13414 = n7502 & n7741;
  assign n17756 = (n7273 & n13413) | (n7273 & n13414) | (n13413 & n13414);
  assign n17757 = n13413 | n13414;
  assign n17758 = (n16332 & n17756) | (n16332 & n17757) | (n17756 & n17757);
  assign n17759 = (n13413 & n13414) | (n13413 & n16387) | (n13414 & n16387);
  assign n17760 = (n13413 & n13414) | (n13413 & n17740) | (n13414 & n17740);
  assign n17761 = (n16282 & n17759) | (n16282 & n17760) | (n17759 & n17760);
  assign n16462 = (n16123 & n17758) | (n16123 & n17761) | (n17758 & n17761);
  assign n13416 = n7741 | n13411;
  assign n13417 = n7502 | n7741;
  assign n17762 = (n7273 & n13416) | (n7273 & n13417) | (n13416 & n13417);
  assign n17763 = n13416 | n13417;
  assign n17764 = (n16332 & n17762) | (n16332 & n17763) | (n17762 & n17763);
  assign n17765 = (n13416 & n13417) | (n13416 & n16387) | (n13417 & n16387);
  assign n17766 = (n13416 & n13417) | (n13416 & n17740) | (n13417 & n17740);
  assign n17767 = (n16282 & n17765) | (n16282 & n17766) | (n17765 & n17766);
  assign n16465 = (n16123 & n17764) | (n16123 & n17767) | (n17764 & n17767);
  assign n7744 = ~n16462 & n16465;
  assign n7745 = x77 & x82;
  assign n7746 = n7744 & n7745;
  assign n7747 = n7744 | n7745;
  assign n7748 = ~n7746 & n7747;
  assign n16466 = n7509 | n7511;
  assign n16467 = (n7509 & n13319) | (n7509 & n16466) | (n13319 & n16466);
  assign n13419 = n7748 & n16467;
  assign n16468 = n7280 | n7509;
  assign n16469 = (n7509 & n7511) | (n7509 & n16468) | (n7511 & n16468);
  assign n13420 = n7748 & n16469;
  assign n16470 = (n13419 & n13420) | (n13419 & n16325) | (n13420 & n16325);
  assign n16471 = (n13419 & n13420) | (n13419 & n16326) | (n13420 & n16326);
  assign n16472 = (n16182 & n16470) | (n16182 & n16471) | (n16470 & n16471);
  assign n13422 = n7748 | n16467;
  assign n13423 = n7748 | n16469;
  assign n16473 = (n13422 & n13423) | (n13422 & n16325) | (n13423 & n16325);
  assign n16474 = (n13422 & n13423) | (n13422 & n16326) | (n13423 & n16326);
  assign n16475 = (n16182 & n16473) | (n16182 & n16474) | (n16473 & n16474);
  assign n7751 = ~n16472 & n16475;
  assign n7752 = x76 & x83;
  assign n7753 = n7751 & n7752;
  assign n7754 = n7751 | n7752;
  assign n7755 = ~n7753 & n7754;
  assign n16476 = n7287 | n7516;
  assign n16477 = (n7516 & n7518) | (n7516 & n16476) | (n7518 & n16476);
  assign n13425 = n7755 & n16477;
  assign n13406 = n7516 | n7518;
  assign n13426 = n7755 & n13406;
  assign n16478 = (n13244 & n13425) | (n13244 & n13426) | (n13425 & n13426);
  assign n16479 = (n13245 & n13425) | (n13245 & n13426) | (n13425 & n13426);
  assign n16480 = (n16233 & n16478) | (n16233 & n16479) | (n16478 & n16479);
  assign n13428 = n7755 | n16477;
  assign n13429 = n7755 | n13406;
  assign n16481 = (n13244 & n13428) | (n13244 & n13429) | (n13428 & n13429);
  assign n16482 = (n13245 & n13428) | (n13245 & n13429) | (n13428 & n13429);
  assign n16483 = (n16233 & n16481) | (n16233 & n16482) | (n16481 & n16482);
  assign n7758 = ~n16480 & n16483;
  assign n7759 = x75 & x84;
  assign n7760 = n7758 & n7759;
  assign n7761 = n7758 | n7759;
  assign n7762 = ~n7760 & n7761;
  assign n16484 = n7523 | n7525;
  assign n16485 = (n7523 & n13317) | (n7523 & n16484) | (n13317 & n16484);
  assign n13431 = n7762 & n16485;
  assign n16486 = n7294 | n7523;
  assign n16487 = (n7523 & n7525) | (n7523 & n16486) | (n7525 & n16486);
  assign n13432 = n7762 & n16487;
  assign n13433 = (n13228 & n13431) | (n13228 & n13432) | (n13431 & n13432);
  assign n13434 = n7762 | n16485;
  assign n13435 = n7762 | n16487;
  assign n13436 = (n13228 & n13434) | (n13228 & n13435) | (n13434 & n13435);
  assign n7765 = ~n13433 & n13436;
  assign n7766 = x74 & x85;
  assign n7767 = n7765 & n7766;
  assign n7768 = n7765 | n7766;
  assign n7769 = ~n7767 & n7768;
  assign n13400 = n7530 | n7532;
  assign n13437 = n7769 & n13400;
  assign n13438 = n7530 & n7769;
  assign n16488 = (n13437 & n13438) | (n13437 & n16385) | (n13438 & n16385);
  assign n16489 = (n13437 & n13438) | (n13437 & n16383) | (n13438 & n16383);
  assign n16490 = (n13130 & n16488) | (n13130 & n16489) | (n16488 & n16489);
  assign n13440 = n7769 | n13400;
  assign n13441 = n7530 | n7769;
  assign n16491 = (n13440 & n13441) | (n13440 & n16385) | (n13441 & n16385);
  assign n16492 = (n13440 & n13441) | (n13440 & n16383) | (n13441 & n16383);
  assign n16493 = (n13130 & n16491) | (n13130 & n16492) | (n16491 & n16492);
  assign n7772 = ~n16490 & n16493;
  assign n7773 = x73 & x86;
  assign n7774 = n7772 & n7773;
  assign n7775 = n7772 | n7773;
  assign n7776 = ~n7774 & n7775;
  assign n13398 = n7537 | n7539;
  assign n16494 = n7776 & n13398;
  assign n16458 = n7308 | n7537;
  assign n16459 = (n7537 & n7539) | (n7537 & n16458) | (n7539 & n16458);
  assign n16495 = n7776 & n16459;
  assign n16496 = (n13258 & n16494) | (n13258 & n16495) | (n16494 & n16495);
  assign n16497 = n7776 | n13398;
  assign n16498 = n7776 | n16459;
  assign n16499 = (n13258 & n16497) | (n13258 & n16498) | (n16497 & n16498);
  assign n7779 = ~n16496 & n16499;
  assign n7780 = x72 & x87;
  assign n7781 = n7779 & n7780;
  assign n7782 = n7779 | n7780;
  assign n7783 = ~n7781 & n7782;
  assign n13395 = n7544 | n7546;
  assign n13443 = n7783 & n13395;
  assign n13444 = n7544 & n7783;
  assign n13445 = (n16381 & n13443) | (n16381 & n13444) | (n13443 & n13444);
  assign n13446 = n7783 | n13395;
  assign n13447 = n7544 | n7783;
  assign n13448 = (n16381 & n13446) | (n16381 & n13447) | (n13446 & n13447);
  assign n7786 = ~n13445 & n13448;
  assign n7787 = x71 & x88;
  assign n7788 = n7786 & n7787;
  assign n7789 = n7786 | n7787;
  assign n7790 = ~n7788 & n7789;
  assign n13449 = n7551 & n7790;
  assign n16500 = (n7790 & n13345) | (n7790 & n13449) | (n13345 & n13449);
  assign n16501 = (n7790 & n13344) | (n7790 & n13449) | (n13344 & n13449);
  assign n16502 = (n16319 & n16500) | (n16319 & n16501) | (n16500 & n16501);
  assign n13451 = n7551 | n7790;
  assign n16503 = n13345 | n13451;
  assign n16504 = n13344 | n13451;
  assign n16505 = (n16319 & n16503) | (n16319 & n16504) | (n16503 & n16504);
  assign n7793 = ~n16502 & n16505;
  assign n7794 = x70 & x89;
  assign n7795 = n7793 & n7794;
  assign n7796 = n7793 | n7794;
  assign n7797 = ~n7795 & n7796;
  assign n7798 = n16457 & n7797;
  assign n7799 = n16457 | n7797;
  assign n7800 = ~n7798 & n7799;
  assign n7801 = x69 & x90;
  assign n7802 = n7800 & n7801;
  assign n7803 = n7800 | n7801;
  assign n7804 = ~n7802 & n7803;
  assign n13390 = n7565 | n7567;
  assign n13453 = n7804 & n13390;
  assign n13454 = n7565 & n7804;
  assign n16506 = (n13307 & n13453) | (n13307 & n13454) | (n13453 & n13454);
  assign n16507 = (n13453 & n13454) | (n13453 & n16376) | (n13454 & n16376);
  assign n16508 = (n16299 & n16506) | (n16299 & n16507) | (n16506 & n16507);
  assign n13456 = n7804 | n13390;
  assign n13457 = n7565 | n7804;
  assign n16509 = (n13307 & n13456) | (n13307 & n13457) | (n13456 & n13457);
  assign n16510 = (n13456 & n13457) | (n13456 & n16376) | (n13457 & n16376);
  assign n16511 = (n16299 & n16509) | (n16299 & n16510) | (n16509 & n16510);
  assign n7807 = ~n16508 & n16511;
  assign n7808 = x68 & x91;
  assign n7809 = n7807 & n7808;
  assign n7810 = n7807 | n7808;
  assign n7811 = ~n7809 & n7810;
  assign n13459 = n7572 & n7811;
  assign n13460 = (n7811 & n16433) | (n7811 & n13459) | (n16433 & n13459);
  assign n13461 = n7572 | n7811;
  assign n13462 = n16433 | n13461;
  assign n7814 = ~n13460 & n13462;
  assign n7815 = x67 & x92;
  assign n7816 = n7814 & n7815;
  assign n7817 = n7814 | n7815;
  assign n7818 = ~n7816 & n7817;
  assign n13463 = n7579 & n7818;
  assign n13464 = (n7818 & n13359) | (n7818 & n13463) | (n13359 & n13463);
  assign n13465 = n7579 | n7818;
  assign n13466 = n13359 | n13465;
  assign n7821 = ~n13464 & n13466;
  assign n7822 = x66 & x93;
  assign n7823 = n7821 & n7822;
  assign n7824 = n7821 | n7822;
  assign n7825 = ~n7823 & n7824;
  assign n13467 = n7586 & n7825;
  assign n13468 = (n7825 & n13364) | (n7825 & n13467) | (n13364 & n13467);
  assign n13469 = n7586 | n7825;
  assign n13470 = n13364 | n13469;
  assign n7828 = ~n13468 & n13470;
  assign n7829 = x65 & x94;
  assign n7830 = n7828 & n7829;
  assign n7831 = n7828 | n7829;
  assign n7832 = ~n7830 & n7831;
  assign n13388 = n7593 | n7595;
  assign n13471 = n7832 & n13388;
  assign n13472 = n7593 & n7832;
  assign n13473 = (n13303 & n13471) | (n13303 & n13472) | (n13471 & n13472);
  assign n13474 = n7832 | n13388;
  assign n13475 = n7593 | n7832;
  assign n13476 = (n13303 & n13474) | (n13303 & n13475) | (n13474 & n13475);
  assign n7835 = ~n13473 & n13476;
  assign n7836 = x64 & x95;
  assign n7837 = n7835 & n7836;
  assign n7838 = n7835 | n7836;
  assign n7839 = ~n7837 & n7838;
  assign n13386 = n7600 | n7602;
  assign n16512 = n7839 & n13386;
  assign n16513 = n7600 & n7839;
  assign n16514 = (n13301 & n16512) | (n13301 & n16513) | (n16512 & n16513);
  assign n16515 = n7839 | n13386;
  assign n16516 = n7600 | n7839;
  assign n16517 = (n13301 & n16515) | (n13301 & n16516) | (n16515 & n16516);
  assign n7842 = ~n16514 & n16517;
  assign n7843 = x63 & x96;
  assign n7844 = n7842 & n7843;
  assign n7845 = n7842 | n7843;
  assign n7846 = ~n7844 & n7845;
  assign n13384 = n7607 | n7609;
  assign n16518 = n7846 & n13384;
  assign n16519 = n7607 & n7846;
  assign n16520 = (n13299 & n16518) | (n13299 & n16519) | (n16518 & n16519);
  assign n16521 = n7846 | n13384;
  assign n16522 = n7607 | n7846;
  assign n16523 = (n13299 & n16521) | (n13299 & n16522) | (n16521 & n16522);
  assign n7849 = ~n16520 & n16523;
  assign n7850 = x62 & x97;
  assign n7851 = n7849 & n7850;
  assign n7852 = n7849 | n7850;
  assign n7853 = ~n7851 & n7852;
  assign n7854 = n13383 & n7853;
  assign n7855 = n13383 | n7853;
  assign n7856 = ~n7854 & n7855;
  assign n7857 = x61 & x98;
  assign n7858 = n7856 & n7857;
  assign n7859 = n7856 | n7857;
  assign n7860 = ~n7858 & n7859;
  assign n7861 = n13381 & n7860;
  assign n7862 = n13381 | n7860;
  assign n7863 = ~n7861 & n7862;
  assign n7864 = x60 & x99;
  assign n7865 = n7863 & n7864;
  assign n7866 = n7863 | n7864;
  assign n7867 = ~n7865 & n7866;
  assign n7868 = n13379 & n7867;
  assign n7869 = n13379 | n7867;
  assign n7870 = ~n7868 & n7869;
  assign n7871 = x59 & x100;
  assign n7872 = n7870 & n7871;
  assign n7873 = n7870 | n7871;
  assign n7874 = ~n7872 & n7873;
  assign n7875 = n13377 & n7874;
  assign n7876 = n13377 | n7874;
  assign n7877 = ~n7875 & n7876;
  assign n7878 = x58 & x101;
  assign n7879 = n7877 & n7878;
  assign n7880 = n7877 | n7878;
  assign n7881 = ~n7879 & n7880;
  assign n7882 = n13375 & n7881;
  assign n7883 = n13375 | n7881;
  assign n7884 = ~n7882 & n7883;
  assign n7885 = x57 & x102;
  assign n7886 = n7884 & n7885;
  assign n7887 = n7884 | n7885;
  assign n7888 = ~n7886 & n7887;
  assign n7889 = n13373 & n7888;
  assign n7890 = n13373 | n7888;
  assign n7891 = ~n7889 & n7890;
  assign n7892 = x56 & x103;
  assign n7893 = n7891 & n7892;
  assign n7894 = n7891 | n7892;
  assign n7895 = ~n7893 & n7894;
  assign n7896 = n7714 & n7895;
  assign n7897 = n7714 | n7895;
  assign n7898 = ~n7896 & n7897;
  assign n7899 = x55 & x104;
  assign n7900 = n7898 & n7899;
  assign n7901 = n7898 | n7899;
  assign n7902 = ~n7900 & n7901;
  assign n7903 = n7713 & n7902;
  assign n7904 = n7713 | n7902;
  assign n7905 = ~n7903 & n7904;
  assign n7906 = x54 & x105;
  assign n7907 = n7905 & n7906;
  assign n7908 = n7905 | n7906;
  assign n7909 = ~n7907 & n7908;
  assign n7910 = n7712 & n7909;
  assign n7911 = n7712 | n7909;
  assign n7912 = ~n7910 & n7911;
  assign n7913 = x53 & x106;
  assign n7914 = n7912 & n7913;
  assign n7915 = n7912 | n7913;
  assign n7916 = ~n7914 & n7915;
  assign n7917 = n7711 & n7916;
  assign n7918 = n7711 | n7916;
  assign n7919 = ~n7917 & n7918;
  assign n7920 = x52 & x107;
  assign n7921 = n7919 & n7920;
  assign n7922 = n7919 | n7920;
  assign n7923 = ~n7921 & n7922;
  assign n7924 = n16452 & n7923;
  assign n7925 = n16452 | n7923;
  assign n7926 = ~n7924 & n7925;
  assign n7927 = x51 & x108;
  assign n7928 = n7926 & n7927;
  assign n7929 = n7926 | n7927;
  assign n7930 = ~n7928 & n7929;
  assign n7931 = n13371 & n7930;
  assign n7932 = n13371 | n7930;
  assign n7933 = ~n7931 & n7932;
  assign n7934 = x50 & x109;
  assign n7935 = n7933 & n7934;
  assign n7936 = n7933 | n7934;
  assign n7937 = ~n7935 & n7936;
  assign n7938 = n13369 & n7937;
  assign n7939 = n13369 | n7937;
  assign n7940 = ~n7938 & n7939;
  assign n7941 = x49 & x110;
  assign n7942 = n7940 & n7941;
  assign n7943 = n7940 | n7941;
  assign n7944 = ~n7942 & n7943;
  assign n7945 = n7705 & n7944;
  assign n7946 = n7705 | n7944;
  assign n7947 = ~n7945 & n7946;
  assign n7948 = x48 & x111;
  assign n7949 = n7947 & n7948;
  assign n7950 = n7947 | n7948;
  assign n7951 = ~n7949 & n7950;
  assign n17768 = n7704 | n7941;
  assign n17769 = (n7703 & n7941) | (n7703 & n17768) | (n7941 & n17768);
  assign n16525 = (n7705 & n7940) | (n7705 & n17769) | (n7940 & n17769);
  assign n13478 = (n7942 & n7944) | (n7942 & n16525) | (n7944 & n16525);
  assign n13479 = n7935 | n13369;
  assign n13480 = (n7935 & n7937) | (n7935 & n13479) | (n7937 & n13479);
  assign n13481 = n7928 | n13371;
  assign n13482 = (n7928 & n7930) | (n7928 & n13481) | (n7930 & n13481);
  assign n16526 = n7921 | n16452;
  assign n16527 = (n7921 & n7923) | (n7921 & n16526) | (n7923 & n16526);
  assign n7956 = n7914 | n7917;
  assign n7957 = n7907 | n7910;
  assign n7958 = n7900 | n7903;
  assign n13483 = n7893 | n7895;
  assign n13484 = (n7714 & n7893) | (n7714 & n13483) | (n7893 & n13483);
  assign n13485 = n7886 | n7888;
  assign n13486 = (n7886 & n13373) | (n7886 & n13485) | (n13373 & n13485);
  assign n13487 = n7879 | n7881;
  assign n13488 = (n7879 & n13375) | (n7879 & n13487) | (n13375 & n13487);
  assign n13489 = n7872 | n7874;
  assign n13490 = (n7872 & n13377) | (n7872 & n13489) | (n13377 & n13489);
  assign n13491 = n7865 | n7867;
  assign n13492 = (n7865 & n13379) | (n7865 & n13491) | (n13379 & n13491);
  assign n13493 = n7858 | n7860;
  assign n13494 = (n7858 & n13381) | (n7858 & n13493) | (n13381 & n13493);
  assign n13385 = (n7607 & n13299) | (n7607 & n13384) | (n13299 & n13384);
  assign n13387 = (n7600 & n13301) | (n7600 & n13386) | (n13301 & n13386);
  assign n13507 = n7788 | n7790;
  assign n16530 = n7551 | n7788;
  assign n16531 = (n7788 & n7790) | (n7788 & n16530) | (n7790 & n16530);
  assign n16532 = (n13345 & n13507) | (n13345 & n16531) | (n13507 & n16531);
  assign n16533 = (n13344 & n13507) | (n13344 & n16531) | (n13507 & n16531);
  assign n16534 = (n16319 & n16532) | (n16319 & n16533) | (n16532 & n16533);
  assign n13316 = (n13130 & n16383) | (n13130 & n16385) | (n16383 & n16385);
  assign n16537 = n7753 | n7755;
  assign n16538 = (n7753 & n16477) | (n7753 & n16537) | (n16477 & n16537);
  assign n16539 = (n7753 & n13406) | (n7753 & n16537) | (n13406 & n16537);
  assign n16540 = (n13244 & n16538) | (n13244 & n16539) | (n16538 & n16539);
  assign n16541 = (n13245 & n16538) | (n13245 & n16539) | (n16538 & n16539);
  assign n16542 = (n16233 & n16540) | (n16233 & n16541) | (n16540 & n16541);
  assign n13322 = n7273 | n16332;
  assign n7982 = x79 & x81;
  assign n16543 = n7739 | n7741;
  assign n16544 = (n7739 & n13411) | (n7739 & n16543) | (n13411 & n16543);
  assign n13523 = n7982 & n16544;
  assign n16545 = n7502 | n7739;
  assign n16546 = (n7739 & n7741) | (n7739 & n16545) | (n7741 & n16545);
  assign n13524 = n7982 & n16546;
  assign n16547 = (n13322 & n13523) | (n13322 & n13524) | (n13523 & n13524);
  assign n16388 = (n16282 & n17740) | (n16282 & n16387) | (n17740 & n16387);
  assign n16548 = (n13523 & n13524) | (n13523 & n16388) | (n13524 & n16388);
  assign n16549 = (n16123 & n16547) | (n16123 & n16548) | (n16547 & n16548);
  assign n13526 = n7982 | n16544;
  assign n13527 = n7982 | n16546;
  assign n16550 = (n13322 & n13526) | (n13322 & n13527) | (n13526 & n13527);
  assign n16551 = (n13526 & n13527) | (n13526 & n16388) | (n13527 & n16388);
  assign n16552 = (n16123 & n16550) | (n16123 & n16551) | (n16550 & n16551);
  assign n7985 = ~n16549 & n16552;
  assign n7986 = x78 & x82;
  assign n7987 = n7985 & n7986;
  assign n7988 = n7985 | n7986;
  assign n7989 = ~n7987 & n7988;
  assign n16553 = n7746 | n7748;
  assign n16558 = (n7746 & n16469) | (n7746 & n16553) | (n16469 & n16553);
  assign n13530 = n7989 & n16558;
  assign n16555 = n7989 & n16553;
  assign n16556 = n7746 & n7989;
  assign n16557 = (n16467 & n16555) | (n16467 & n16556) | (n16555 & n16556);
  assign n16559 = (n13530 & n16325) | (n13530 & n16557) | (n16325 & n16557);
  assign n16560 = (n13530 & n16326) | (n13530 & n16557) | (n16326 & n16557);
  assign n16561 = (n16182 & n16559) | (n16182 & n16560) | (n16559 & n16560);
  assign n13533 = n7989 | n16558;
  assign n16562 = n7989 | n16553;
  assign n16563 = n7746 | n7989;
  assign n16564 = (n16467 & n16562) | (n16467 & n16563) | (n16562 & n16563);
  assign n16565 = (n13533 & n16325) | (n13533 & n16564) | (n16325 & n16564);
  assign n16566 = (n13533 & n16326) | (n13533 & n16564) | (n16326 & n16564);
  assign n16567 = (n16182 & n16565) | (n16182 & n16566) | (n16565 & n16566);
  assign n7992 = ~n16561 & n16567;
  assign n7993 = x77 & x83;
  assign n7994 = n7992 & n7993;
  assign n7995 = n7992 | n7993;
  assign n7996 = ~n7994 & n7995;
  assign n7997 = n16542 & n7996;
  assign n7998 = n16542 | n7996;
  assign n7999 = ~n7997 & n7998;
  assign n8000 = x76 & x84;
  assign n8001 = n7999 & n8000;
  assign n8002 = n7999 | n8000;
  assign n8003 = ~n8001 & n8002;
  assign n13535 = n7760 & n8003;
  assign n16568 = (n8003 & n13431) | (n8003 & n13535) | (n13431 & n13535);
  assign n16569 = (n8003 & n13432) | (n8003 & n13535) | (n13432 & n13535);
  assign n16570 = (n13228 & n16568) | (n13228 & n16569) | (n16568 & n16569);
  assign n13537 = n7760 | n8003;
  assign n16571 = n13431 | n13537;
  assign n16572 = n13432 | n13537;
  assign n16573 = (n13228 & n16571) | (n13228 & n16572) | (n16571 & n16572);
  assign n8006 = ~n16570 & n16573;
  assign n8007 = x75 & x85;
  assign n8008 = n8006 & n8007;
  assign n8009 = n8006 | n8007;
  assign n8010 = ~n8008 & n8009;
  assign n17770 = n7767 & n8010;
  assign n17771 = (n8010 & n13437) | (n8010 & n17770) | (n13437 & n17770);
  assign n16535 = n7530 | n7767;
  assign n16536 = (n7767 & n7769) | (n7767 & n16535) | (n7769 & n16535);
  assign n16575 = n8010 & n16536;
  assign n16576 = (n13316 & n17771) | (n13316 & n16575) | (n17771 & n16575);
  assign n17772 = n7767 | n8010;
  assign n17773 = n13437 | n17772;
  assign n16578 = n8010 | n16536;
  assign n16579 = (n13316 & n17773) | (n13316 & n16578) | (n17773 & n16578);
  assign n8013 = ~n16576 & n16579;
  assign n8014 = x74 & x86;
  assign n8015 = n8013 & n8014;
  assign n8016 = n8013 | n8014;
  assign n8017 = ~n8015 & n8016;
  assign n13509 = n7774 | n7776;
  assign n13539 = n8017 & n13509;
  assign n13540 = n7774 & n8017;
  assign n16580 = (n13398 & n13539) | (n13398 & n13540) | (n13539 & n13540);
  assign n16581 = (n13539 & n13540) | (n13539 & n16459) | (n13540 & n16459);
  assign n16582 = (n13258 & n16580) | (n13258 & n16581) | (n16580 & n16581);
  assign n13542 = n8017 | n13509;
  assign n13543 = n7774 | n8017;
  assign n16583 = (n13398 & n13542) | (n13398 & n13543) | (n13542 & n13543);
  assign n16584 = (n13542 & n13543) | (n13542 & n16459) | (n13543 & n16459);
  assign n16585 = (n13258 & n16583) | (n13258 & n16584) | (n16583 & n16584);
  assign n8020 = ~n16582 & n16585;
  assign n8021 = x73 & x87;
  assign n8022 = n8020 & n8021;
  assign n8023 = n8020 | n8021;
  assign n8024 = ~n8022 & n8023;
  assign n13545 = n7781 & n8024;
  assign n13546 = (n8024 & n13445) | (n8024 & n13545) | (n13445 & n13545);
  assign n13547 = n7781 | n8024;
  assign n13548 = n13445 | n13547;
  assign n8027 = ~n13546 & n13548;
  assign n8028 = x72 & x88;
  assign n8029 = n8027 & n8028;
  assign n8030 = n8027 | n8028;
  assign n8031 = ~n8029 & n8030;
  assign n8032 = n16534 & n8031;
  assign n8033 = n16534 | n8031;
  assign n8034 = ~n8032 & n8033;
  assign n8035 = x71 & x89;
  assign n8036 = n8034 & n8035;
  assign n8037 = n8034 | n8035;
  assign n8038 = ~n8036 & n8037;
  assign n13504 = n7795 | n7797;
  assign n13549 = n8038 & n13504;
  assign n13550 = n7795 & n8038;
  assign n13551 = (n16457 & n13549) | (n16457 & n13550) | (n13549 & n13550);
  assign n13552 = n8038 | n13504;
  assign n13553 = n7795 | n8038;
  assign n13554 = (n16457 & n13552) | (n16457 & n13553) | (n13552 & n13553);
  assign n8041 = ~n13551 & n13554;
  assign n8042 = x70 & x90;
  assign n8043 = n8041 & n8042;
  assign n8044 = n8041 | n8042;
  assign n8045 = ~n8043 & n8044;
  assign n13555 = n7802 & n8045;
  assign n13556 = (n8045 & n16508) | (n8045 & n13555) | (n16508 & n13555);
  assign n13557 = n7802 | n8045;
  assign n13558 = n16508 | n13557;
  assign n8048 = ~n13556 & n13558;
  assign n8049 = x69 & x91;
  assign n8050 = n8048 & n8049;
  assign n8051 = n8048 | n8049;
  assign n8052 = ~n8050 & n8051;
  assign n13502 = n7809 | n7811;
  assign n16586 = n8052 & n13502;
  assign n16528 = n7572 | n7809;
  assign n16529 = (n7809 & n7811) | (n7809 & n16528) | (n7811 & n16528);
  assign n16587 = n8052 & n16529;
  assign n16588 = (n16433 & n16586) | (n16433 & n16587) | (n16586 & n16587);
  assign n16589 = n8052 | n13502;
  assign n16590 = n8052 | n16529;
  assign n16591 = (n16433 & n16589) | (n16433 & n16590) | (n16589 & n16590);
  assign n8055 = ~n16588 & n16591;
  assign n8056 = x68 & x92;
  assign n8057 = n8055 & n8056;
  assign n8058 = n8055 | n8056;
  assign n8059 = ~n8057 & n8058;
  assign n13559 = n7816 & n8059;
  assign n16592 = (n8059 & n13463) | (n8059 & n13559) | (n13463 & n13559);
  assign n16593 = (n7818 & n8059) | (n7818 & n13559) | (n8059 & n13559);
  assign n16594 = (n13359 & n16592) | (n13359 & n16593) | (n16592 & n16593);
  assign n13561 = n7816 | n8059;
  assign n16595 = n13463 | n13561;
  assign n16596 = n7818 | n13561;
  assign n16597 = (n13359 & n16595) | (n13359 & n16596) | (n16595 & n16596);
  assign n8062 = ~n16594 & n16597;
  assign n8063 = x67 & x93;
  assign n8064 = n8062 & n8063;
  assign n8065 = n8062 | n8063;
  assign n8066 = ~n8064 & n8065;
  assign n13563 = n7823 & n8066;
  assign n13564 = (n8066 & n13468) | (n8066 & n13563) | (n13468 & n13563);
  assign n13565 = n7823 | n8066;
  assign n13566 = n13468 | n13565;
  assign n8069 = ~n13564 & n13566;
  assign n8070 = x66 & x94;
  assign n8071 = n8069 & n8070;
  assign n8072 = n8069 | n8070;
  assign n8073 = ~n8071 & n8072;
  assign n13567 = n7830 & n8073;
  assign n13568 = (n8073 & n13473) | (n8073 & n13567) | (n13473 & n13567);
  assign n13569 = n7830 | n8073;
  assign n13570 = n13473 | n13569;
  assign n8076 = ~n13568 & n13570;
  assign n8077 = x65 & x95;
  assign n8078 = n8076 & n8077;
  assign n8079 = n8076 | n8077;
  assign n8080 = ~n8078 & n8079;
  assign n13499 = n7837 | n7839;
  assign n13571 = n8080 & n13499;
  assign n13572 = n7837 & n8080;
  assign n13573 = (n13387 & n13571) | (n13387 & n13572) | (n13571 & n13572);
  assign n13574 = n8080 | n13499;
  assign n13575 = n7837 | n8080;
  assign n13576 = (n13387 & n13574) | (n13387 & n13575) | (n13574 & n13575);
  assign n8083 = ~n13573 & n13576;
  assign n8084 = x64 & x96;
  assign n8085 = n8083 & n8084;
  assign n8086 = n8083 | n8084;
  assign n8087 = ~n8085 & n8086;
  assign n13497 = n7844 | n7846;
  assign n16598 = n8087 & n13497;
  assign n16599 = n7844 & n8087;
  assign n16600 = (n13385 & n16598) | (n13385 & n16599) | (n16598 & n16599);
  assign n16601 = n8087 | n13497;
  assign n16602 = n7844 | n8087;
  assign n16603 = (n13385 & n16601) | (n13385 & n16602) | (n16601 & n16602);
  assign n8090 = ~n16600 & n16603;
  assign n8091 = x63 & x97;
  assign n8092 = n8090 & n8091;
  assign n8093 = n8090 | n8091;
  assign n8094 = ~n8092 & n8093;
  assign n13495 = n7851 | n7853;
  assign n16604 = n8094 & n13495;
  assign n16605 = n7851 & n8094;
  assign n16606 = (n13383 & n16604) | (n13383 & n16605) | (n16604 & n16605);
  assign n16607 = n8094 | n13495;
  assign n16608 = n7851 | n8094;
  assign n16609 = (n13383 & n16607) | (n13383 & n16608) | (n16607 & n16608);
  assign n8097 = ~n16606 & n16609;
  assign n8098 = x62 & x98;
  assign n8099 = n8097 & n8098;
  assign n8100 = n8097 | n8098;
  assign n8101 = ~n8099 & n8100;
  assign n8102 = n13494 & n8101;
  assign n8103 = n13494 | n8101;
  assign n8104 = ~n8102 & n8103;
  assign n8105 = x61 & x99;
  assign n8106 = n8104 & n8105;
  assign n8107 = n8104 | n8105;
  assign n8108 = ~n8106 & n8107;
  assign n8109 = n13492 & n8108;
  assign n8110 = n13492 | n8108;
  assign n8111 = ~n8109 & n8110;
  assign n8112 = x60 & x100;
  assign n8113 = n8111 & n8112;
  assign n8114 = n8111 | n8112;
  assign n8115 = ~n8113 & n8114;
  assign n8116 = n13490 & n8115;
  assign n8117 = n13490 | n8115;
  assign n8118 = ~n8116 & n8117;
  assign n8119 = x59 & x101;
  assign n8120 = n8118 & n8119;
  assign n8121 = n8118 | n8119;
  assign n8122 = ~n8120 & n8121;
  assign n8123 = n13488 & n8122;
  assign n8124 = n13488 | n8122;
  assign n8125 = ~n8123 & n8124;
  assign n8126 = x58 & x102;
  assign n8127 = n8125 & n8126;
  assign n8128 = n8125 | n8126;
  assign n8129 = ~n8127 & n8128;
  assign n8130 = n13486 & n8129;
  assign n8131 = n13486 | n8129;
  assign n8132 = ~n8130 & n8131;
  assign n8133 = x57 & x103;
  assign n8134 = n8132 & n8133;
  assign n8135 = n8132 | n8133;
  assign n8136 = ~n8134 & n8135;
  assign n8137 = n13484 & n8136;
  assign n8138 = n13484 | n8136;
  assign n8139 = ~n8137 & n8138;
  assign n8140 = x56 & x104;
  assign n8141 = n8139 & n8140;
  assign n8142 = n8139 | n8140;
  assign n8143 = ~n8141 & n8142;
  assign n8144 = n7958 & n8143;
  assign n8145 = n7958 | n8143;
  assign n8146 = ~n8144 & n8145;
  assign n8147 = x55 & x105;
  assign n8148 = n8146 & n8147;
  assign n8149 = n8146 | n8147;
  assign n8150 = ~n8148 & n8149;
  assign n8151 = n7957 & n8150;
  assign n8152 = n7957 | n8150;
  assign n8153 = ~n8151 & n8152;
  assign n8154 = x54 & x106;
  assign n8155 = n8153 & n8154;
  assign n8156 = n8153 | n8154;
  assign n8157 = ~n8155 & n8156;
  assign n8158 = n7956 & n8157;
  assign n8159 = n7956 | n8157;
  assign n8160 = ~n8158 & n8159;
  assign n8161 = x53 & x107;
  assign n8162 = n8160 & n8161;
  assign n8163 = n8160 | n8161;
  assign n8164 = ~n8162 & n8163;
  assign n8165 = n16527 & n8164;
  assign n8166 = n16527 | n8164;
  assign n8167 = ~n8165 & n8166;
  assign n8168 = x52 & x108;
  assign n8169 = n8167 & n8168;
  assign n8170 = n8167 | n8168;
  assign n8171 = ~n8169 & n8170;
  assign n8172 = n13482 & n8171;
  assign n8173 = n13482 | n8171;
  assign n8174 = ~n8172 & n8173;
  assign n8175 = x51 & x109;
  assign n8176 = n8174 & n8175;
  assign n8177 = n8174 | n8175;
  assign n8178 = ~n8176 & n8177;
  assign n8179 = n13480 & n8178;
  assign n8180 = n13480 | n8178;
  assign n8181 = ~n8179 & n8180;
  assign n8182 = x50 & x110;
  assign n8183 = n8181 & n8182;
  assign n8184 = n8181 | n8182;
  assign n8185 = ~n8183 & n8184;
  assign n8186 = n13478 & n8185;
  assign n8187 = n13478 | n8185;
  assign n8188 = ~n8186 & n8187;
  assign n8189 = x49 & x111;
  assign n8190 = n8188 & n8189;
  assign n8191 = n8188 | n8189;
  assign n8192 = ~n8190 & n8191;
  assign n8193 = n7949 & n8192;
  assign n8194 = n7949 | n8192;
  assign n8195 = ~n8193 & n8194;
  assign n17774 = n7948 | n8189;
  assign n17775 = (n7947 & n8189) | (n7947 & n17774) | (n8189 & n17774);
  assign n16611 = (n7949 & n8188) | (n7949 & n17775) | (n8188 & n17775);
  assign n13578 = (n8190 & n8192) | (n8190 & n16611) | (n8192 & n16611);
  assign n13579 = n8183 | n13478;
  assign n13580 = (n8183 & n8185) | (n8183 & n13579) | (n8185 & n13579);
  assign n13581 = n8176 | n13480;
  assign n13582 = (n8176 & n8178) | (n8176 & n13581) | (n8178 & n13581);
  assign n13583 = n8169 | n13482;
  assign n13584 = (n8169 & n8171) | (n8169 & n13583) | (n8171 & n13583);
  assign n16612 = n8162 | n16527;
  assign n16613 = (n8162 & n8164) | (n8162 & n16612) | (n8164 & n16612);
  assign n8201 = n8155 | n8158;
  assign n8202 = n8148 | n8151;
  assign n13585 = n8141 | n8143;
  assign n13586 = (n7958 & n8141) | (n7958 & n13585) | (n8141 & n13585);
  assign n13587 = n8134 | n8136;
  assign n13588 = (n8134 & n13484) | (n8134 & n13587) | (n13484 & n13587);
  assign n13589 = n8127 | n8129;
  assign n13590 = (n8127 & n13486) | (n8127 & n13589) | (n13486 & n13589);
  assign n13591 = n8120 | n8122;
  assign n13592 = (n8120 & n13488) | (n8120 & n13591) | (n13488 & n13591);
  assign n13593 = n8113 | n8115;
  assign n13594 = (n8113 & n13490) | (n8113 & n13593) | (n13490 & n13593);
  assign n13595 = n8106 | n8108;
  assign n13596 = (n8106 & n13492) | (n8106 & n13595) | (n13492 & n13595);
  assign n13496 = (n7851 & n13383) | (n7851 & n13495) | (n13383 & n13495);
  assign n13498 = (n7844 & n13385) | (n7844 & n13497) | (n13385 & n13497);
  assign n13503 = (n16433 & n16529) | (n16433 & n13502) | (n16529 & n13502);
  assign n13399 = (n13258 & n16459) | (n13258 & n13398) | (n16459 & n13398);
  assign n13511 = n7767 | n13437;
  assign n8226 = x79 & x82;
  assign n16620 = n7982 & n8226;
  assign n16621 = n16544 & n16620;
  assign n16622 = n16546 & n16620;
  assign n16623 = (n13322 & n16621) | (n13322 & n16622) | (n16621 & n16622);
  assign n16624 = (n16388 & n16621) | (n16388 & n16622) | (n16621 & n16622);
  assign n16625 = (n16123 & n16623) | (n16123 & n16624) | (n16623 & n16624);
  assign n16626 = n7982 | n8226;
  assign n16627 = (n8226 & n16544) | (n8226 & n16626) | (n16544 & n16626);
  assign n16628 = (n8226 & n16546) | (n8226 & n16626) | (n16546 & n16626);
  assign n16629 = (n13322 & n16627) | (n13322 & n16628) | (n16627 & n16628);
  assign n16630 = (n16388 & n16627) | (n16388 & n16628) | (n16627 & n16628);
  assign n16631 = (n16123 & n16629) | (n16123 & n16630) | (n16629 & n16630);
  assign n8229 = ~n16625 & n16631;
  assign n13629 = n7987 & n8229;
  assign n13630 = (n8229 & n16561) | (n8229 & n13629) | (n16561 & n13629);
  assign n13631 = n7987 | n8229;
  assign n13632 = n16561 | n13631;
  assign n8232 = ~n13630 & n13632;
  assign n8233 = x78 & x83;
  assign n8234 = n8232 & n8233;
  assign n8235 = n8232 | n8233;
  assign n8236 = ~n8234 & n8235;
  assign n13621 = n7994 | n7996;
  assign n13633 = n8236 & n13621;
  assign n13634 = n7994 & n8236;
  assign n13635 = (n16542 & n13633) | (n16542 & n13634) | (n13633 & n13634);
  assign n13636 = n8236 | n13621;
  assign n13637 = n7994 | n8236;
  assign n13638 = (n16542 & n13636) | (n16542 & n13637) | (n13636 & n13637);
  assign n8239 = ~n13635 & n13638;
  assign n8240 = x77 & x84;
  assign n8241 = n8239 & n8240;
  assign n8242 = n8239 | n8240;
  assign n8243 = ~n8241 & n8242;
  assign n16632 = n7760 | n8001;
  assign n16633 = (n8001 & n8003) | (n8001 & n16632) | (n8003 & n16632);
  assign n13639 = n8243 & n16633;
  assign n13619 = n8001 | n8003;
  assign n13640 = n8243 & n13619;
  assign n16634 = (n13431 & n13639) | (n13431 & n13640) | (n13639 & n13640);
  assign n16635 = (n13432 & n13639) | (n13432 & n13640) | (n13639 & n13640);
  assign n16636 = (n13228 & n16634) | (n13228 & n16635) | (n16634 & n16635);
  assign n13642 = n8243 | n16633;
  assign n13643 = n8243 | n13619;
  assign n16637 = (n13431 & n13642) | (n13431 & n13643) | (n13642 & n13643);
  assign n16638 = (n13432 & n13642) | (n13432 & n13643) | (n13642 & n13643);
  assign n16639 = (n13228 & n16637) | (n13228 & n16638) | (n16637 & n16638);
  assign n8246 = ~n16636 & n16639;
  assign n8247 = x76 & x85;
  assign n8248 = n8246 & n8247;
  assign n8249 = n8246 | n8247;
  assign n8250 = ~n8248 & n8249;
  assign n13616 = n8008 | n8010;
  assign n13645 = n8250 & n13616;
  assign n13646 = n8008 & n8250;
  assign n16640 = (n13511 & n13645) | (n13511 & n13646) | (n13645 & n13646);
  assign n16641 = (n13645 & n13646) | (n13645 & n16536) | (n13646 & n16536);
  assign n16642 = (n13316 & n16640) | (n13316 & n16641) | (n16640 & n16641);
  assign n13648 = n8250 | n13616;
  assign n13649 = n8008 | n8250;
  assign n16643 = (n13511 & n13648) | (n13511 & n13649) | (n13648 & n13649);
  assign n16644 = (n13648 & n13649) | (n13648 & n16536) | (n13649 & n16536);
  assign n16645 = (n13316 & n16643) | (n13316 & n16644) | (n16643 & n16644);
  assign n8253 = ~n16642 & n16645;
  assign n8254 = x75 & x86;
  assign n8255 = n8253 & n8254;
  assign n8256 = n8253 | n8254;
  assign n8257 = ~n8255 & n8256;
  assign n17776 = n8015 & n8257;
  assign n17777 = (n8257 & n13539) | (n8257 & n17776) | (n13539 & n17776);
  assign n16618 = n7774 | n8015;
  assign n16619 = (n8015 & n8017) | (n8015 & n16618) | (n8017 & n16618);
  assign n16647 = n8257 & n16619;
  assign n16648 = (n13399 & n17777) | (n13399 & n16647) | (n17777 & n16647);
  assign n17778 = n8015 | n8257;
  assign n17779 = n13539 | n17778;
  assign n16650 = n8257 | n16619;
  assign n16651 = (n13399 & n17779) | (n13399 & n16650) | (n17779 & n16650);
  assign n8260 = ~n16648 & n16651;
  assign n8261 = x74 & x87;
  assign n8262 = n8260 & n8261;
  assign n8263 = n8260 | n8261;
  assign n8264 = ~n8262 & n8263;
  assign n13611 = n8022 | n8024;
  assign n16652 = n8264 & n13611;
  assign n16616 = n7781 | n8022;
  assign n16617 = (n8022 & n8024) | (n8022 & n16616) | (n8024 & n16616);
  assign n16653 = n8264 & n16617;
  assign n16654 = (n13445 & n16652) | (n13445 & n16653) | (n16652 & n16653);
  assign n16655 = n8264 | n13611;
  assign n16656 = n8264 | n16617;
  assign n16657 = (n13445 & n16655) | (n13445 & n16656) | (n16655 & n16656);
  assign n8267 = ~n16654 & n16657;
  assign n8268 = x73 & x88;
  assign n8269 = n8267 & n8268;
  assign n8270 = n8267 | n8268;
  assign n8271 = ~n8269 & n8270;
  assign n13608 = n8029 | n8031;
  assign n13651 = n8271 & n13608;
  assign n13652 = n8029 & n8271;
  assign n13653 = (n16534 & n13651) | (n16534 & n13652) | (n13651 & n13652);
  assign n13654 = n8271 | n13608;
  assign n13655 = n8029 | n8271;
  assign n13656 = (n16534 & n13654) | (n16534 & n13655) | (n13654 & n13655);
  assign n8274 = ~n13653 & n13656;
  assign n8275 = x72 & x89;
  assign n8276 = n8274 & n8275;
  assign n8277 = n8274 | n8275;
  assign n8278 = ~n8276 & n8277;
  assign n13657 = n8036 & n8278;
  assign n16658 = (n8278 & n13550) | (n8278 & n13657) | (n13550 & n13657);
  assign n16659 = (n8278 & n13549) | (n8278 & n13657) | (n13549 & n13657);
  assign n16660 = (n16457 & n16658) | (n16457 & n16659) | (n16658 & n16659);
  assign n13659 = n8036 | n8278;
  assign n16661 = n13550 | n13659;
  assign n16662 = n13549 | n13659;
  assign n16663 = (n16457 & n16661) | (n16457 & n16662) | (n16661 & n16662);
  assign n8281 = ~n16660 & n16663;
  assign n8282 = x71 & x90;
  assign n8283 = n8281 & n8282;
  assign n8284 = n8281 | n8282;
  assign n8285 = ~n8283 & n8284;
  assign n13606 = n8043 | n8045;
  assign n16664 = n8285 & n13606;
  assign n16614 = n7802 | n8043;
  assign n16615 = (n8043 & n8045) | (n8043 & n16614) | (n8045 & n16614);
  assign n16665 = n8285 & n16615;
  assign n16666 = (n16508 & n16664) | (n16508 & n16665) | (n16664 & n16665);
  assign n16667 = n8285 | n13606;
  assign n16668 = n8285 | n16615;
  assign n16669 = (n16508 & n16667) | (n16508 & n16668) | (n16667 & n16668);
  assign n8288 = ~n16666 & n16669;
  assign n8289 = x70 & x91;
  assign n8290 = n8288 & n8289;
  assign n8291 = n8288 | n8289;
  assign n8292 = ~n8290 & n8291;
  assign n13603 = n8050 | n8052;
  assign n13661 = n8292 & n13603;
  assign n13662 = n8050 & n8292;
  assign n13663 = (n13503 & n13661) | (n13503 & n13662) | (n13661 & n13662);
  assign n13664 = n8292 | n13603;
  assign n13665 = n8050 | n8292;
  assign n13666 = (n13503 & n13664) | (n13503 & n13665) | (n13664 & n13665);
  assign n8295 = ~n13663 & n13666;
  assign n8296 = x69 & x92;
  assign n8297 = n8295 & n8296;
  assign n8298 = n8295 | n8296;
  assign n8299 = ~n8297 & n8298;
  assign n13667 = n8057 & n8299;
  assign n13668 = (n8299 & n16594) | (n8299 & n13667) | (n16594 & n13667);
  assign n13669 = n8057 | n8299;
  assign n13670 = n16594 | n13669;
  assign n8302 = ~n13668 & n13670;
  assign n8303 = x68 & x93;
  assign n8304 = n8302 & n8303;
  assign n8305 = n8302 | n8303;
  assign n8306 = ~n8304 & n8305;
  assign n13671 = n8064 & n8306;
  assign n13672 = (n8306 & n13564) | (n8306 & n13671) | (n13564 & n13671);
  assign n13673 = n8064 | n8306;
  assign n13674 = n13564 | n13673;
  assign n8309 = ~n13672 & n13674;
  assign n8310 = x67 & x94;
  assign n8311 = n8309 & n8310;
  assign n8312 = n8309 | n8310;
  assign n8313 = ~n8311 & n8312;
  assign n13675 = n8071 & n8313;
  assign n13676 = (n8313 & n13568) | (n8313 & n13675) | (n13568 & n13675);
  assign n13677 = n8071 | n8313;
  assign n13678 = n13568 | n13677;
  assign n8316 = ~n13676 & n13678;
  assign n8317 = x66 & x95;
  assign n8318 = n8316 & n8317;
  assign n8319 = n8316 | n8317;
  assign n8320 = ~n8318 & n8319;
  assign n13679 = n8078 & n8320;
  assign n13680 = (n8320 & n13573) | (n8320 & n13679) | (n13573 & n13679);
  assign n13681 = n8078 | n8320;
  assign n13682 = n13573 | n13681;
  assign n8323 = ~n13680 & n13682;
  assign n8324 = x65 & x96;
  assign n8325 = n8323 & n8324;
  assign n8326 = n8323 | n8324;
  assign n8327 = ~n8325 & n8326;
  assign n13601 = n8085 | n8087;
  assign n13683 = n8327 & n13601;
  assign n13684 = n8085 & n8327;
  assign n13685 = (n13498 & n13683) | (n13498 & n13684) | (n13683 & n13684);
  assign n13686 = n8327 | n13601;
  assign n13687 = n8085 | n8327;
  assign n13688 = (n13498 & n13686) | (n13498 & n13687) | (n13686 & n13687);
  assign n8330 = ~n13685 & n13688;
  assign n8331 = x64 & x97;
  assign n8332 = n8330 & n8331;
  assign n8333 = n8330 | n8331;
  assign n8334 = ~n8332 & n8333;
  assign n13599 = n8092 | n8094;
  assign n16670 = n8334 & n13599;
  assign n16671 = n8092 & n8334;
  assign n16672 = (n13496 & n16670) | (n13496 & n16671) | (n16670 & n16671);
  assign n16673 = n8334 | n13599;
  assign n16674 = n8092 | n8334;
  assign n16675 = (n13496 & n16673) | (n13496 & n16674) | (n16673 & n16674);
  assign n8337 = ~n16672 & n16675;
  assign n8338 = x63 & x98;
  assign n8339 = n8337 & n8338;
  assign n8340 = n8337 | n8338;
  assign n8341 = ~n8339 & n8340;
  assign n13597 = n8099 | n8101;
  assign n16676 = n8341 & n13597;
  assign n16677 = n8099 & n8341;
  assign n16678 = (n13494 & n16676) | (n13494 & n16677) | (n16676 & n16677);
  assign n16679 = n8341 | n13597;
  assign n16680 = n8099 | n8341;
  assign n16681 = (n13494 & n16679) | (n13494 & n16680) | (n16679 & n16680);
  assign n8344 = ~n16678 & n16681;
  assign n8345 = x62 & x99;
  assign n8346 = n8344 & n8345;
  assign n8347 = n8344 | n8345;
  assign n8348 = ~n8346 & n8347;
  assign n8349 = n13596 & n8348;
  assign n8350 = n13596 | n8348;
  assign n8351 = ~n8349 & n8350;
  assign n8352 = x61 & x100;
  assign n8353 = n8351 & n8352;
  assign n8354 = n8351 | n8352;
  assign n8355 = ~n8353 & n8354;
  assign n8356 = n13594 & n8355;
  assign n8357 = n13594 | n8355;
  assign n8358 = ~n8356 & n8357;
  assign n8359 = x60 & x101;
  assign n8360 = n8358 & n8359;
  assign n8361 = n8358 | n8359;
  assign n8362 = ~n8360 & n8361;
  assign n8363 = n13592 & n8362;
  assign n8364 = n13592 | n8362;
  assign n8365 = ~n8363 & n8364;
  assign n8366 = x59 & x102;
  assign n8367 = n8365 & n8366;
  assign n8368 = n8365 | n8366;
  assign n8369 = ~n8367 & n8368;
  assign n8370 = n13590 & n8369;
  assign n8371 = n13590 | n8369;
  assign n8372 = ~n8370 & n8371;
  assign n8373 = x58 & x103;
  assign n8374 = n8372 & n8373;
  assign n8375 = n8372 | n8373;
  assign n8376 = ~n8374 & n8375;
  assign n8377 = n13588 & n8376;
  assign n8378 = n13588 | n8376;
  assign n8379 = ~n8377 & n8378;
  assign n8380 = x57 & x104;
  assign n8381 = n8379 & n8380;
  assign n8382 = n8379 | n8380;
  assign n8383 = ~n8381 & n8382;
  assign n8384 = n13586 & n8383;
  assign n8385 = n13586 | n8383;
  assign n8386 = ~n8384 & n8385;
  assign n8387 = x56 & x105;
  assign n8388 = n8386 & n8387;
  assign n8389 = n8386 | n8387;
  assign n8390 = ~n8388 & n8389;
  assign n8391 = n8202 & n8390;
  assign n8392 = n8202 | n8390;
  assign n8393 = ~n8391 & n8392;
  assign n8394 = x55 & x106;
  assign n8395 = n8393 & n8394;
  assign n8396 = n8393 | n8394;
  assign n8397 = ~n8395 & n8396;
  assign n8398 = n8201 & n8397;
  assign n8399 = n8201 | n8397;
  assign n8400 = ~n8398 & n8399;
  assign n8401 = x54 & x107;
  assign n8402 = n8400 & n8401;
  assign n8403 = n8400 | n8401;
  assign n8404 = ~n8402 & n8403;
  assign n8405 = n16613 & n8404;
  assign n8406 = n16613 | n8404;
  assign n8407 = ~n8405 & n8406;
  assign n8408 = x53 & x108;
  assign n8409 = n8407 & n8408;
  assign n8410 = n8407 | n8408;
  assign n8411 = ~n8409 & n8410;
  assign n8412 = n13584 & n8411;
  assign n8413 = n13584 | n8411;
  assign n8414 = ~n8412 & n8413;
  assign n8415 = x52 & x109;
  assign n8416 = n8414 & n8415;
  assign n8417 = n8414 | n8415;
  assign n8418 = ~n8416 & n8417;
  assign n8419 = n13582 & n8418;
  assign n8420 = n13582 | n8418;
  assign n8421 = ~n8419 & n8420;
  assign n8422 = x51 & x110;
  assign n8423 = n8421 & n8422;
  assign n8424 = n8421 | n8422;
  assign n8425 = ~n8423 & n8424;
  assign n8426 = n13580 & n8425;
  assign n8427 = n13580 | n8425;
  assign n8428 = ~n8426 & n8427;
  assign n8429 = x50 & x111;
  assign n8430 = n8428 & n8429;
  assign n8431 = n8428 | n8429;
  assign n8432 = ~n8430 & n8431;
  assign n8433 = n13578 & n8432;
  assign n8434 = n13578 | n8432;
  assign n8435 = ~n8433 & n8434;
  assign n13689 = n8430 | n13578;
  assign n13690 = (n8430 & n8432) | (n8430 & n13689) | (n8432 & n13689);
  assign n13691 = n8423 | n13580;
  assign n13692 = (n8423 & n8425) | (n8423 & n13691) | (n8425 & n13691);
  assign n13693 = n8416 | n13582;
  assign n13694 = (n8416 & n8418) | (n8416 & n13693) | (n8418 & n13693);
  assign n13695 = n8409 | n13584;
  assign n13696 = (n8409 & n8411) | (n8409 & n13695) | (n8411 & n13695);
  assign n16682 = n8402 | n16613;
  assign n16683 = (n8402 & n8404) | (n8402 & n16682) | (n8404 & n16682);
  assign n8441 = n8395 | n8398;
  assign n13697 = n8388 | n8390;
  assign n13698 = (n8202 & n8388) | (n8202 & n13697) | (n8388 & n13697);
  assign n13699 = n8381 | n8383;
  assign n13700 = (n8381 & n13586) | (n8381 & n13699) | (n13586 & n13699);
  assign n13701 = n8374 | n8376;
  assign n13702 = (n8374 & n13588) | (n8374 & n13701) | (n13588 & n13701);
  assign n13703 = n8367 | n8369;
  assign n13704 = (n8367 & n13590) | (n8367 & n13703) | (n13590 & n13703);
  assign n13705 = n8360 | n8362;
  assign n13706 = (n8360 & n13592) | (n8360 & n13705) | (n13592 & n13705);
  assign n13707 = n8353 | n8355;
  assign n13708 = (n8353 & n13594) | (n8353 & n13707) | (n13594 & n13707);
  assign n13598 = (n8099 & n13494) | (n8099 & n13597) | (n13494 & n13597);
  assign n13600 = (n8092 & n13496) | (n8092 & n13599) | (n13496 & n13599);
  assign n13721 = n8276 | n8278;
  assign n16686 = n8036 | n8276;
  assign n16687 = (n8276 & n8278) | (n8276 & n16686) | (n8278 & n16686);
  assign n16688 = (n13550 & n13721) | (n13550 & n16687) | (n13721 & n16687);
  assign n16689 = (n13549 & n13721) | (n13549 & n16687) | (n13721 & n16687);
  assign n16690 = (n16457 & n16688) | (n16457 & n16689) | (n16688 & n16689);
  assign n13612 = (n13445 & n16617) | (n13445 & n13611) | (n16617 & n13611);
  assign n13614 = n8015 | n13539;
  assign n16691 = n8248 | n8250;
  assign n16692 = (n8248 & n13616) | (n8248 & n16691) | (n13616 & n16691);
  assign n16693 = n8008 | n8248;
  assign n16694 = (n8248 & n8250) | (n8248 & n16693) | (n8250 & n16693);
  assign n16695 = (n13511 & n16692) | (n13511 & n16694) | (n16692 & n16694);
  assign n16696 = (n16536 & n16692) | (n16536 & n16694) | (n16692 & n16694);
  assign n16697 = (n13316 & n16695) | (n13316 & n16696) | (n16695 & n16696);
  assign n8466 = x79 & x83;
  assign n16698 = n8229 | n16625;
  assign n16699 = (n7987 & n16625) | (n7987 & n16698) | (n16625 & n16698);
  assign n13736 = n8466 & n16699;
  assign n17780 = n8466 & n16624;
  assign n17781 = n8466 & n16623;
  assign n17782 = (n16123 & n17780) | (n16123 & n17781) | (n17780 & n17781);
  assign n16701 = (n8229 & n8466) | (n8229 & n17782) | (n8466 & n17782);
  assign n13738 = (n16561 & n13736) | (n16561 & n16701) | (n13736 & n16701);
  assign n13739 = n8466 | n16699;
  assign n17783 = n8466 | n16624;
  assign n17784 = n8466 | n16623;
  assign n17785 = (n16123 & n17783) | (n16123 & n17784) | (n17783 & n17784);
  assign n16703 = n8229 | n17785;
  assign n13741 = (n16561 & n13739) | (n16561 & n16703) | (n13739 & n16703);
  assign n8469 = ~n13738 & n13741;
  assign n16704 = n8234 & n8469;
  assign n16705 = (n8469 & n13633) | (n8469 & n16704) | (n13633 & n16704);
  assign n16706 = n7994 | n8234;
  assign n16707 = (n8234 & n8236) | (n8234 & n16706) | (n8236 & n16706);
  assign n13743 = n8469 & n16707;
  assign n13744 = (n16542 & n16705) | (n16542 & n13743) | (n16705 & n13743);
  assign n16708 = n8234 | n8469;
  assign n16709 = n13633 | n16708;
  assign n13746 = n8469 | n16707;
  assign n13747 = (n16542 & n16709) | (n16542 & n13746) | (n16709 & n13746);
  assign n8472 = ~n13744 & n13747;
  assign n8473 = x78 & x84;
  assign n8474 = n8472 & n8473;
  assign n8475 = n8472 | n8473;
  assign n8476 = ~n8474 & n8475;
  assign n13748 = n8241 & n8476;
  assign n13749 = (n8476 & n16636) | (n8476 & n13748) | (n16636 & n13748);
  assign n13750 = n8241 | n8476;
  assign n13751 = n16636 | n13750;
  assign n8479 = ~n13749 & n13751;
  assign n8480 = x77 & x85;
  assign n8481 = n8479 & n8480;
  assign n8482 = n8479 | n8480;
  assign n8483 = ~n8481 & n8482;
  assign n8484 = n16697 & n8483;
  assign n8485 = n16697 | n8483;
  assign n8486 = ~n8484 & n8485;
  assign n8487 = x76 & x86;
  assign n8488 = n8486 & n8487;
  assign n8489 = n8486 | n8487;
  assign n8490 = ~n8488 & n8489;
  assign n13725 = n8255 | n8257;
  assign n13752 = n8490 & n13725;
  assign n13753 = n8255 & n8490;
  assign n16710 = (n13614 & n13752) | (n13614 & n13753) | (n13752 & n13753);
  assign n16711 = (n13752 & n13753) | (n13752 & n16619) | (n13753 & n16619);
  assign n16712 = (n13399 & n16710) | (n13399 & n16711) | (n16710 & n16711);
  assign n13755 = n8490 | n13725;
  assign n13756 = n8255 | n8490;
  assign n16713 = (n13614 & n13755) | (n13614 & n13756) | (n13755 & n13756);
  assign n16714 = (n13755 & n13756) | (n13755 & n16619) | (n13756 & n16619);
  assign n16715 = (n13399 & n16713) | (n13399 & n16714) | (n16713 & n16714);
  assign n8493 = ~n16712 & n16715;
  assign n8494 = x75 & x87;
  assign n8495 = n8493 & n8494;
  assign n8496 = n8493 | n8494;
  assign n8497 = ~n8495 & n8496;
  assign n13723 = n8262 | n8264;
  assign n13758 = n8497 & n13723;
  assign n13759 = n8262 & n8497;
  assign n13760 = (n13612 & n13758) | (n13612 & n13759) | (n13758 & n13759);
  assign n13761 = n8497 | n13723;
  assign n13762 = n8262 | n8497;
  assign n13763 = (n13612 & n13761) | (n13612 & n13762) | (n13761 & n13762);
  assign n8500 = ~n13760 & n13763;
  assign n8501 = x74 & x88;
  assign n8502 = n8500 & n8501;
  assign n8503 = n8500 | n8501;
  assign n8504 = ~n8502 & n8503;
  assign n13764 = n8269 & n8504;
  assign n13765 = (n8504 & n13653) | (n8504 & n13764) | (n13653 & n13764);
  assign n13766 = n8269 | n8504;
  assign n13767 = n13653 | n13766;
  assign n8507 = ~n13765 & n13767;
  assign n8508 = x73 & x89;
  assign n8509 = n8507 & n8508;
  assign n8510 = n8507 | n8508;
  assign n8511 = ~n8509 & n8510;
  assign n8512 = n16690 & n8511;
  assign n8513 = n16690 | n8511;
  assign n8514 = ~n8512 & n8513;
  assign n8515 = x72 & x90;
  assign n8516 = n8514 & n8515;
  assign n8517 = n8514 | n8515;
  assign n8518 = ~n8516 & n8517;
  assign n13718 = n8283 | n8285;
  assign n13768 = n8518 & n13718;
  assign n13769 = n8283 & n8518;
  assign n16716 = (n13606 & n13768) | (n13606 & n13769) | (n13768 & n13769);
  assign n16717 = (n13768 & n13769) | (n13768 & n16615) | (n13769 & n16615);
  assign n16718 = (n16508 & n16716) | (n16508 & n16717) | (n16716 & n16717);
  assign n13771 = n8518 | n13718;
  assign n13772 = n8283 | n8518;
  assign n16719 = (n13606 & n13771) | (n13606 & n13772) | (n13771 & n13772);
  assign n16720 = (n13771 & n13772) | (n13771 & n16615) | (n13772 & n16615);
  assign n16721 = (n16508 & n16719) | (n16508 & n16720) | (n16719 & n16720);
  assign n8521 = ~n16718 & n16721;
  assign n8522 = x71 & x91;
  assign n8523 = n8521 & n8522;
  assign n8524 = n8521 | n8522;
  assign n8525 = ~n8523 & n8524;
  assign n13774 = n8290 & n8525;
  assign n16722 = (n8525 & n13661) | (n8525 & n13774) | (n13661 & n13774);
  assign n16723 = (n8525 & n13662) | (n8525 & n13774) | (n13662 & n13774);
  assign n16724 = (n13503 & n16722) | (n13503 & n16723) | (n16722 & n16723);
  assign n13776 = n8290 | n8525;
  assign n16725 = n13661 | n13776;
  assign n16726 = n13662 | n13776;
  assign n16727 = (n13503 & n16725) | (n13503 & n16726) | (n16725 & n16726);
  assign n8528 = ~n16724 & n16727;
  assign n8529 = x70 & x92;
  assign n8530 = n8528 & n8529;
  assign n8531 = n8528 | n8529;
  assign n8532 = ~n8530 & n8531;
  assign n13716 = n8297 | n8299;
  assign n16728 = n8532 & n13716;
  assign n16684 = n8057 | n8297;
  assign n16685 = (n8297 & n8299) | (n8297 & n16684) | (n8299 & n16684);
  assign n16729 = n8532 & n16685;
  assign n16730 = (n16594 & n16728) | (n16594 & n16729) | (n16728 & n16729);
  assign n16731 = n8532 | n13716;
  assign n16732 = n8532 | n16685;
  assign n16733 = (n16594 & n16731) | (n16594 & n16732) | (n16731 & n16732);
  assign n8535 = ~n16730 & n16733;
  assign n8536 = x69 & x93;
  assign n8537 = n8535 & n8536;
  assign n8538 = n8535 | n8536;
  assign n8539 = ~n8537 & n8538;
  assign n13778 = n8304 & n8539;
  assign n16734 = (n8539 & n13671) | (n8539 & n13778) | (n13671 & n13778);
  assign n16735 = (n8306 & n8539) | (n8306 & n13778) | (n8539 & n13778);
  assign n16736 = (n13564 & n16734) | (n13564 & n16735) | (n16734 & n16735);
  assign n13780 = n8304 | n8539;
  assign n16737 = n13671 | n13780;
  assign n16738 = n8306 | n13780;
  assign n16739 = (n13564 & n16737) | (n13564 & n16738) | (n16737 & n16738);
  assign n8542 = ~n16736 & n16739;
  assign n8543 = x68 & x94;
  assign n8544 = n8542 & n8543;
  assign n8545 = n8542 | n8543;
  assign n8546 = ~n8544 & n8545;
  assign n13782 = n8311 & n8546;
  assign n13783 = (n8546 & n13676) | (n8546 & n13782) | (n13676 & n13782);
  assign n13784 = n8311 | n8546;
  assign n13785 = n13676 | n13784;
  assign n8549 = ~n13783 & n13785;
  assign n8550 = x67 & x95;
  assign n8551 = n8549 & n8550;
  assign n8552 = n8549 | n8550;
  assign n8553 = ~n8551 & n8552;
  assign n13786 = n8318 & n8553;
  assign n13787 = (n8553 & n13680) | (n8553 & n13786) | (n13680 & n13786);
  assign n13788 = n8318 | n8553;
  assign n13789 = n13680 | n13788;
  assign n8556 = ~n13787 & n13789;
  assign n8557 = x66 & x96;
  assign n8558 = n8556 & n8557;
  assign n8559 = n8556 | n8557;
  assign n8560 = ~n8558 & n8559;
  assign n13790 = n8325 & n8560;
  assign n13791 = (n8560 & n13685) | (n8560 & n13790) | (n13685 & n13790);
  assign n13792 = n8325 | n8560;
  assign n13793 = n13685 | n13792;
  assign n8563 = ~n13791 & n13793;
  assign n8564 = x65 & x97;
  assign n8565 = n8563 & n8564;
  assign n8566 = n8563 | n8564;
  assign n8567 = ~n8565 & n8566;
  assign n13713 = n8332 | n8334;
  assign n13794 = n8567 & n13713;
  assign n13795 = n8332 & n8567;
  assign n13796 = (n13600 & n13794) | (n13600 & n13795) | (n13794 & n13795);
  assign n13797 = n8567 | n13713;
  assign n13798 = n8332 | n8567;
  assign n13799 = (n13600 & n13797) | (n13600 & n13798) | (n13797 & n13798);
  assign n8570 = ~n13796 & n13799;
  assign n8571 = x64 & x98;
  assign n8572 = n8570 & n8571;
  assign n8573 = n8570 | n8571;
  assign n8574 = ~n8572 & n8573;
  assign n13711 = n8339 | n8341;
  assign n16740 = n8574 & n13711;
  assign n16741 = n8339 & n8574;
  assign n16742 = (n13598 & n16740) | (n13598 & n16741) | (n16740 & n16741);
  assign n16743 = n8574 | n13711;
  assign n16744 = n8339 | n8574;
  assign n16745 = (n13598 & n16743) | (n13598 & n16744) | (n16743 & n16744);
  assign n8577 = ~n16742 & n16745;
  assign n8578 = x63 & x99;
  assign n8579 = n8577 & n8578;
  assign n8580 = n8577 | n8578;
  assign n8581 = ~n8579 & n8580;
  assign n13709 = n8346 | n8348;
  assign n16746 = n8581 & n13709;
  assign n16747 = n8346 & n8581;
  assign n16748 = (n13596 & n16746) | (n13596 & n16747) | (n16746 & n16747);
  assign n16749 = n8581 | n13709;
  assign n16750 = n8346 | n8581;
  assign n16751 = (n13596 & n16749) | (n13596 & n16750) | (n16749 & n16750);
  assign n8584 = ~n16748 & n16751;
  assign n8585 = x62 & x100;
  assign n8586 = n8584 & n8585;
  assign n8587 = n8584 | n8585;
  assign n8588 = ~n8586 & n8587;
  assign n8589 = n13708 & n8588;
  assign n8590 = n13708 | n8588;
  assign n8591 = ~n8589 & n8590;
  assign n8592 = x61 & x101;
  assign n8593 = n8591 & n8592;
  assign n8594 = n8591 | n8592;
  assign n8595 = ~n8593 & n8594;
  assign n8596 = n13706 & n8595;
  assign n8597 = n13706 | n8595;
  assign n8598 = ~n8596 & n8597;
  assign n8599 = x60 & x102;
  assign n8600 = n8598 & n8599;
  assign n8601 = n8598 | n8599;
  assign n8602 = ~n8600 & n8601;
  assign n8603 = n13704 & n8602;
  assign n8604 = n13704 | n8602;
  assign n8605 = ~n8603 & n8604;
  assign n8606 = x59 & x103;
  assign n8607 = n8605 & n8606;
  assign n8608 = n8605 | n8606;
  assign n8609 = ~n8607 & n8608;
  assign n8610 = n13702 & n8609;
  assign n8611 = n13702 | n8609;
  assign n8612 = ~n8610 & n8611;
  assign n8613 = x58 & x104;
  assign n8614 = n8612 & n8613;
  assign n8615 = n8612 | n8613;
  assign n8616 = ~n8614 & n8615;
  assign n8617 = n13700 & n8616;
  assign n8618 = n13700 | n8616;
  assign n8619 = ~n8617 & n8618;
  assign n8620 = x57 & x105;
  assign n8621 = n8619 & n8620;
  assign n8622 = n8619 | n8620;
  assign n8623 = ~n8621 & n8622;
  assign n8624 = n13698 & n8623;
  assign n8625 = n13698 | n8623;
  assign n8626 = ~n8624 & n8625;
  assign n8627 = x56 & x106;
  assign n8628 = n8626 & n8627;
  assign n8629 = n8626 | n8627;
  assign n8630 = ~n8628 & n8629;
  assign n8631 = n8441 & n8630;
  assign n8632 = n8441 | n8630;
  assign n8633 = ~n8631 & n8632;
  assign n8634 = x55 & x107;
  assign n8635 = n8633 & n8634;
  assign n8636 = n8633 | n8634;
  assign n8637 = ~n8635 & n8636;
  assign n8638 = n16683 & n8637;
  assign n8639 = n16683 | n8637;
  assign n8640 = ~n8638 & n8639;
  assign n8641 = x54 & x108;
  assign n8642 = n8640 & n8641;
  assign n8643 = n8640 | n8641;
  assign n8644 = ~n8642 & n8643;
  assign n8645 = n13696 & n8644;
  assign n8646 = n13696 | n8644;
  assign n8647 = ~n8645 & n8646;
  assign n8648 = x53 & x109;
  assign n8649 = n8647 & n8648;
  assign n8650 = n8647 | n8648;
  assign n8651 = ~n8649 & n8650;
  assign n8652 = n13694 & n8651;
  assign n8653 = n13694 | n8651;
  assign n8654 = ~n8652 & n8653;
  assign n8655 = x52 & x110;
  assign n8656 = n8654 & n8655;
  assign n8657 = n8654 | n8655;
  assign n8658 = ~n8656 & n8657;
  assign n8659 = n13692 & n8658;
  assign n8660 = n13692 | n8658;
  assign n8661 = ~n8659 & n8660;
  assign n8662 = x51 & x111;
  assign n8663 = n8661 & n8662;
  assign n8664 = n8661 | n8662;
  assign n8665 = ~n8663 & n8664;
  assign n8666 = n13690 & n8665;
  assign n8667 = n13690 | n8665;
  assign n8668 = ~n8666 & n8667;
  assign n13800 = n8663 | n13690;
  assign n13801 = (n8663 & n8665) | (n8663 & n13800) | (n8665 & n13800);
  assign n13802 = n8656 | n13692;
  assign n13803 = (n8656 & n8658) | (n8656 & n13802) | (n8658 & n13802);
  assign n13804 = n8649 | n13694;
  assign n13805 = (n8649 & n8651) | (n8649 & n13804) | (n8651 & n13804);
  assign n13806 = n8642 | n13696;
  assign n13807 = (n8642 & n8644) | (n8642 & n13806) | (n8644 & n13806);
  assign n16752 = n8635 | n16683;
  assign n16753 = (n8635 & n8637) | (n8635 & n16752) | (n8637 & n16752);
  assign n13808 = n8628 | n8630;
  assign n13809 = (n8441 & n8628) | (n8441 & n13808) | (n8628 & n13808);
  assign n13810 = n8621 | n8623;
  assign n13811 = (n8621 & n13698) | (n8621 & n13810) | (n13698 & n13810);
  assign n13812 = n8614 | n8616;
  assign n13813 = (n8614 & n13700) | (n8614 & n13812) | (n13700 & n13812);
  assign n13814 = n8607 | n8609;
  assign n13815 = (n8607 & n13702) | (n8607 & n13814) | (n13702 & n13814);
  assign n13816 = n8600 | n8602;
  assign n13817 = (n8600 & n13704) | (n8600 & n13816) | (n13704 & n13816);
  assign n13818 = n8593 | n8595;
  assign n13819 = (n8593 & n13706) | (n8593 & n13818) | (n13706 & n13818);
  assign n13710 = (n8346 & n13596) | (n8346 & n13709) | (n13596 & n13709);
  assign n13712 = (n8339 & n13598) | (n8339 & n13711) | (n13598 & n13711);
  assign n13717 = (n16594 & n16685) | (n16594 & n13716) | (n16685 & n13716);
  assign n13829 = n8523 | n8525;
  assign n16754 = n8290 | n8523;
  assign n16755 = (n8523 & n8525) | (n8523 & n16754) | (n8525 & n16754);
  assign n16756 = (n13661 & n13829) | (n13661 & n16755) | (n13829 & n16755);
  assign n16757 = (n13662 & n13829) | (n13662 & n16755) | (n13829 & n16755);
  assign n16758 = (n13503 & n16756) | (n13503 & n16757) | (n16756 & n16757);
  assign n13615 = (n13399 & n16619) | (n13399 & n13614) | (n16619 & n13614);
  assign n8698 = x79 & x84;
  assign n16763 = n8469 | n13738;
  assign n17786 = (n8234 & n13738) | (n8234 & n16763) | (n13738 & n16763);
  assign n17787 = n8698 & n17786;
  assign n17788 = n8698 & n16763;
  assign n17789 = (n13633 & n17787) | (n13633 & n17788) | (n17787 & n17788);
  assign n17790 = n8698 & n13738;
  assign n17791 = (n16707 & n17788) | (n16707 & n17790) | (n17788 & n17790);
  assign n16769 = (n16542 & n17789) | (n16542 & n17791) | (n17789 & n17791);
  assign n17792 = n8698 | n17786;
  assign n17793 = n8698 | n16763;
  assign n17794 = (n13633 & n17792) | (n13633 & n17793) | (n17792 & n17793);
  assign n17795 = n8698 | n13738;
  assign n17796 = (n16707 & n17793) | (n16707 & n17795) | (n17793 & n17795);
  assign n16772 = (n16542 & n17794) | (n16542 & n17796) | (n17794 & n17796);
  assign n8701 = ~n16769 & n16772;
  assign n16773 = n8241 | n8474;
  assign n16774 = (n8474 & n8476) | (n8474 & n16773) | (n8476 & n16773);
  assign n13847 = n8701 & n16774;
  assign n16775 = n8474 & n8701;
  assign n16776 = (n8476 & n8701) | (n8476 & n16775) | (n8701 & n16775);
  assign n13849 = (n16636 & n13847) | (n16636 & n16776) | (n13847 & n16776);
  assign n13850 = n8701 | n16774;
  assign n16777 = n8474 | n8701;
  assign n16778 = n8476 | n16777;
  assign n13852 = (n16636 & n13850) | (n16636 & n16778) | (n13850 & n16778);
  assign n8704 = ~n13849 & n13852;
  assign n8705 = x78 & x85;
  assign n8706 = n8704 & n8705;
  assign n8707 = n8704 | n8705;
  assign n8708 = ~n8706 & n8707;
  assign n13839 = n8481 | n8483;
  assign n13853 = n8708 & n13839;
  assign n13854 = n8481 & n8708;
  assign n13855 = (n16697 & n13853) | (n16697 & n13854) | (n13853 & n13854);
  assign n13856 = n8708 | n13839;
  assign n13857 = n8481 | n8708;
  assign n13858 = (n16697 & n13856) | (n16697 & n13857) | (n13856 & n13857);
  assign n8711 = ~n13855 & n13858;
  assign n8712 = x77 & x86;
  assign n8713 = n8711 & n8712;
  assign n8714 = n8711 | n8712;
  assign n8715 = ~n8713 & n8714;
  assign n17797 = n8488 & n8715;
  assign n17798 = (n8715 & n13752) | (n8715 & n17797) | (n13752 & n17797);
  assign n16761 = n8255 | n8488;
  assign n16762 = (n8488 & n8490) | (n8488 & n16761) | (n8490 & n16761);
  assign n16780 = n8715 & n16762;
  assign n16781 = (n13615 & n17798) | (n13615 & n16780) | (n17798 & n16780);
  assign n17799 = n8488 | n8715;
  assign n17800 = n13752 | n17799;
  assign n16783 = n8715 | n16762;
  assign n16784 = (n13615 & n17800) | (n13615 & n16783) | (n17800 & n16783);
  assign n8718 = ~n16781 & n16784;
  assign n8719 = x76 & x87;
  assign n8720 = n8718 & n8719;
  assign n8721 = n8718 | n8719;
  assign n8722 = ~n8720 & n8721;
  assign n13859 = n8495 & n8722;
  assign n16785 = (n8722 & n13758) | (n8722 & n13859) | (n13758 & n13859);
  assign n16786 = (n8722 & n13759) | (n8722 & n13859) | (n13759 & n13859);
  assign n16787 = (n13612 & n16785) | (n13612 & n16786) | (n16785 & n16786);
  assign n13861 = n8495 | n8722;
  assign n16788 = n13758 | n13861;
  assign n16789 = n13759 | n13861;
  assign n16790 = (n13612 & n16788) | (n13612 & n16789) | (n16788 & n16789);
  assign n8725 = ~n16787 & n16790;
  assign n8726 = x75 & x88;
  assign n8727 = n8725 & n8726;
  assign n8728 = n8725 | n8726;
  assign n8729 = ~n8727 & n8728;
  assign n13834 = n8502 | n8504;
  assign n16791 = n8729 & n13834;
  assign n16759 = n8269 | n8502;
  assign n16760 = (n8502 & n8504) | (n8502 & n16759) | (n8504 & n16759);
  assign n16792 = n8729 & n16760;
  assign n16793 = (n13653 & n16791) | (n13653 & n16792) | (n16791 & n16792);
  assign n16794 = n8729 | n13834;
  assign n16795 = n8729 | n16760;
  assign n16796 = (n13653 & n16794) | (n13653 & n16795) | (n16794 & n16795);
  assign n8732 = ~n16793 & n16796;
  assign n8733 = x74 & x89;
  assign n8734 = n8732 & n8733;
  assign n8735 = n8732 | n8733;
  assign n8736 = ~n8734 & n8735;
  assign n13831 = n8509 | n8511;
  assign n13863 = n8736 & n13831;
  assign n13864 = n8509 & n8736;
  assign n13865 = (n16690 & n13863) | (n16690 & n13864) | (n13863 & n13864);
  assign n13866 = n8736 | n13831;
  assign n13867 = n8509 | n8736;
  assign n13868 = (n16690 & n13866) | (n16690 & n13867) | (n13866 & n13867);
  assign n8739 = ~n13865 & n13868;
  assign n8740 = x73 & x90;
  assign n8741 = n8739 & n8740;
  assign n8742 = n8739 | n8740;
  assign n8743 = ~n8741 & n8742;
  assign n13869 = n8516 & n8743;
  assign n13870 = (n8743 & n16718) | (n8743 & n13869) | (n16718 & n13869);
  assign n13871 = n8516 | n8743;
  assign n13872 = n16718 | n13871;
  assign n8746 = ~n13870 & n13872;
  assign n8747 = x72 & x91;
  assign n8748 = n8746 & n8747;
  assign n8749 = n8746 | n8747;
  assign n8750 = ~n8748 & n8749;
  assign n8751 = n16758 & n8750;
  assign n8752 = n16758 | n8750;
  assign n8753 = ~n8751 & n8752;
  assign n8754 = x71 & x92;
  assign n8755 = n8753 & n8754;
  assign n8756 = n8753 | n8754;
  assign n8757 = ~n8755 & n8756;
  assign n13826 = n8530 | n8532;
  assign n13873 = n8757 & n13826;
  assign n13874 = n8530 & n8757;
  assign n13875 = (n13717 & n13873) | (n13717 & n13874) | (n13873 & n13874);
  assign n13876 = n8757 | n13826;
  assign n13877 = n8530 | n8757;
  assign n13878 = (n13717 & n13876) | (n13717 & n13877) | (n13876 & n13877);
  assign n8760 = ~n13875 & n13878;
  assign n8761 = x70 & x93;
  assign n8762 = n8760 & n8761;
  assign n8763 = n8760 | n8761;
  assign n8764 = ~n8762 & n8763;
  assign n13879 = n8537 & n8764;
  assign n13880 = (n8764 & n16736) | (n8764 & n13879) | (n16736 & n13879);
  assign n13881 = n8537 | n8764;
  assign n13882 = n16736 | n13881;
  assign n8767 = ~n13880 & n13882;
  assign n8768 = x69 & x94;
  assign n8769 = n8767 & n8768;
  assign n8770 = n8767 | n8768;
  assign n8771 = ~n8769 & n8770;
  assign n13883 = n8544 & n8771;
  assign n13884 = (n8771 & n13783) | (n8771 & n13883) | (n13783 & n13883);
  assign n13885 = n8544 | n8771;
  assign n13886 = n13783 | n13885;
  assign n8774 = ~n13884 & n13886;
  assign n8775 = x68 & x95;
  assign n8776 = n8774 & n8775;
  assign n8777 = n8774 | n8775;
  assign n8778 = ~n8776 & n8777;
  assign n13887 = n8551 & n8778;
  assign n13888 = (n8778 & n13787) | (n8778 & n13887) | (n13787 & n13887);
  assign n13889 = n8551 | n8778;
  assign n13890 = n13787 | n13889;
  assign n8781 = ~n13888 & n13890;
  assign n8782 = x67 & x96;
  assign n8783 = n8781 & n8782;
  assign n8784 = n8781 | n8782;
  assign n8785 = ~n8783 & n8784;
  assign n13891 = n8558 & n8785;
  assign n13892 = (n8785 & n13791) | (n8785 & n13891) | (n13791 & n13891);
  assign n13893 = n8558 | n8785;
  assign n13894 = n13791 | n13893;
  assign n8788 = ~n13892 & n13894;
  assign n8789 = x66 & x97;
  assign n8790 = n8788 & n8789;
  assign n8791 = n8788 | n8789;
  assign n8792 = ~n8790 & n8791;
  assign n13895 = n8565 & n8792;
  assign n13896 = (n8792 & n13796) | (n8792 & n13895) | (n13796 & n13895);
  assign n13897 = n8565 | n8792;
  assign n13898 = n13796 | n13897;
  assign n8795 = ~n13896 & n13898;
  assign n8796 = x65 & x98;
  assign n8797 = n8795 & n8796;
  assign n8798 = n8795 | n8796;
  assign n8799 = ~n8797 & n8798;
  assign n13824 = n8572 | n8574;
  assign n13899 = n8799 & n13824;
  assign n13900 = n8572 & n8799;
  assign n13901 = (n13712 & n13899) | (n13712 & n13900) | (n13899 & n13900);
  assign n13902 = n8799 | n13824;
  assign n13903 = n8572 | n8799;
  assign n13904 = (n13712 & n13902) | (n13712 & n13903) | (n13902 & n13903);
  assign n8802 = ~n13901 & n13904;
  assign n8803 = x64 & x99;
  assign n8804 = n8802 & n8803;
  assign n8805 = n8802 | n8803;
  assign n8806 = ~n8804 & n8805;
  assign n13822 = n8579 | n8581;
  assign n16797 = n8806 & n13822;
  assign n16798 = n8579 & n8806;
  assign n16799 = (n13710 & n16797) | (n13710 & n16798) | (n16797 & n16798);
  assign n16800 = n8806 | n13822;
  assign n16801 = n8579 | n8806;
  assign n16802 = (n13710 & n16800) | (n13710 & n16801) | (n16800 & n16801);
  assign n8809 = ~n16799 & n16802;
  assign n8810 = x63 & x100;
  assign n8811 = n8809 & n8810;
  assign n8812 = n8809 | n8810;
  assign n8813 = ~n8811 & n8812;
  assign n13820 = n8586 | n8588;
  assign n16803 = n8813 & n13820;
  assign n16804 = n8586 & n8813;
  assign n16805 = (n13708 & n16803) | (n13708 & n16804) | (n16803 & n16804);
  assign n16806 = n8813 | n13820;
  assign n16807 = n8586 | n8813;
  assign n16808 = (n13708 & n16806) | (n13708 & n16807) | (n16806 & n16807);
  assign n8816 = ~n16805 & n16808;
  assign n8817 = x62 & x101;
  assign n8818 = n8816 & n8817;
  assign n8819 = n8816 | n8817;
  assign n8820 = ~n8818 & n8819;
  assign n8821 = n13819 & n8820;
  assign n8822 = n13819 | n8820;
  assign n8823 = ~n8821 & n8822;
  assign n8824 = x61 & x102;
  assign n8825 = n8823 & n8824;
  assign n8826 = n8823 | n8824;
  assign n8827 = ~n8825 & n8826;
  assign n8828 = n13817 & n8827;
  assign n8829 = n13817 | n8827;
  assign n8830 = ~n8828 & n8829;
  assign n8831 = x60 & x103;
  assign n8832 = n8830 & n8831;
  assign n8833 = n8830 | n8831;
  assign n8834 = ~n8832 & n8833;
  assign n8835 = n13815 & n8834;
  assign n8836 = n13815 | n8834;
  assign n8837 = ~n8835 & n8836;
  assign n8838 = x59 & x104;
  assign n8839 = n8837 & n8838;
  assign n8840 = n8837 | n8838;
  assign n8841 = ~n8839 & n8840;
  assign n8842 = n13813 & n8841;
  assign n8843 = n13813 | n8841;
  assign n8844 = ~n8842 & n8843;
  assign n8845 = x58 & x105;
  assign n8846 = n8844 & n8845;
  assign n8847 = n8844 | n8845;
  assign n8848 = ~n8846 & n8847;
  assign n8849 = n13811 & n8848;
  assign n8850 = n13811 | n8848;
  assign n8851 = ~n8849 & n8850;
  assign n8852 = x57 & x106;
  assign n8853 = n8851 & n8852;
  assign n8854 = n8851 | n8852;
  assign n8855 = ~n8853 & n8854;
  assign n8856 = n13809 & n8855;
  assign n8857 = n13809 | n8855;
  assign n8858 = ~n8856 & n8857;
  assign n8859 = x56 & x107;
  assign n8860 = n8858 & n8859;
  assign n8861 = n8858 | n8859;
  assign n8862 = ~n8860 & n8861;
  assign n8863 = n16753 & n8862;
  assign n8864 = n16753 | n8862;
  assign n8865 = ~n8863 & n8864;
  assign n8866 = x55 & x108;
  assign n8867 = n8865 & n8866;
  assign n8868 = n8865 | n8866;
  assign n8869 = ~n8867 & n8868;
  assign n8870 = n13807 & n8869;
  assign n8871 = n13807 | n8869;
  assign n8872 = ~n8870 & n8871;
  assign n8873 = x54 & x109;
  assign n8874 = n8872 & n8873;
  assign n8875 = n8872 | n8873;
  assign n8876 = ~n8874 & n8875;
  assign n8877 = n13805 & n8876;
  assign n8878 = n13805 | n8876;
  assign n8879 = ~n8877 & n8878;
  assign n8880 = x53 & x110;
  assign n8881 = n8879 & n8880;
  assign n8882 = n8879 | n8880;
  assign n8883 = ~n8881 & n8882;
  assign n8884 = n13803 & n8883;
  assign n8885 = n13803 | n8883;
  assign n8886 = ~n8884 & n8885;
  assign n8887 = x52 & x111;
  assign n8888 = n8886 & n8887;
  assign n8889 = n8886 | n8887;
  assign n8890 = ~n8888 & n8889;
  assign n8891 = n13801 & n8890;
  assign n8892 = n13801 | n8890;
  assign n8893 = ~n8891 & n8892;
  assign n13905 = n8888 | n13801;
  assign n13906 = (n8888 & n8890) | (n8888 & n13905) | (n8890 & n13905);
  assign n13907 = n8881 | n13803;
  assign n13908 = (n8881 & n8883) | (n8881 & n13907) | (n8883 & n13907);
  assign n13909 = n8874 | n13805;
  assign n13910 = (n8874 & n8876) | (n8874 & n13909) | (n8876 & n13909);
  assign n13911 = n8867 | n13807;
  assign n13912 = (n8867 & n8869) | (n8867 & n13911) | (n8869 & n13911);
  assign n13913 = n8860 | n8862;
  assign n13914 = (n16753 & n8860) | (n16753 & n13913) | (n8860 & n13913);
  assign n13915 = n8853 | n8855;
  assign n13916 = (n8853 & n13809) | (n8853 & n13915) | (n13809 & n13915);
  assign n13917 = n8846 | n8848;
  assign n13918 = (n8846 & n13811) | (n8846 & n13917) | (n13811 & n13917);
  assign n13919 = n8839 | n8841;
  assign n13920 = (n8839 & n13813) | (n8839 & n13919) | (n13813 & n13919);
  assign n13921 = n8832 | n8834;
  assign n13922 = (n8832 & n13815) | (n8832 & n13921) | (n13815 & n13921);
  assign n13923 = n8825 | n8827;
  assign n13924 = (n8825 & n13817) | (n8825 & n13923) | (n13817 & n13923);
  assign n13821 = (n8586 & n13708) | (n8586 & n13820) | (n13708 & n13820);
  assign n13823 = (n8579 & n13710) | (n8579 & n13822) | (n13710 & n13822);
  assign n13835 = (n13653 & n16760) | (n13653 & n13834) | (n16760 & n13834);
  assign n13942 = n8720 | n8722;
  assign n16813 = n8495 | n8720;
  assign n16814 = (n8720 & n8722) | (n8720 & n16813) | (n8722 & n16813);
  assign n16815 = (n13758 & n13942) | (n13758 & n16814) | (n13942 & n16814);
  assign n16816 = (n13759 & n13942) | (n13759 & n16814) | (n13942 & n16814);
  assign n16817 = (n13612 & n16815) | (n13612 & n16816) | (n16815 & n16816);
  assign n13837 = n8488 | n13752;
  assign n8922 = x79 & x85;
  assign n17801 = n8922 & n16769;
  assign n17802 = (n8922 & n16776) | (n8922 & n17801) | (n16776 & n17801);
  assign n16822 = n8701 | n16769;
  assign n17803 = n8922 & n16822;
  assign n17804 = (n16774 & n17801) | (n16774 & n17803) | (n17801 & n17803);
  assign n16826 = (n16636 & n17802) | (n16636 & n17804) | (n17802 & n17804);
  assign n17805 = n8922 | n16769;
  assign n17806 = n16776 | n17805;
  assign n17807 = n8922 | n16822;
  assign n17808 = (n16774 & n17805) | (n16774 & n17807) | (n17805 & n17807);
  assign n16829 = (n16636 & n17806) | (n16636 & n17808) | (n17806 & n17808);
  assign n8925 = ~n16826 & n16829;
  assign n16818 = n8706 | n8708;
  assign n16819 = (n8706 & n13839) | (n8706 & n16818) | (n13839 & n16818);
  assign n16830 = n8925 & n16819;
  assign n16820 = n8481 | n8706;
  assign n16821 = (n8706 & n8708) | (n8706 & n16820) | (n8708 & n16820);
  assign n16831 = n8925 & n16821;
  assign n16832 = (n16697 & n16830) | (n16697 & n16831) | (n16830 & n16831);
  assign n16833 = n8925 | n16819;
  assign n16834 = n8925 | n16821;
  assign n16835 = (n16697 & n16833) | (n16697 & n16834) | (n16833 & n16834);
  assign n8928 = ~n16832 & n16835;
  assign n8929 = x78 & x86;
  assign n8930 = n8928 & n8929;
  assign n8931 = n8928 | n8929;
  assign n8932 = ~n8930 & n8931;
  assign n13944 = n8713 | n8715;
  assign n13952 = n8932 & n13944;
  assign n13953 = n8713 & n8932;
  assign n16836 = (n13837 & n13952) | (n13837 & n13953) | (n13952 & n13953);
  assign n16837 = (n13952 & n13953) | (n13952 & n16762) | (n13953 & n16762);
  assign n16838 = (n13615 & n16836) | (n13615 & n16837) | (n16836 & n16837);
  assign n13955 = n8932 | n13944;
  assign n13956 = n8713 | n8932;
  assign n16839 = (n13837 & n13955) | (n13837 & n13956) | (n13955 & n13956);
  assign n16840 = (n13955 & n13956) | (n13955 & n16762) | (n13956 & n16762);
  assign n16841 = (n13615 & n16839) | (n13615 & n16840) | (n16839 & n16840);
  assign n8935 = ~n16838 & n16841;
  assign n8936 = x77 & x87;
  assign n8937 = n8935 & n8936;
  assign n8938 = n8935 | n8936;
  assign n8939 = ~n8937 & n8938;
  assign n8940 = n16817 & n8939;
  assign n8941 = n16817 | n8939;
  assign n8942 = ~n8940 & n8941;
  assign n8943 = x76 & x88;
  assign n8944 = n8942 & n8943;
  assign n8945 = n8942 | n8943;
  assign n8946 = ~n8944 & n8945;
  assign n13939 = n8727 | n8729;
  assign n13958 = n8946 & n13939;
  assign n13959 = n8727 & n8946;
  assign n13960 = (n13835 & n13958) | (n13835 & n13959) | (n13958 & n13959);
  assign n13961 = n8946 | n13939;
  assign n13962 = n8727 | n8946;
  assign n13963 = (n13835 & n13961) | (n13835 & n13962) | (n13961 & n13962);
  assign n8949 = ~n13960 & n13963;
  assign n8950 = x75 & x89;
  assign n8951 = n8949 & n8950;
  assign n8952 = n8949 | n8950;
  assign n8953 = ~n8951 & n8952;
  assign n13964 = n8734 & n8953;
  assign n13965 = (n8953 & n13865) | (n8953 & n13964) | (n13865 & n13964);
  assign n13966 = n8734 | n8953;
  assign n13967 = n13865 | n13966;
  assign n8956 = ~n13965 & n13967;
  assign n8957 = x74 & x90;
  assign n8958 = n8956 & n8957;
  assign n8959 = n8956 | n8957;
  assign n8960 = ~n8958 & n8959;
  assign n13937 = n8741 | n8743;
  assign n16842 = n8960 & n13937;
  assign n16811 = n8516 | n8741;
  assign n16812 = (n8741 & n8743) | (n8741 & n16811) | (n8743 & n16811);
  assign n16843 = n8960 & n16812;
  assign n16844 = (n16718 & n16842) | (n16718 & n16843) | (n16842 & n16843);
  assign n16845 = n8960 | n13937;
  assign n16846 = n8960 | n16812;
  assign n16847 = (n16718 & n16845) | (n16718 & n16846) | (n16845 & n16846);
  assign n8963 = ~n16844 & n16847;
  assign n8964 = x73 & x91;
  assign n8965 = n8963 & n8964;
  assign n8966 = n8963 | n8964;
  assign n8967 = ~n8965 & n8966;
  assign n13934 = n8748 | n8750;
  assign n13968 = n8967 & n13934;
  assign n13969 = n8748 & n8967;
  assign n13970 = (n16758 & n13968) | (n16758 & n13969) | (n13968 & n13969);
  assign n13971 = n8967 | n13934;
  assign n13972 = n8748 | n8967;
  assign n13973 = (n16758 & n13971) | (n16758 & n13972) | (n13971 & n13972);
  assign n8970 = ~n13970 & n13973;
  assign n8971 = x72 & x92;
  assign n8972 = n8970 & n8971;
  assign n8973 = n8970 | n8971;
  assign n8974 = ~n8972 & n8973;
  assign n13974 = n8755 & n8974;
  assign n16848 = (n8974 & n13874) | (n8974 & n13974) | (n13874 & n13974);
  assign n16849 = (n8974 & n13873) | (n8974 & n13974) | (n13873 & n13974);
  assign n16850 = (n13717 & n16848) | (n13717 & n16849) | (n16848 & n16849);
  assign n13976 = n8755 | n8974;
  assign n16851 = n13874 | n13976;
  assign n16852 = n13873 | n13976;
  assign n16853 = (n13717 & n16851) | (n13717 & n16852) | (n16851 & n16852);
  assign n8977 = ~n16850 & n16853;
  assign n8978 = x71 & x93;
  assign n8979 = n8977 & n8978;
  assign n8980 = n8977 | n8978;
  assign n8981 = ~n8979 & n8980;
  assign n13932 = n8762 | n8764;
  assign n16854 = n8981 & n13932;
  assign n16809 = n8537 | n8762;
  assign n16810 = (n8762 & n8764) | (n8762 & n16809) | (n8764 & n16809);
  assign n16855 = n8981 & n16810;
  assign n16856 = (n16736 & n16854) | (n16736 & n16855) | (n16854 & n16855);
  assign n16857 = n8981 | n13932;
  assign n16858 = n8981 | n16810;
  assign n16859 = (n16736 & n16857) | (n16736 & n16858) | (n16857 & n16858);
  assign n8984 = ~n16856 & n16859;
  assign n8985 = x70 & x94;
  assign n8986 = n8984 & n8985;
  assign n8987 = n8984 | n8985;
  assign n8988 = ~n8986 & n8987;
  assign n13978 = n8769 & n8988;
  assign n16860 = (n8988 & n13883) | (n8988 & n13978) | (n13883 & n13978);
  assign n16861 = (n8771 & n8988) | (n8771 & n13978) | (n8988 & n13978);
  assign n16862 = (n13783 & n16860) | (n13783 & n16861) | (n16860 & n16861);
  assign n13980 = n8769 | n8988;
  assign n16863 = n13883 | n13980;
  assign n16864 = n8771 | n13980;
  assign n16865 = (n13783 & n16863) | (n13783 & n16864) | (n16863 & n16864);
  assign n8991 = ~n16862 & n16865;
  assign n8992 = x69 & x95;
  assign n8993 = n8991 & n8992;
  assign n8994 = n8991 | n8992;
  assign n8995 = ~n8993 & n8994;
  assign n13982 = n8776 & n8995;
  assign n13983 = (n8995 & n13888) | (n8995 & n13982) | (n13888 & n13982);
  assign n13984 = n8776 | n8995;
  assign n13985 = n13888 | n13984;
  assign n8998 = ~n13983 & n13985;
  assign n8999 = x68 & x96;
  assign n9000 = n8998 & n8999;
  assign n9001 = n8998 | n8999;
  assign n9002 = ~n9000 & n9001;
  assign n13986 = n8783 & n9002;
  assign n13987 = (n9002 & n13892) | (n9002 & n13986) | (n13892 & n13986);
  assign n13988 = n8783 | n9002;
  assign n13989 = n13892 | n13988;
  assign n9005 = ~n13987 & n13989;
  assign n9006 = x67 & x97;
  assign n9007 = n9005 & n9006;
  assign n9008 = n9005 | n9006;
  assign n9009 = ~n9007 & n9008;
  assign n13990 = n8790 & n9009;
  assign n13991 = (n9009 & n13896) | (n9009 & n13990) | (n13896 & n13990);
  assign n13992 = n8790 | n9009;
  assign n13993 = n13896 | n13992;
  assign n9012 = ~n13991 & n13993;
  assign n9013 = x66 & x98;
  assign n9014 = n9012 & n9013;
  assign n9015 = n9012 | n9013;
  assign n9016 = ~n9014 & n9015;
  assign n13994 = n8797 & n9016;
  assign n13995 = (n9016 & n13901) | (n9016 & n13994) | (n13901 & n13994);
  assign n13996 = n8797 | n9016;
  assign n13997 = n13901 | n13996;
  assign n9019 = ~n13995 & n13997;
  assign n9020 = x65 & x99;
  assign n9021 = n9019 & n9020;
  assign n9022 = n9019 | n9020;
  assign n9023 = ~n9021 & n9022;
  assign n13929 = n8804 | n8806;
  assign n13998 = n9023 & n13929;
  assign n13999 = n8804 & n9023;
  assign n14000 = (n13823 & n13998) | (n13823 & n13999) | (n13998 & n13999);
  assign n14001 = n9023 | n13929;
  assign n14002 = n8804 | n9023;
  assign n14003 = (n13823 & n14001) | (n13823 & n14002) | (n14001 & n14002);
  assign n9026 = ~n14000 & n14003;
  assign n9027 = x64 & x100;
  assign n9028 = n9026 & n9027;
  assign n9029 = n9026 | n9027;
  assign n9030 = ~n9028 & n9029;
  assign n13927 = n8811 | n8813;
  assign n16866 = n9030 & n13927;
  assign n16867 = n8811 & n9030;
  assign n16868 = (n13821 & n16866) | (n13821 & n16867) | (n16866 & n16867);
  assign n16869 = n9030 | n13927;
  assign n16870 = n8811 | n9030;
  assign n16871 = (n13821 & n16869) | (n13821 & n16870) | (n16869 & n16870);
  assign n9033 = ~n16868 & n16871;
  assign n9034 = x63 & x101;
  assign n9035 = n9033 & n9034;
  assign n9036 = n9033 | n9034;
  assign n9037 = ~n9035 & n9036;
  assign n13925 = n8818 | n8820;
  assign n16872 = n9037 & n13925;
  assign n16873 = n8818 & n9037;
  assign n16874 = (n13819 & n16872) | (n13819 & n16873) | (n16872 & n16873);
  assign n16875 = n9037 | n13925;
  assign n16876 = n8818 | n9037;
  assign n16877 = (n13819 & n16875) | (n13819 & n16876) | (n16875 & n16876);
  assign n9040 = ~n16874 & n16877;
  assign n9041 = x62 & x102;
  assign n9042 = n9040 & n9041;
  assign n9043 = n9040 | n9041;
  assign n9044 = ~n9042 & n9043;
  assign n9045 = n13924 & n9044;
  assign n9046 = n13924 | n9044;
  assign n9047 = ~n9045 & n9046;
  assign n9048 = x61 & x103;
  assign n9049 = n9047 & n9048;
  assign n9050 = n9047 | n9048;
  assign n9051 = ~n9049 & n9050;
  assign n9052 = n13922 & n9051;
  assign n9053 = n13922 | n9051;
  assign n9054 = ~n9052 & n9053;
  assign n9055 = x60 & x104;
  assign n9056 = n9054 & n9055;
  assign n9057 = n9054 | n9055;
  assign n9058 = ~n9056 & n9057;
  assign n9059 = n13920 & n9058;
  assign n9060 = n13920 | n9058;
  assign n9061 = ~n9059 & n9060;
  assign n9062 = x59 & x105;
  assign n9063 = n9061 & n9062;
  assign n9064 = n9061 | n9062;
  assign n9065 = ~n9063 & n9064;
  assign n9066 = n13918 & n9065;
  assign n9067 = n13918 | n9065;
  assign n9068 = ~n9066 & n9067;
  assign n9069 = x58 & x106;
  assign n9070 = n9068 & n9069;
  assign n9071 = n9068 | n9069;
  assign n9072 = ~n9070 & n9071;
  assign n9073 = n13916 & n9072;
  assign n9074 = n13916 | n9072;
  assign n9075 = ~n9073 & n9074;
  assign n9076 = x57 & x107;
  assign n9077 = n9075 & n9076;
  assign n9078 = n9075 | n9076;
  assign n9079 = ~n9077 & n9078;
  assign n9080 = n13914 & n9079;
  assign n9081 = n13914 | n9079;
  assign n9082 = ~n9080 & n9081;
  assign n9083 = x56 & x108;
  assign n9084 = n9082 & n9083;
  assign n9085 = n9082 | n9083;
  assign n9086 = ~n9084 & n9085;
  assign n9087 = n13912 & n9086;
  assign n9088 = n13912 | n9086;
  assign n9089 = ~n9087 & n9088;
  assign n9090 = x55 & x109;
  assign n9091 = n9089 & n9090;
  assign n9092 = n9089 | n9090;
  assign n9093 = ~n9091 & n9092;
  assign n9094 = n13910 & n9093;
  assign n9095 = n13910 | n9093;
  assign n9096 = ~n9094 & n9095;
  assign n9097 = x54 & x110;
  assign n9098 = n9096 & n9097;
  assign n9099 = n9096 | n9097;
  assign n9100 = ~n9098 & n9099;
  assign n9101 = n13908 & n9100;
  assign n9102 = n13908 | n9100;
  assign n9103 = ~n9101 & n9102;
  assign n9104 = x53 & x111;
  assign n9105 = n9103 & n9104;
  assign n9106 = n9103 | n9104;
  assign n9107 = ~n9105 & n9106;
  assign n9108 = n13906 & n9107;
  assign n9109 = n13906 | n9107;
  assign n9110 = ~n9108 & n9109;
  assign n9111 = n9105 | n9108;
  assign n9112 = n9098 | n9101;
  assign n9113 = n9091 | n9094;
  assign n9114 = n9084 | n9087;
  assign n14004 = n9077 | n9079;
  assign n14005 = (n9077 & n13914) | (n9077 & n14004) | (n13914 & n14004);
  assign n14006 = n9070 | n9072;
  assign n14007 = (n9070 & n13916) | (n9070 & n14006) | (n13916 & n14006);
  assign n14008 = n9063 | n9065;
  assign n14009 = (n9063 & n13918) | (n9063 & n14008) | (n13918 & n14008);
  assign n14010 = n9056 | n9058;
  assign n14011 = (n9056 & n13920) | (n9056 & n14010) | (n13920 & n14010);
  assign n14012 = n9049 | n9051;
  assign n14013 = (n9049 & n13922) | (n9049 & n14012) | (n13922 & n14012);
  assign n13926 = (n8818 & n13819) | (n8818 & n13925) | (n13819 & n13925);
  assign n13928 = (n8811 & n13821) | (n8811 & n13927) | (n13821 & n13927);
  assign n13933 = (n16736 & n16810) | (n16736 & n13932) | (n16810 & n13932);
  assign n14023 = n8972 | n8974;
  assign n16878 = n8755 | n8972;
  assign n16879 = (n8972 & n8974) | (n8972 & n16878) | (n8974 & n16878);
  assign n16880 = (n13874 & n14023) | (n13874 & n16879) | (n14023 & n16879);
  assign n16881 = (n13873 & n14023) | (n13873 & n16879) | (n14023 & n16879);
  assign n16882 = (n13717 & n16880) | (n13717 & n16881) | (n16880 & n16881);
  assign n13938 = (n16718 & n16812) | (n16718 & n13937) | (n16812 & n13937);
  assign n16885 = n8713 | n8930;
  assign n16886 = (n8930 & n8932) | (n8930 & n16885) | (n8932 & n16885);
  assign n16887 = n8930 | n8932;
  assign n16888 = (n8930 & n13944) | (n8930 & n16887) | (n13944 & n16887);
  assign n16889 = (n13837 & n16886) | (n13837 & n16888) | (n16886 & n16888);
  assign n16890 = (n16762 & n16886) | (n16762 & n16888) | (n16886 & n16888);
  assign n16891 = (n13615 & n16889) | (n13615 & n16890) | (n16889 & n16890);
  assign n9138 = x79 & x86;
  assign n17809 = n9138 & n17804;
  assign n17810 = n9138 & n17802;
  assign n17811 = (n16636 & n17809) | (n16636 & n17810) | (n17809 & n17810);
  assign n16893 = (n8925 & n9138) | (n8925 & n17811) | (n9138 & n17811);
  assign n17812 = n9138 & n17803;
  assign n17813 = n9138 & n17801;
  assign n17814 = (n16774 & n17812) | (n16774 & n17813) | (n17812 & n17813);
  assign n17815 = n8922 & n9138;
  assign n17816 = (n16776 & n17813) | (n16776 & n17815) | (n17813 & n17815);
  assign n16896 = (n16636 & n17814) | (n16636 & n17816) | (n17814 & n17816);
  assign n16897 = (n16819 & n16893) | (n16819 & n16896) | (n16893 & n16896);
  assign n16898 = (n16821 & n16893) | (n16821 & n16896) | (n16893 & n16896);
  assign n16899 = (n16697 & n16897) | (n16697 & n16898) | (n16897 & n16898);
  assign n17817 = n9138 | n17804;
  assign n17818 = n9138 | n17802;
  assign n17819 = (n16636 & n17817) | (n16636 & n17818) | (n17817 & n17818);
  assign n16901 = n8925 | n17819;
  assign n17820 = n9138 | n17803;
  assign n17821 = n9138 | n17801;
  assign n17822 = (n16774 & n17820) | (n16774 & n17821) | (n17820 & n17821);
  assign n17823 = n8922 | n9138;
  assign n17824 = (n16776 & n17821) | (n16776 & n17823) | (n17821 & n17823);
  assign n16904 = (n16636 & n17822) | (n16636 & n17824) | (n17822 & n17824);
  assign n16905 = (n16819 & n16901) | (n16819 & n16904) | (n16901 & n16904);
  assign n16906 = (n16821 & n16901) | (n16821 & n16904) | (n16901 & n16904);
  assign n16907 = (n16697 & n16905) | (n16697 & n16906) | (n16905 & n16906);
  assign n9141 = ~n16899 & n16907;
  assign n9142 = n16891 & n9141;
  assign n9143 = n16891 | n9141;
  assign n9144 = ~n9142 & n9143;
  assign n9145 = x78 & x87;
  assign n9146 = n9144 & n9145;
  assign n9147 = n9144 | n9145;
  assign n9148 = ~n9146 & n9147;
  assign n14030 = n8937 | n8939;
  assign n14043 = n9148 & n14030;
  assign n14044 = n8937 & n9148;
  assign n14045 = (n16817 & n14043) | (n16817 & n14044) | (n14043 & n14044);
  assign n14046 = n9148 | n14030;
  assign n14047 = n8937 | n9148;
  assign n14048 = (n16817 & n14046) | (n16817 & n14047) | (n14046 & n14047);
  assign n9151 = ~n14045 & n14048;
  assign n9152 = x77 & x88;
  assign n9153 = n9151 & n9152;
  assign n9154 = n9151 | n9152;
  assign n9155 = ~n9153 & n9154;
  assign n14049 = n8944 & n9155;
  assign n16908 = (n9155 & n13959) | (n9155 & n14049) | (n13959 & n14049);
  assign n16909 = (n9155 & n13958) | (n9155 & n14049) | (n13958 & n14049);
  assign n16910 = (n13835 & n16908) | (n13835 & n16909) | (n16908 & n16909);
  assign n14051 = n8944 | n9155;
  assign n16911 = n13959 | n14051;
  assign n16912 = n13958 | n14051;
  assign n16913 = (n13835 & n16911) | (n13835 & n16912) | (n16911 & n16912);
  assign n9158 = ~n16910 & n16913;
  assign n9159 = x76 & x89;
  assign n9160 = n9158 & n9159;
  assign n9161 = n9158 | n9159;
  assign n9162 = ~n9160 & n9161;
  assign n14028 = n8951 | n8953;
  assign n16914 = n9162 & n14028;
  assign n16883 = n8734 | n8951;
  assign n16884 = (n8951 & n8953) | (n8951 & n16883) | (n8953 & n16883);
  assign n16915 = n9162 & n16884;
  assign n16916 = (n13865 & n16914) | (n13865 & n16915) | (n16914 & n16915);
  assign n16917 = n9162 | n14028;
  assign n16918 = n9162 | n16884;
  assign n16919 = (n13865 & n16917) | (n13865 & n16918) | (n16917 & n16918);
  assign n9165 = ~n16916 & n16919;
  assign n9166 = x75 & x90;
  assign n9167 = n9165 & n9166;
  assign n9168 = n9165 | n9166;
  assign n9169 = ~n9167 & n9168;
  assign n14025 = n8958 | n8960;
  assign n14053 = n9169 & n14025;
  assign n14054 = n8958 & n9169;
  assign n14055 = (n13938 & n14053) | (n13938 & n14054) | (n14053 & n14054);
  assign n14056 = n9169 | n14025;
  assign n14057 = n8958 | n9169;
  assign n14058 = (n13938 & n14056) | (n13938 & n14057) | (n14056 & n14057);
  assign n9172 = ~n14055 & n14058;
  assign n9173 = x74 & x91;
  assign n9174 = n9172 & n9173;
  assign n9175 = n9172 | n9173;
  assign n9176 = ~n9174 & n9175;
  assign n14059 = n8965 & n9176;
  assign n16920 = (n9176 & n13968) | (n9176 & n14059) | (n13968 & n14059);
  assign n16921 = (n9176 & n13969) | (n9176 & n14059) | (n13969 & n14059);
  assign n16922 = (n16758 & n16920) | (n16758 & n16921) | (n16920 & n16921);
  assign n14061 = n8965 | n9176;
  assign n16923 = n13968 | n14061;
  assign n16924 = n13969 | n14061;
  assign n16925 = (n16758 & n16923) | (n16758 & n16924) | (n16923 & n16924);
  assign n9179 = ~n16922 & n16925;
  assign n9180 = x73 & x92;
  assign n9181 = n9179 & n9180;
  assign n9182 = n9179 | n9180;
  assign n9183 = ~n9181 & n9182;
  assign n9184 = n16882 & n9183;
  assign n9185 = n16882 | n9183;
  assign n9186 = ~n9184 & n9185;
  assign n9187 = x72 & x93;
  assign n9188 = n9186 & n9187;
  assign n9189 = n9186 | n9187;
  assign n9190 = ~n9188 & n9189;
  assign n14020 = n8979 | n8981;
  assign n14063 = n9190 & n14020;
  assign n14064 = n8979 & n9190;
  assign n14065 = (n13933 & n14063) | (n13933 & n14064) | (n14063 & n14064);
  assign n14066 = n9190 | n14020;
  assign n14067 = n8979 | n9190;
  assign n14068 = (n13933 & n14066) | (n13933 & n14067) | (n14066 & n14067);
  assign n9193 = ~n14065 & n14068;
  assign n9194 = x71 & x94;
  assign n9195 = n9193 & n9194;
  assign n9196 = n9193 | n9194;
  assign n9197 = ~n9195 & n9196;
  assign n14069 = n8986 & n9197;
  assign n14070 = (n9197 & n16862) | (n9197 & n14069) | (n16862 & n14069);
  assign n14071 = n8986 | n9197;
  assign n14072 = n16862 | n14071;
  assign n9200 = ~n14070 & n14072;
  assign n9201 = x70 & x95;
  assign n9202 = n9200 & n9201;
  assign n9203 = n9200 | n9201;
  assign n9204 = ~n9202 & n9203;
  assign n14073 = n8993 & n9204;
  assign n14074 = (n9204 & n13983) | (n9204 & n14073) | (n13983 & n14073);
  assign n14075 = n8993 | n9204;
  assign n14076 = n13983 | n14075;
  assign n9207 = ~n14074 & n14076;
  assign n9208 = x69 & x96;
  assign n9209 = n9207 & n9208;
  assign n9210 = n9207 | n9208;
  assign n9211 = ~n9209 & n9210;
  assign n14077 = n9000 & n9211;
  assign n14078 = (n9211 & n13987) | (n9211 & n14077) | (n13987 & n14077);
  assign n14079 = n9000 | n9211;
  assign n14080 = n13987 | n14079;
  assign n9214 = ~n14078 & n14080;
  assign n9215 = x68 & x97;
  assign n9216 = n9214 & n9215;
  assign n9217 = n9214 | n9215;
  assign n9218 = ~n9216 & n9217;
  assign n14081 = n9007 & n9218;
  assign n14082 = (n9218 & n13991) | (n9218 & n14081) | (n13991 & n14081);
  assign n14083 = n9007 | n9218;
  assign n14084 = n13991 | n14083;
  assign n9221 = ~n14082 & n14084;
  assign n9222 = x67 & x98;
  assign n9223 = n9221 & n9222;
  assign n9224 = n9221 | n9222;
  assign n9225 = ~n9223 & n9224;
  assign n14085 = n9014 & n9225;
  assign n14086 = (n9225 & n13995) | (n9225 & n14085) | (n13995 & n14085);
  assign n14087 = n9014 | n9225;
  assign n14088 = n13995 | n14087;
  assign n9228 = ~n14086 & n14088;
  assign n9229 = x66 & x99;
  assign n9230 = n9228 & n9229;
  assign n9231 = n9228 | n9229;
  assign n9232 = ~n9230 & n9231;
  assign n14089 = n9021 & n9232;
  assign n14090 = (n9232 & n14000) | (n9232 & n14089) | (n14000 & n14089);
  assign n14091 = n9021 | n9232;
  assign n14092 = n14000 | n14091;
  assign n9235 = ~n14090 & n14092;
  assign n9236 = x65 & x100;
  assign n9237 = n9235 & n9236;
  assign n9238 = n9235 | n9236;
  assign n9239 = ~n9237 & n9238;
  assign n14018 = n9028 | n9030;
  assign n14093 = n9239 & n14018;
  assign n14094 = n9028 & n9239;
  assign n14095 = (n13928 & n14093) | (n13928 & n14094) | (n14093 & n14094);
  assign n14096 = n9239 | n14018;
  assign n14097 = n9028 | n9239;
  assign n14098 = (n13928 & n14096) | (n13928 & n14097) | (n14096 & n14097);
  assign n9242 = ~n14095 & n14098;
  assign n9243 = x64 & x101;
  assign n9244 = n9242 & n9243;
  assign n9245 = n9242 | n9243;
  assign n9246 = ~n9244 & n9245;
  assign n14016 = n9035 | n9037;
  assign n16926 = n9246 & n14016;
  assign n16927 = n9035 & n9246;
  assign n16928 = (n13926 & n16926) | (n13926 & n16927) | (n16926 & n16927);
  assign n16929 = n9246 | n14016;
  assign n16930 = n9035 | n9246;
  assign n16931 = (n13926 & n16929) | (n13926 & n16930) | (n16929 & n16930);
  assign n9249 = ~n16928 & n16931;
  assign n9250 = x63 & x102;
  assign n9251 = n9249 & n9250;
  assign n9252 = n9249 | n9250;
  assign n9253 = ~n9251 & n9252;
  assign n14014 = n9042 | n9044;
  assign n16932 = n9253 & n14014;
  assign n16933 = n9042 & n9253;
  assign n16934 = (n13924 & n16932) | (n13924 & n16933) | (n16932 & n16933);
  assign n16935 = n9253 | n14014;
  assign n16936 = n9042 | n9253;
  assign n16937 = (n13924 & n16935) | (n13924 & n16936) | (n16935 & n16936);
  assign n9256 = ~n16934 & n16937;
  assign n9257 = x62 & x103;
  assign n9258 = n9256 & n9257;
  assign n9259 = n9256 | n9257;
  assign n9260 = ~n9258 & n9259;
  assign n9261 = n14013 & n9260;
  assign n9262 = n14013 | n9260;
  assign n9263 = ~n9261 & n9262;
  assign n9264 = x61 & x104;
  assign n9265 = n9263 & n9264;
  assign n9266 = n9263 | n9264;
  assign n9267 = ~n9265 & n9266;
  assign n9268 = n14011 & n9267;
  assign n9269 = n14011 | n9267;
  assign n9270 = ~n9268 & n9269;
  assign n9271 = x60 & x105;
  assign n9272 = n9270 & n9271;
  assign n9273 = n9270 | n9271;
  assign n9274 = ~n9272 & n9273;
  assign n9275 = n14009 & n9274;
  assign n9276 = n14009 | n9274;
  assign n9277 = ~n9275 & n9276;
  assign n9278 = x59 & x106;
  assign n9279 = n9277 & n9278;
  assign n9280 = n9277 | n9278;
  assign n9281 = ~n9279 & n9280;
  assign n9282 = n14007 & n9281;
  assign n9283 = n14007 | n9281;
  assign n9284 = ~n9282 & n9283;
  assign n9285 = x58 & x107;
  assign n9286 = n9284 & n9285;
  assign n9287 = n9284 | n9285;
  assign n9288 = ~n9286 & n9287;
  assign n9289 = n14005 & n9288;
  assign n9290 = n14005 | n9288;
  assign n9291 = ~n9289 & n9290;
  assign n9292 = x57 & x108;
  assign n9293 = n9291 & n9292;
  assign n9294 = n9291 | n9292;
  assign n9295 = ~n9293 & n9294;
  assign n9296 = n9114 & n9295;
  assign n9297 = n9114 | n9295;
  assign n9298 = ~n9296 & n9297;
  assign n9299 = x56 & x109;
  assign n9300 = n9298 & n9299;
  assign n9301 = n9298 | n9299;
  assign n9302 = ~n9300 & n9301;
  assign n9303 = n9113 & n9302;
  assign n9304 = n9113 | n9302;
  assign n9305 = ~n9303 & n9304;
  assign n9306 = x55 & x110;
  assign n9307 = n9305 & n9306;
  assign n9308 = n9305 | n9306;
  assign n9309 = ~n9307 & n9308;
  assign n9310 = n9112 & n9309;
  assign n9311 = n9112 | n9309;
  assign n9312 = ~n9310 & n9311;
  assign n9313 = x54 & x111;
  assign n9314 = n9312 & n9313;
  assign n9315 = n9312 | n9313;
  assign n9316 = ~n9314 & n9315;
  assign n9317 = n9111 & n9316;
  assign n9318 = n9111 | n9316;
  assign n9319 = ~n9317 & n9318;
  assign n9320 = n9314 | n9317;
  assign n9321 = n9307 | n9310;
  assign n9322 = n9300 | n9303;
  assign n14099 = n9293 | n9295;
  assign n14100 = (n9114 & n9293) | (n9114 & n14099) | (n9293 & n14099);
  assign n14101 = n9286 | n9288;
  assign n14102 = (n9286 & n14005) | (n9286 & n14101) | (n14005 & n14101);
  assign n14103 = n9279 | n9281;
  assign n14104 = (n9279 & n14007) | (n9279 & n14103) | (n14007 & n14103);
  assign n14105 = n9272 | n9274;
  assign n14106 = (n9272 & n14009) | (n9272 & n14105) | (n14009 & n14105);
  assign n14107 = n9265 | n9267;
  assign n14108 = (n9265 & n14011) | (n9265 & n14107) | (n14011 & n14107);
  assign n14015 = (n9042 & n13924) | (n9042 & n14014) | (n13924 & n14014);
  assign n14017 = (n9035 & n13926) | (n9035 & n14016) | (n13926 & n14016);
  assign n14121 = n9174 | n9176;
  assign n16940 = n8965 | n9174;
  assign n16941 = (n9174 & n9176) | (n9174 & n16940) | (n9176 & n16940);
  assign n16942 = (n13968 & n14121) | (n13968 & n16941) | (n14121 & n16941);
  assign n16943 = (n13969 & n14121) | (n13969 & n16941) | (n14121 & n16941);
  assign n16944 = (n16758 & n16942) | (n16758 & n16943) | (n16942 & n16943);
  assign n14029 = (n13865 & n16884) | (n13865 & n14028) | (n16884 & n14028);
  assign n14126 = n9153 | n9155;
  assign n16945 = n8944 | n9153;
  assign n16946 = (n9153 & n9155) | (n9153 & n16945) | (n9155 & n16945);
  assign n16947 = (n13959 & n14126) | (n13959 & n16946) | (n14126 & n16946);
  assign n16948 = (n13958 & n14126) | (n13958 & n16946) | (n14126 & n16946);
  assign n16949 = (n13835 & n16947) | (n13835 & n16948) | (n16947 & n16948);
  assign n16950 = n8937 | n9146;
  assign n16951 = (n9146 & n9148) | (n9146 & n16950) | (n9148 & n16950);
  assign n14129 = n9146 | n14043;
  assign n14130 = (n16817 & n16951) | (n16817 & n14129) | (n16951 & n14129);
  assign n9346 = x79 & x87;
  assign n16952 = n9346 & n16899;
  assign n16953 = (n9141 & n9346) | (n9141 & n16952) | (n9346 & n16952);
  assign n14134 = n9346 & n16899;
  assign n14135 = (n16891 & n16953) | (n16891 & n14134) | (n16953 & n14134);
  assign n16954 = n9346 | n16899;
  assign n16955 = n9141 | n16954;
  assign n14137 = n9346 | n16899;
  assign n14138 = (n16891 & n16955) | (n16891 & n14137) | (n16955 & n14137);
  assign n9349 = ~n14135 & n14138;
  assign n9350 = n14130 & n9349;
  assign n9351 = n14130 | n9349;
  assign n9352 = ~n9350 & n9351;
  assign n9353 = x78 & x88;
  assign n9354 = n9352 & n9353;
  assign n9355 = n9352 | n9353;
  assign n9356 = ~n9354 & n9355;
  assign n9357 = n16949 & n9356;
  assign n9358 = n16949 | n9356;
  assign n9359 = ~n9357 & n9358;
  assign n9360 = x77 & x89;
  assign n9361 = n9359 & n9360;
  assign n9362 = n9359 | n9360;
  assign n9363 = ~n9361 & n9362;
  assign n14123 = n9160 | n9162;
  assign n14139 = n9363 & n14123;
  assign n14140 = n9160 & n9363;
  assign n14141 = (n14029 & n14139) | (n14029 & n14140) | (n14139 & n14140);
  assign n14142 = n9363 | n14123;
  assign n14143 = n9160 | n9363;
  assign n14144 = (n14029 & n14142) | (n14029 & n14143) | (n14142 & n14143);
  assign n9366 = ~n14141 & n14144;
  assign n9367 = x76 & x90;
  assign n9368 = n9366 & n9367;
  assign n9369 = n9366 | n9367;
  assign n9370 = ~n9368 & n9369;
  assign n14145 = n9167 & n9370;
  assign n16956 = (n9370 & n14053) | (n9370 & n14145) | (n14053 & n14145);
  assign n16957 = (n9370 & n14054) | (n9370 & n14145) | (n14054 & n14145);
  assign n16958 = (n13938 & n16956) | (n13938 & n16957) | (n16956 & n16957);
  assign n14147 = n9167 | n9370;
  assign n16959 = n14053 | n14147;
  assign n16960 = n14054 | n14147;
  assign n16961 = (n13938 & n16959) | (n13938 & n16960) | (n16959 & n16960);
  assign n9373 = ~n16958 & n16961;
  assign n9374 = x75 & x91;
  assign n9375 = n9373 & n9374;
  assign n9376 = n9373 | n9374;
  assign n9377 = ~n9375 & n9376;
  assign n9378 = n16944 & n9377;
  assign n9379 = n16944 | n9377;
  assign n9380 = ~n9378 & n9379;
  assign n9381 = x74 & x92;
  assign n9382 = n9380 & n9381;
  assign n9383 = n9380 | n9381;
  assign n9384 = ~n9382 & n9383;
  assign n14118 = n9181 | n9183;
  assign n14149 = n9384 & n14118;
  assign n14150 = n9181 & n9384;
  assign n14151 = (n16882 & n14149) | (n16882 & n14150) | (n14149 & n14150);
  assign n14152 = n9384 | n14118;
  assign n14153 = n9181 | n9384;
  assign n14154 = (n16882 & n14152) | (n16882 & n14153) | (n14152 & n14153);
  assign n9387 = ~n14151 & n14154;
  assign n9388 = x73 & x93;
  assign n9389 = n9387 & n9388;
  assign n9390 = n9387 | n9388;
  assign n9391 = ~n9389 & n9390;
  assign n14155 = n9188 & n9391;
  assign n16962 = (n9391 & n14064) | (n9391 & n14155) | (n14064 & n14155);
  assign n16963 = (n9391 & n14063) | (n9391 & n14155) | (n14063 & n14155);
  assign n16964 = (n13933 & n16962) | (n13933 & n16963) | (n16962 & n16963);
  assign n14157 = n9188 | n9391;
  assign n16965 = n14064 | n14157;
  assign n16966 = n14063 | n14157;
  assign n16967 = (n13933 & n16965) | (n13933 & n16966) | (n16965 & n16966);
  assign n9394 = ~n16964 & n16967;
  assign n9395 = x72 & x94;
  assign n9396 = n9394 & n9395;
  assign n9397 = n9394 | n9395;
  assign n9398 = ~n9396 & n9397;
  assign n14116 = n9195 | n9197;
  assign n16968 = n9398 & n14116;
  assign n16938 = n8986 | n9195;
  assign n16939 = (n9195 & n9197) | (n9195 & n16938) | (n9197 & n16938);
  assign n16969 = n9398 & n16939;
  assign n16970 = (n16862 & n16968) | (n16862 & n16969) | (n16968 & n16969);
  assign n16971 = n9398 | n14116;
  assign n16972 = n9398 | n16939;
  assign n16973 = (n16862 & n16971) | (n16862 & n16972) | (n16971 & n16972);
  assign n9401 = ~n16970 & n16973;
  assign n9402 = x71 & x95;
  assign n9403 = n9401 & n9402;
  assign n9404 = n9401 | n9402;
  assign n9405 = ~n9403 & n9404;
  assign n14159 = n9202 & n9405;
  assign n16974 = (n9405 & n14073) | (n9405 & n14159) | (n14073 & n14159);
  assign n16975 = (n9204 & n9405) | (n9204 & n14159) | (n9405 & n14159);
  assign n16976 = (n13983 & n16974) | (n13983 & n16975) | (n16974 & n16975);
  assign n14161 = n9202 | n9405;
  assign n16977 = n14073 | n14161;
  assign n16978 = n9204 | n14161;
  assign n16979 = (n13983 & n16977) | (n13983 & n16978) | (n16977 & n16978);
  assign n9408 = ~n16976 & n16979;
  assign n9409 = x70 & x96;
  assign n9410 = n9408 & n9409;
  assign n9411 = n9408 | n9409;
  assign n9412 = ~n9410 & n9411;
  assign n14163 = n9209 & n9412;
  assign n14164 = (n9412 & n14078) | (n9412 & n14163) | (n14078 & n14163);
  assign n14165 = n9209 | n9412;
  assign n14166 = n14078 | n14165;
  assign n9415 = ~n14164 & n14166;
  assign n9416 = x69 & x97;
  assign n9417 = n9415 & n9416;
  assign n9418 = n9415 | n9416;
  assign n9419 = ~n9417 & n9418;
  assign n14167 = n9216 & n9419;
  assign n14168 = (n9419 & n14082) | (n9419 & n14167) | (n14082 & n14167);
  assign n14169 = n9216 | n9419;
  assign n14170 = n14082 | n14169;
  assign n9422 = ~n14168 & n14170;
  assign n9423 = x68 & x98;
  assign n9424 = n9422 & n9423;
  assign n9425 = n9422 | n9423;
  assign n9426 = ~n9424 & n9425;
  assign n14171 = n9223 & n9426;
  assign n14172 = (n9426 & n14086) | (n9426 & n14171) | (n14086 & n14171);
  assign n14173 = n9223 | n9426;
  assign n14174 = n14086 | n14173;
  assign n9429 = ~n14172 & n14174;
  assign n9430 = x67 & x99;
  assign n9431 = n9429 & n9430;
  assign n9432 = n9429 | n9430;
  assign n9433 = ~n9431 & n9432;
  assign n14175 = n9230 & n9433;
  assign n14176 = (n9433 & n14090) | (n9433 & n14175) | (n14090 & n14175);
  assign n14177 = n9230 | n9433;
  assign n14178 = n14090 | n14177;
  assign n9436 = ~n14176 & n14178;
  assign n9437 = x66 & x100;
  assign n9438 = n9436 & n9437;
  assign n9439 = n9436 | n9437;
  assign n9440 = ~n9438 & n9439;
  assign n14179 = n9237 & n9440;
  assign n14180 = (n9440 & n14095) | (n9440 & n14179) | (n14095 & n14179);
  assign n14181 = n9237 | n9440;
  assign n14182 = n14095 | n14181;
  assign n9443 = ~n14180 & n14182;
  assign n9444 = x65 & x101;
  assign n9445 = n9443 & n9444;
  assign n9446 = n9443 | n9444;
  assign n9447 = ~n9445 & n9446;
  assign n14113 = n9244 | n9246;
  assign n14183 = n9447 & n14113;
  assign n14184 = n9244 & n9447;
  assign n14185 = (n14017 & n14183) | (n14017 & n14184) | (n14183 & n14184);
  assign n14186 = n9447 | n14113;
  assign n14187 = n9244 | n9447;
  assign n14188 = (n14017 & n14186) | (n14017 & n14187) | (n14186 & n14187);
  assign n9450 = ~n14185 & n14188;
  assign n9451 = x64 & x102;
  assign n9452 = n9450 & n9451;
  assign n9453 = n9450 | n9451;
  assign n9454 = ~n9452 & n9453;
  assign n14111 = n9251 | n9253;
  assign n16980 = n9454 & n14111;
  assign n16981 = n9251 & n9454;
  assign n16982 = (n14015 & n16980) | (n14015 & n16981) | (n16980 & n16981);
  assign n16983 = n9454 | n14111;
  assign n16984 = n9251 | n9454;
  assign n16985 = (n14015 & n16983) | (n14015 & n16984) | (n16983 & n16984);
  assign n9457 = ~n16982 & n16985;
  assign n9458 = x63 & x103;
  assign n9459 = n9457 & n9458;
  assign n9460 = n9457 | n9458;
  assign n9461 = ~n9459 & n9460;
  assign n14109 = n9258 | n9260;
  assign n16986 = n9461 & n14109;
  assign n16987 = n9258 & n9461;
  assign n16988 = (n14013 & n16986) | (n14013 & n16987) | (n16986 & n16987);
  assign n16989 = n9461 | n14109;
  assign n16990 = n9258 | n9461;
  assign n16991 = (n14013 & n16989) | (n14013 & n16990) | (n16989 & n16990);
  assign n9464 = ~n16988 & n16991;
  assign n9465 = x62 & x104;
  assign n9466 = n9464 & n9465;
  assign n9467 = n9464 | n9465;
  assign n9468 = ~n9466 & n9467;
  assign n9469 = n14108 & n9468;
  assign n9470 = n14108 | n9468;
  assign n9471 = ~n9469 & n9470;
  assign n9472 = x61 & x105;
  assign n9473 = n9471 & n9472;
  assign n9474 = n9471 | n9472;
  assign n9475 = ~n9473 & n9474;
  assign n9476 = n14106 & n9475;
  assign n9477 = n14106 | n9475;
  assign n9478 = ~n9476 & n9477;
  assign n9479 = x60 & x106;
  assign n9480 = n9478 & n9479;
  assign n9481 = n9478 | n9479;
  assign n9482 = ~n9480 & n9481;
  assign n9483 = n14104 & n9482;
  assign n9484 = n14104 | n9482;
  assign n9485 = ~n9483 & n9484;
  assign n9486 = x59 & x107;
  assign n9487 = n9485 & n9486;
  assign n9488 = n9485 | n9486;
  assign n9489 = ~n9487 & n9488;
  assign n9490 = n14102 & n9489;
  assign n9491 = n14102 | n9489;
  assign n9492 = ~n9490 & n9491;
  assign n9493 = x58 & x108;
  assign n9494 = n9492 & n9493;
  assign n9495 = n9492 | n9493;
  assign n9496 = ~n9494 & n9495;
  assign n9497 = n14100 & n9496;
  assign n9498 = n14100 | n9496;
  assign n9499 = ~n9497 & n9498;
  assign n9500 = x57 & x109;
  assign n9501 = n9499 & n9500;
  assign n9502 = n9499 | n9500;
  assign n9503 = ~n9501 & n9502;
  assign n9504 = n9322 & n9503;
  assign n9505 = n9322 | n9503;
  assign n9506 = ~n9504 & n9505;
  assign n9507 = x56 & x110;
  assign n9508 = n9506 & n9507;
  assign n9509 = n9506 | n9507;
  assign n9510 = ~n9508 & n9509;
  assign n9511 = n9321 & n9510;
  assign n9512 = n9321 | n9510;
  assign n9513 = ~n9511 & n9512;
  assign n9514 = x55 & x111;
  assign n9515 = n9513 & n9514;
  assign n9516 = n9513 | n9514;
  assign n9517 = ~n9515 & n9516;
  assign n9518 = n9320 & n9517;
  assign n9519 = n9320 | n9517;
  assign n9520 = ~n9518 & n9519;
  assign n9521 = n9515 | n9518;
  assign n9522 = n9508 | n9511;
  assign n14189 = n9501 | n9503;
  assign n14190 = (n9322 & n9501) | (n9322 & n14189) | (n9501 & n14189);
  assign n14191 = n9494 | n9496;
  assign n14192 = (n9494 & n14100) | (n9494 & n14191) | (n14100 & n14191);
  assign n14193 = n9487 | n9489;
  assign n14194 = (n9487 & n14102) | (n9487 & n14193) | (n14102 & n14193);
  assign n14195 = n9480 | n9482;
  assign n14196 = (n9480 & n14104) | (n9480 & n14195) | (n14104 & n14195);
  assign n14197 = n9473 | n9475;
  assign n14198 = (n9473 & n14106) | (n9473 & n14197) | (n14106 & n14197);
  assign n14110 = (n9258 & n14013) | (n9258 & n14109) | (n14013 & n14109);
  assign n14112 = (n9251 & n14015) | (n9251 & n14111) | (n14015 & n14111);
  assign n14117 = (n16862 & n16939) | (n16862 & n14116) | (n16939 & n14116);
  assign n14208 = n9389 | n9391;
  assign n16992 = n9188 | n9389;
  assign n16993 = (n9389 & n9391) | (n9389 & n16992) | (n9391 & n16992);
  assign n16994 = (n14064 & n14208) | (n14064 & n16993) | (n14208 & n16993);
  assign n16995 = (n14063 & n14208) | (n14063 & n16993) | (n14208 & n16993);
  assign n16996 = (n13933 & n16994) | (n13933 & n16995) | (n16994 & n16995);
  assign n14213 = n9368 | n9370;
  assign n16997 = n9167 | n9368;
  assign n16998 = (n9368 & n9370) | (n9368 & n16997) | (n9370 & n16997);
  assign n16999 = (n14053 & n14213) | (n14053 & n16998) | (n14213 & n16998);
  assign n17000 = (n14054 & n14213) | (n14054 & n16998) | (n14213 & n16998);
  assign n17001 = (n13938 & n16999) | (n13938 & n17000) | (n16999 & n17000);
  assign n9546 = x79 & x88;
  assign n17003 = n9546 & n16953;
  assign n17825 = n9346 & n9546;
  assign n17826 = n16899 & n17825;
  assign n17005 = (n16891 & n17003) | (n16891 & n17826) | (n17003 & n17826);
  assign n17002 = (n9349 & n9546) | (n9349 & n17005) | (n9546 & n17005);
  assign n14221 = (n14130 & n17002) | (n14130 & n17005) | (n17002 & n17005);
  assign n17007 = n9546 | n16953;
  assign n17827 = n9346 | n9546;
  assign n17828 = (n9546 & n16899) | (n9546 & n17827) | (n16899 & n17827);
  assign n17009 = (n16891 & n17007) | (n16891 & n17828) | (n17007 & n17828);
  assign n17006 = n9349 | n17009;
  assign n14224 = (n14130 & n17006) | (n14130 & n17009) | (n17006 & n17009);
  assign n9549 = ~n14221 & n14224;
  assign n14226 = n9354 & n9549;
  assign n17010 = (n9356 & n9549) | (n9356 & n14226) | (n9549 & n14226);
  assign n14227 = (n16949 & n17010) | (n16949 & n14226) | (n17010 & n14226);
  assign n14229 = n9354 | n9549;
  assign n17011 = n9356 | n14229;
  assign n14230 = (n16949 & n17011) | (n16949 & n14229) | (n17011 & n14229);
  assign n9552 = ~n14227 & n14230;
  assign n9553 = x78 & x89;
  assign n9554 = n9552 & n9553;
  assign n9555 = n9552 | n9553;
  assign n9556 = ~n9554 & n9555;
  assign n14231 = n9361 & n9556;
  assign n17012 = (n9556 & n14140) | (n9556 & n14231) | (n14140 & n14231);
  assign n17013 = (n9556 & n14139) | (n9556 & n14231) | (n14139 & n14231);
  assign n17014 = (n14029 & n17012) | (n14029 & n17013) | (n17012 & n17013);
  assign n14233 = n9361 | n9556;
  assign n17015 = n14140 | n14233;
  assign n17016 = n14139 | n14233;
  assign n17017 = (n14029 & n17015) | (n14029 & n17016) | (n17015 & n17016);
  assign n9559 = ~n17014 & n17017;
  assign n9560 = x77 & x90;
  assign n9561 = n9559 & n9560;
  assign n9562 = n9559 | n9560;
  assign n9563 = ~n9561 & n9562;
  assign n9564 = n17001 & n9563;
  assign n9565 = n17001 | n9563;
  assign n9566 = ~n9564 & n9565;
  assign n9567 = x76 & x91;
  assign n9568 = n9566 & n9567;
  assign n9569 = n9566 | n9567;
  assign n9570 = ~n9568 & n9569;
  assign n14210 = n9375 | n9377;
  assign n14235 = n9570 & n14210;
  assign n14236 = n9375 & n9570;
  assign n14237 = (n16944 & n14235) | (n16944 & n14236) | (n14235 & n14236);
  assign n14238 = n9570 | n14210;
  assign n14239 = n9375 | n9570;
  assign n14240 = (n16944 & n14238) | (n16944 & n14239) | (n14238 & n14239);
  assign n9573 = ~n14237 & n14240;
  assign n9574 = x75 & x92;
  assign n9575 = n9573 & n9574;
  assign n9576 = n9573 | n9574;
  assign n9577 = ~n9575 & n9576;
  assign n14241 = n9382 & n9577;
  assign n17018 = (n9577 & n14150) | (n9577 & n14241) | (n14150 & n14241);
  assign n17019 = (n9577 & n14149) | (n9577 & n14241) | (n14149 & n14241);
  assign n17020 = (n16882 & n17018) | (n16882 & n17019) | (n17018 & n17019);
  assign n14243 = n9382 | n9577;
  assign n17021 = n14150 | n14243;
  assign n17022 = n14149 | n14243;
  assign n17023 = (n16882 & n17021) | (n16882 & n17022) | (n17021 & n17022);
  assign n9580 = ~n17020 & n17023;
  assign n9581 = x74 & x93;
  assign n9582 = n9580 & n9581;
  assign n9583 = n9580 | n9581;
  assign n9584 = ~n9582 & n9583;
  assign n9585 = n16996 & n9584;
  assign n9586 = n16996 | n9584;
  assign n9587 = ~n9585 & n9586;
  assign n9588 = x73 & x94;
  assign n9589 = n9587 & n9588;
  assign n9590 = n9587 | n9588;
  assign n9591 = ~n9589 & n9590;
  assign n14205 = n9396 | n9398;
  assign n14245 = n9591 & n14205;
  assign n14246 = n9396 & n9591;
  assign n14247 = (n14117 & n14245) | (n14117 & n14246) | (n14245 & n14246);
  assign n14248 = n9591 | n14205;
  assign n14249 = n9396 | n9591;
  assign n14250 = (n14117 & n14248) | (n14117 & n14249) | (n14248 & n14249);
  assign n9594 = ~n14247 & n14250;
  assign n9595 = x72 & x95;
  assign n9596 = n9594 & n9595;
  assign n9597 = n9594 | n9595;
  assign n9598 = ~n9596 & n9597;
  assign n14251 = n9403 & n9598;
  assign n14252 = (n9598 & n16976) | (n9598 & n14251) | (n16976 & n14251);
  assign n14253 = n9403 | n9598;
  assign n14254 = n16976 | n14253;
  assign n9601 = ~n14252 & n14254;
  assign n9602 = x71 & x96;
  assign n9603 = n9601 & n9602;
  assign n9604 = n9601 | n9602;
  assign n9605 = ~n9603 & n9604;
  assign n14255 = n9410 & n9605;
  assign n14256 = (n9605 & n14164) | (n9605 & n14255) | (n14164 & n14255);
  assign n14257 = n9410 | n9605;
  assign n14258 = n14164 | n14257;
  assign n9608 = ~n14256 & n14258;
  assign n9609 = x70 & x97;
  assign n9610 = n9608 & n9609;
  assign n9611 = n9608 | n9609;
  assign n9612 = ~n9610 & n9611;
  assign n14259 = n9417 & n9612;
  assign n14260 = (n9612 & n14168) | (n9612 & n14259) | (n14168 & n14259);
  assign n14261 = n9417 | n9612;
  assign n14262 = n14168 | n14261;
  assign n9615 = ~n14260 & n14262;
  assign n9616 = x69 & x98;
  assign n9617 = n9615 & n9616;
  assign n9618 = n9615 | n9616;
  assign n9619 = ~n9617 & n9618;
  assign n14263 = n9424 & n9619;
  assign n14264 = (n9619 & n14172) | (n9619 & n14263) | (n14172 & n14263);
  assign n14265 = n9424 | n9619;
  assign n14266 = n14172 | n14265;
  assign n9622 = ~n14264 & n14266;
  assign n9623 = x68 & x99;
  assign n9624 = n9622 & n9623;
  assign n9625 = n9622 | n9623;
  assign n9626 = ~n9624 & n9625;
  assign n14267 = n9431 & n9626;
  assign n14268 = (n9626 & n14176) | (n9626 & n14267) | (n14176 & n14267);
  assign n14269 = n9431 | n9626;
  assign n14270 = n14176 | n14269;
  assign n9629 = ~n14268 & n14270;
  assign n9630 = x67 & x100;
  assign n9631 = n9629 & n9630;
  assign n9632 = n9629 | n9630;
  assign n9633 = ~n9631 & n9632;
  assign n14271 = n9438 & n9633;
  assign n14272 = (n9633 & n14180) | (n9633 & n14271) | (n14180 & n14271);
  assign n14273 = n9438 | n9633;
  assign n14274 = n14180 | n14273;
  assign n9636 = ~n14272 & n14274;
  assign n9637 = x66 & x101;
  assign n9638 = n9636 & n9637;
  assign n9639 = n9636 | n9637;
  assign n9640 = ~n9638 & n9639;
  assign n14275 = n9445 & n9640;
  assign n14276 = (n9640 & n14185) | (n9640 & n14275) | (n14185 & n14275);
  assign n14277 = n9445 | n9640;
  assign n14278 = n14185 | n14277;
  assign n9643 = ~n14276 & n14278;
  assign n9644 = x65 & x102;
  assign n9645 = n9643 & n9644;
  assign n9646 = n9643 | n9644;
  assign n9647 = ~n9645 & n9646;
  assign n14203 = n9452 | n9454;
  assign n14279 = n9647 & n14203;
  assign n14280 = n9452 & n9647;
  assign n14281 = (n14112 & n14279) | (n14112 & n14280) | (n14279 & n14280);
  assign n14282 = n9647 | n14203;
  assign n14283 = n9452 | n9647;
  assign n14284 = (n14112 & n14282) | (n14112 & n14283) | (n14282 & n14283);
  assign n9650 = ~n14281 & n14284;
  assign n9651 = x64 & x103;
  assign n9652 = n9650 & n9651;
  assign n9653 = n9650 | n9651;
  assign n9654 = ~n9652 & n9653;
  assign n14201 = n9459 | n9461;
  assign n17024 = n9654 & n14201;
  assign n17025 = n9459 & n9654;
  assign n17026 = (n14110 & n17024) | (n14110 & n17025) | (n17024 & n17025);
  assign n17027 = n9654 | n14201;
  assign n17028 = n9459 | n9654;
  assign n17029 = (n14110 & n17027) | (n14110 & n17028) | (n17027 & n17028);
  assign n9657 = ~n17026 & n17029;
  assign n9658 = x63 & x104;
  assign n9659 = n9657 & n9658;
  assign n9660 = n9657 | n9658;
  assign n9661 = ~n9659 & n9660;
  assign n14199 = n9466 | n9468;
  assign n17030 = n9661 & n14199;
  assign n17031 = n9466 & n9661;
  assign n17032 = (n14108 & n17030) | (n14108 & n17031) | (n17030 & n17031);
  assign n17033 = n9661 | n14199;
  assign n17034 = n9466 | n9661;
  assign n17035 = (n14108 & n17033) | (n14108 & n17034) | (n17033 & n17034);
  assign n9664 = ~n17032 & n17035;
  assign n9665 = x62 & x105;
  assign n9666 = n9664 & n9665;
  assign n9667 = n9664 | n9665;
  assign n9668 = ~n9666 & n9667;
  assign n9669 = n14198 & n9668;
  assign n9670 = n14198 | n9668;
  assign n9671 = ~n9669 & n9670;
  assign n9672 = x61 & x106;
  assign n9673 = n9671 & n9672;
  assign n9674 = n9671 | n9672;
  assign n9675 = ~n9673 & n9674;
  assign n9676 = n14196 & n9675;
  assign n9677 = n14196 | n9675;
  assign n9678 = ~n9676 & n9677;
  assign n9679 = x60 & x107;
  assign n9680 = n9678 & n9679;
  assign n9681 = n9678 | n9679;
  assign n9682 = ~n9680 & n9681;
  assign n9683 = n14194 & n9682;
  assign n9684 = n14194 | n9682;
  assign n9685 = ~n9683 & n9684;
  assign n9686 = x59 & x108;
  assign n9687 = n9685 & n9686;
  assign n9688 = n9685 | n9686;
  assign n9689 = ~n9687 & n9688;
  assign n9690 = n14192 & n9689;
  assign n9691 = n14192 | n9689;
  assign n9692 = ~n9690 & n9691;
  assign n9693 = x58 & x109;
  assign n9694 = n9692 & n9693;
  assign n9695 = n9692 | n9693;
  assign n9696 = ~n9694 & n9695;
  assign n9697 = n14190 & n9696;
  assign n9698 = n14190 | n9696;
  assign n9699 = ~n9697 & n9698;
  assign n9700 = x57 & x110;
  assign n9701 = n9699 & n9700;
  assign n9702 = n9699 | n9700;
  assign n9703 = ~n9701 & n9702;
  assign n9704 = n9522 & n9703;
  assign n9705 = n9522 | n9703;
  assign n9706 = ~n9704 & n9705;
  assign n9707 = x56 & x111;
  assign n9708 = n9706 & n9707;
  assign n9709 = n9706 | n9707;
  assign n9710 = ~n9708 & n9709;
  assign n9711 = n9521 & n9710;
  assign n9712 = n9521 | n9710;
  assign n9713 = ~n9711 & n9712;
  assign n9714 = n9708 | n9711;
  assign n14285 = n9701 | n9703;
  assign n14286 = (n9522 & n9701) | (n9522 & n14285) | (n9701 & n14285);
  assign n14287 = n9694 | n9696;
  assign n14288 = (n9694 & n14190) | (n9694 & n14287) | (n14190 & n14287);
  assign n14289 = n9687 | n9689;
  assign n14290 = (n9687 & n14192) | (n9687 & n14289) | (n14192 & n14289);
  assign n14291 = n9680 | n9682;
  assign n14292 = (n9680 & n14194) | (n9680 & n14291) | (n14194 & n14291);
  assign n14293 = n9673 | n9675;
  assign n14294 = (n9673 & n14196) | (n9673 & n14293) | (n14196 & n14293);
  assign n14200 = (n9466 & n14108) | (n9466 & n14199) | (n14108 & n14199);
  assign n14202 = (n9459 & n14110) | (n9459 & n14201) | (n14110 & n14201);
  assign n14307 = n9575 | n9577;
  assign n17038 = n9382 | n9575;
  assign n17039 = (n9575 & n9577) | (n9575 & n17038) | (n9577 & n17038);
  assign n17040 = (n14150 & n14307) | (n14150 & n17039) | (n14307 & n17039);
  assign n17041 = (n14149 & n14307) | (n14149 & n17039) | (n14307 & n17039);
  assign n17042 = (n16882 & n17040) | (n16882 & n17041) | (n17040 & n17041);
  assign n14312 = n9554 | n9556;
  assign n17043 = n9361 | n9554;
  assign n17044 = (n9554 & n9556) | (n9554 & n17043) | (n9556 & n17043);
  assign n17045 = (n14140 & n14312) | (n14140 & n17044) | (n14312 & n17044);
  assign n17046 = (n14139 & n14312) | (n14139 & n17044) | (n14312 & n17044);
  assign n17047 = (n14029 & n17045) | (n14029 & n17046) | (n17045 & n17046);
  assign n9738 = x79 & x89;
  assign n17831 = n9738 & n17003;
  assign n17832 = n9738 & n17826;
  assign n17833 = (n16891 & n17831) | (n16891 & n17832) | (n17831 & n17832);
  assign n17829 = n9546 & n9738;
  assign n17830 = (n9349 & n17833) | (n9349 & n17829) | (n17833 & n17829);
  assign n17050 = (n14130 & n17830) | (n14130 & n17833) | (n17830 & n17833);
  assign n17051 = (n9738 & n17010) | (n9738 & n17050) | (n17010 & n17050);
  assign n17834 = (n9549 & n9738) | (n9549 & n17050) | (n9738 & n17050);
  assign n17835 = n9738 & n17050;
  assign n17836 = (n9354 & n17834) | (n9354 & n17835) | (n17834 & n17835);
  assign n17053 = (n16949 & n17051) | (n16949 & n17836) | (n17051 & n17836);
  assign n17839 = n9738 | n17003;
  assign n17840 = n9738 | n17826;
  assign n17841 = (n16891 & n17839) | (n16891 & n17840) | (n17839 & n17840);
  assign n17837 = n9546 | n9738;
  assign n17838 = (n9349 & n17841) | (n9349 & n17837) | (n17841 & n17837);
  assign n17056 = (n14130 & n17838) | (n14130 & n17841) | (n17838 & n17841);
  assign n17057 = n17010 | n17056;
  assign n17842 = n9549 | n17056;
  assign n17843 = (n9354 & n17056) | (n9354 & n17842) | (n17056 & n17842);
  assign n17059 = (n16949 & n17057) | (n16949 & n17843) | (n17057 & n17843);
  assign n9741 = ~n17053 & n17059;
  assign n9742 = n17047 & n9741;
  assign n9743 = n17047 | n9741;
  assign n9744 = ~n9742 & n9743;
  assign n9745 = x78 & x90;
  assign n9746 = n9744 & n9745;
  assign n9747 = n9744 | n9745;
  assign n9748 = ~n9746 & n9747;
  assign n14309 = n9561 | n9563;
  assign n14318 = n9748 & n14309;
  assign n14319 = n9561 & n9748;
  assign n14320 = (n17001 & n14318) | (n17001 & n14319) | (n14318 & n14319);
  assign n14321 = n9748 | n14309;
  assign n14322 = n9561 | n9748;
  assign n14323 = (n17001 & n14321) | (n17001 & n14322) | (n14321 & n14322);
  assign n9751 = ~n14320 & n14323;
  assign n9752 = x77 & x91;
  assign n9753 = n9751 & n9752;
  assign n9754 = n9751 | n9752;
  assign n9755 = ~n9753 & n9754;
  assign n14324 = n9568 & n9755;
  assign n17060 = (n9755 & n14236) | (n9755 & n14324) | (n14236 & n14324);
  assign n17061 = (n9755 & n14235) | (n9755 & n14324) | (n14235 & n14324);
  assign n17062 = (n16944 & n17060) | (n16944 & n17061) | (n17060 & n17061);
  assign n14326 = n9568 | n9755;
  assign n17063 = n14236 | n14326;
  assign n17064 = n14235 | n14326;
  assign n17065 = (n16944 & n17063) | (n16944 & n17064) | (n17063 & n17064);
  assign n9758 = ~n17062 & n17065;
  assign n9759 = x76 & x92;
  assign n9760 = n9758 & n9759;
  assign n9761 = n9758 | n9759;
  assign n9762 = ~n9760 & n9761;
  assign n9763 = n17042 & n9762;
  assign n9764 = n17042 | n9762;
  assign n9765 = ~n9763 & n9764;
  assign n9766 = x75 & x93;
  assign n9767 = n9765 & n9766;
  assign n9768 = n9765 | n9766;
  assign n9769 = ~n9767 & n9768;
  assign n14304 = n9582 | n9584;
  assign n14328 = n9769 & n14304;
  assign n14329 = n9582 & n9769;
  assign n14330 = (n16996 & n14328) | (n16996 & n14329) | (n14328 & n14329);
  assign n14331 = n9769 | n14304;
  assign n14332 = n9582 | n9769;
  assign n14333 = (n16996 & n14331) | (n16996 & n14332) | (n14331 & n14332);
  assign n9772 = ~n14330 & n14333;
  assign n9773 = x74 & x94;
  assign n9774 = n9772 & n9773;
  assign n9775 = n9772 | n9773;
  assign n9776 = ~n9774 & n9775;
  assign n14334 = n9589 & n9776;
  assign n17066 = (n9776 & n14246) | (n9776 & n14334) | (n14246 & n14334);
  assign n17067 = (n9776 & n14245) | (n9776 & n14334) | (n14245 & n14334);
  assign n17068 = (n14117 & n17066) | (n14117 & n17067) | (n17066 & n17067);
  assign n14336 = n9589 | n9776;
  assign n17069 = n14246 | n14336;
  assign n17070 = n14245 | n14336;
  assign n17071 = (n14117 & n17069) | (n14117 & n17070) | (n17069 & n17070);
  assign n9779 = ~n17068 & n17071;
  assign n9780 = x73 & x95;
  assign n9781 = n9779 & n9780;
  assign n9782 = n9779 | n9780;
  assign n9783 = ~n9781 & n9782;
  assign n14302 = n9596 | n9598;
  assign n17072 = n9783 & n14302;
  assign n17036 = n9403 | n9596;
  assign n17037 = (n9596 & n9598) | (n9596 & n17036) | (n9598 & n17036);
  assign n17073 = n9783 & n17037;
  assign n17074 = (n16976 & n17072) | (n16976 & n17073) | (n17072 & n17073);
  assign n17075 = n9783 | n14302;
  assign n17076 = n9783 | n17037;
  assign n17077 = (n16976 & n17075) | (n16976 & n17076) | (n17075 & n17076);
  assign n9786 = ~n17074 & n17077;
  assign n9787 = x72 & x96;
  assign n9788 = n9786 & n9787;
  assign n9789 = n9786 | n9787;
  assign n9790 = ~n9788 & n9789;
  assign n14338 = n9603 & n9790;
  assign n17078 = (n9790 & n14255) | (n9790 & n14338) | (n14255 & n14338);
  assign n17079 = (n9605 & n9790) | (n9605 & n14338) | (n9790 & n14338);
  assign n17080 = (n14164 & n17078) | (n14164 & n17079) | (n17078 & n17079);
  assign n14340 = n9603 | n9790;
  assign n17081 = n14255 | n14340;
  assign n17082 = n9605 | n14340;
  assign n17083 = (n14164 & n17081) | (n14164 & n17082) | (n17081 & n17082);
  assign n9793 = ~n17080 & n17083;
  assign n9794 = x71 & x97;
  assign n9795 = n9793 & n9794;
  assign n9796 = n9793 | n9794;
  assign n9797 = ~n9795 & n9796;
  assign n14342 = n9610 & n9797;
  assign n14343 = (n9797 & n14260) | (n9797 & n14342) | (n14260 & n14342);
  assign n14344 = n9610 | n9797;
  assign n14345 = n14260 | n14344;
  assign n9800 = ~n14343 & n14345;
  assign n9801 = x70 & x98;
  assign n9802 = n9800 & n9801;
  assign n9803 = n9800 | n9801;
  assign n9804 = ~n9802 & n9803;
  assign n14346 = n9617 & n9804;
  assign n14347 = (n9804 & n14264) | (n9804 & n14346) | (n14264 & n14346);
  assign n14348 = n9617 | n9804;
  assign n14349 = n14264 | n14348;
  assign n9807 = ~n14347 & n14349;
  assign n9808 = x69 & x99;
  assign n9809 = n9807 & n9808;
  assign n9810 = n9807 | n9808;
  assign n9811 = ~n9809 & n9810;
  assign n14350 = n9624 & n9811;
  assign n14351 = (n9811 & n14268) | (n9811 & n14350) | (n14268 & n14350);
  assign n14352 = n9624 | n9811;
  assign n14353 = n14268 | n14352;
  assign n9814 = ~n14351 & n14353;
  assign n9815 = x68 & x100;
  assign n9816 = n9814 & n9815;
  assign n9817 = n9814 | n9815;
  assign n9818 = ~n9816 & n9817;
  assign n14354 = n9631 & n9818;
  assign n14355 = (n9818 & n14272) | (n9818 & n14354) | (n14272 & n14354);
  assign n14356 = n9631 | n9818;
  assign n14357 = n14272 | n14356;
  assign n9821 = ~n14355 & n14357;
  assign n9822 = x67 & x101;
  assign n9823 = n9821 & n9822;
  assign n9824 = n9821 | n9822;
  assign n9825 = ~n9823 & n9824;
  assign n14358 = n9638 & n9825;
  assign n14359 = (n9825 & n14276) | (n9825 & n14358) | (n14276 & n14358);
  assign n14360 = n9638 | n9825;
  assign n14361 = n14276 | n14360;
  assign n9828 = ~n14359 & n14361;
  assign n9829 = x66 & x102;
  assign n9830 = n9828 & n9829;
  assign n9831 = n9828 | n9829;
  assign n9832 = ~n9830 & n9831;
  assign n14362 = n9645 & n9832;
  assign n14363 = (n9832 & n14281) | (n9832 & n14362) | (n14281 & n14362);
  assign n14364 = n9645 | n9832;
  assign n14365 = n14281 | n14364;
  assign n9835 = ~n14363 & n14365;
  assign n9836 = x65 & x103;
  assign n9837 = n9835 & n9836;
  assign n9838 = n9835 | n9836;
  assign n9839 = ~n9837 & n9838;
  assign n14299 = n9652 | n9654;
  assign n14366 = n9839 & n14299;
  assign n14367 = n9652 & n9839;
  assign n14368 = (n14202 & n14366) | (n14202 & n14367) | (n14366 & n14367);
  assign n14369 = n9839 | n14299;
  assign n14370 = n9652 | n9839;
  assign n14371 = (n14202 & n14369) | (n14202 & n14370) | (n14369 & n14370);
  assign n9842 = ~n14368 & n14371;
  assign n9843 = x64 & x104;
  assign n9844 = n9842 & n9843;
  assign n9845 = n9842 | n9843;
  assign n9846 = ~n9844 & n9845;
  assign n14297 = n9659 | n9661;
  assign n17084 = n9846 & n14297;
  assign n17085 = n9659 & n9846;
  assign n17086 = (n14200 & n17084) | (n14200 & n17085) | (n17084 & n17085);
  assign n17087 = n9846 | n14297;
  assign n17088 = n9659 | n9846;
  assign n17089 = (n14200 & n17087) | (n14200 & n17088) | (n17087 & n17088);
  assign n9849 = ~n17086 & n17089;
  assign n9850 = x63 & x105;
  assign n9851 = n9849 & n9850;
  assign n9852 = n9849 | n9850;
  assign n9853 = ~n9851 & n9852;
  assign n14295 = n9666 | n9668;
  assign n17090 = n9853 & n14295;
  assign n17091 = n9666 & n9853;
  assign n17092 = (n14198 & n17090) | (n14198 & n17091) | (n17090 & n17091);
  assign n17093 = n9853 | n14295;
  assign n17094 = n9666 | n9853;
  assign n17095 = (n14198 & n17093) | (n14198 & n17094) | (n17093 & n17094);
  assign n9856 = ~n17092 & n17095;
  assign n9857 = x62 & x106;
  assign n9858 = n9856 & n9857;
  assign n9859 = n9856 | n9857;
  assign n9860 = ~n9858 & n9859;
  assign n9861 = n14294 & n9860;
  assign n9862 = n14294 | n9860;
  assign n9863 = ~n9861 & n9862;
  assign n9864 = x61 & x107;
  assign n9865 = n9863 & n9864;
  assign n9866 = n9863 | n9864;
  assign n9867 = ~n9865 & n9866;
  assign n9868 = n14292 & n9867;
  assign n9869 = n14292 | n9867;
  assign n9870 = ~n9868 & n9869;
  assign n9871 = x60 & x108;
  assign n9872 = n9870 & n9871;
  assign n9873 = n9870 | n9871;
  assign n9874 = ~n9872 & n9873;
  assign n9875 = n14290 & n9874;
  assign n9876 = n14290 | n9874;
  assign n9877 = ~n9875 & n9876;
  assign n9878 = x59 & x109;
  assign n9879 = n9877 & n9878;
  assign n9880 = n9877 | n9878;
  assign n9881 = ~n9879 & n9880;
  assign n9882 = n14288 & n9881;
  assign n9883 = n14288 | n9881;
  assign n9884 = ~n9882 & n9883;
  assign n9885 = x58 & x110;
  assign n9886 = n9884 & n9885;
  assign n9887 = n9884 | n9885;
  assign n9888 = ~n9886 & n9887;
  assign n9889 = n14286 & n9888;
  assign n9890 = n14286 | n9888;
  assign n9891 = ~n9889 & n9890;
  assign n9892 = x57 & x111;
  assign n9893 = n9891 & n9892;
  assign n9894 = n9891 | n9892;
  assign n9895 = ~n9893 & n9894;
  assign n9896 = n9714 & n9895;
  assign n9897 = n9714 | n9895;
  assign n9898 = ~n9896 & n9897;
  assign n14372 = n9893 | n9895;
  assign n14373 = (n9714 & n9893) | (n9714 & n14372) | (n9893 & n14372);
  assign n14374 = n9886 | n9888;
  assign n14375 = (n9886 & n14286) | (n9886 & n14374) | (n14286 & n14374);
  assign n14376 = n9879 | n9881;
  assign n14377 = (n9879 & n14288) | (n9879 & n14376) | (n14288 & n14376);
  assign n14378 = n9872 | n9874;
  assign n14379 = (n9872 & n14290) | (n9872 & n14378) | (n14290 & n14378);
  assign n14380 = n9865 | n9867;
  assign n14381 = (n9865 & n14292) | (n9865 & n14380) | (n14292 & n14380);
  assign n14296 = (n9666 & n14198) | (n9666 & n14295) | (n14198 & n14295);
  assign n14298 = (n9659 & n14200) | (n9659 & n14297) | (n14200 & n14297);
  assign n14303 = (n16976 & n17037) | (n16976 & n14302) | (n17037 & n14302);
  assign n14391 = n9774 | n9776;
  assign n17096 = n9589 | n9774;
  assign n17097 = (n9774 & n9776) | (n9774 & n17096) | (n9776 & n17096);
  assign n17098 = (n14246 & n14391) | (n14246 & n17097) | (n14391 & n17097);
  assign n17099 = (n14245 & n14391) | (n14245 & n17097) | (n14391 & n17097);
  assign n17100 = (n14117 & n17098) | (n14117 & n17099) | (n17098 & n17099);
  assign n14396 = n9753 | n9755;
  assign n17101 = n9568 | n9753;
  assign n17102 = (n9753 & n9755) | (n9753 & n17101) | (n9755 & n17101);
  assign n17103 = (n14236 & n14396) | (n14236 & n17102) | (n14396 & n17102);
  assign n17104 = (n14235 & n14396) | (n14235 & n17102) | (n14396 & n17102);
  assign n17105 = (n16944 & n17103) | (n16944 & n17104) | (n17103 & n17104);
  assign n9922 = x79 & x90;
  assign n17106 = n9922 & n17053;
  assign n17107 = (n9741 & n9922) | (n9741 & n17106) | (n9922 & n17106);
  assign n14401 = n9922 & n17053;
  assign n14402 = (n17047 & n17107) | (n17047 & n14401) | (n17107 & n14401);
  assign n17108 = n9922 | n17053;
  assign n17109 = n9741 | n17108;
  assign n14404 = n9922 | n17053;
  assign n14405 = (n17047 & n17109) | (n17047 & n14404) | (n17109 & n14404);
  assign n9925 = ~n14402 & n14405;
  assign n14406 = n9746 & n9925;
  assign n17110 = (n9925 & n14319) | (n9925 & n14406) | (n14319 & n14406);
  assign n17111 = (n9925 & n14318) | (n9925 & n14406) | (n14318 & n14406);
  assign n17112 = (n17001 & n17110) | (n17001 & n17111) | (n17110 & n17111);
  assign n14408 = n9746 | n9925;
  assign n17113 = n14319 | n14408;
  assign n17114 = n14318 | n14408;
  assign n17115 = (n17001 & n17113) | (n17001 & n17114) | (n17113 & n17114);
  assign n9928 = ~n17112 & n17115;
  assign n9929 = x78 & x91;
  assign n9930 = n9928 & n9929;
  assign n9931 = n9928 | n9929;
  assign n9932 = ~n9930 & n9931;
  assign n9933 = n17105 & n9932;
  assign n9934 = n17105 | n9932;
  assign n9935 = ~n9933 & n9934;
  assign n9936 = x77 & x92;
  assign n9937 = n9935 & n9936;
  assign n9938 = n9935 | n9936;
  assign n9939 = ~n9937 & n9938;
  assign n14393 = n9760 | n9762;
  assign n14410 = n9939 & n14393;
  assign n14411 = n9760 & n9939;
  assign n14412 = (n17042 & n14410) | (n17042 & n14411) | (n14410 & n14411);
  assign n14413 = n9939 | n14393;
  assign n14414 = n9760 | n9939;
  assign n14415 = (n17042 & n14413) | (n17042 & n14414) | (n14413 & n14414);
  assign n9942 = ~n14412 & n14415;
  assign n9943 = x76 & x93;
  assign n9944 = n9942 & n9943;
  assign n9945 = n9942 | n9943;
  assign n9946 = ~n9944 & n9945;
  assign n14416 = n9767 & n9946;
  assign n17116 = (n9946 & n14329) | (n9946 & n14416) | (n14329 & n14416);
  assign n17117 = (n9946 & n14328) | (n9946 & n14416) | (n14328 & n14416);
  assign n17118 = (n16996 & n17116) | (n16996 & n17117) | (n17116 & n17117);
  assign n14418 = n9767 | n9946;
  assign n17119 = n14329 | n14418;
  assign n17120 = n14328 | n14418;
  assign n17121 = (n16996 & n17119) | (n16996 & n17120) | (n17119 & n17120);
  assign n9949 = ~n17118 & n17121;
  assign n9950 = x75 & x94;
  assign n9951 = n9949 & n9950;
  assign n9952 = n9949 | n9950;
  assign n9953 = ~n9951 & n9952;
  assign n9954 = n17100 & n9953;
  assign n9955 = n17100 | n9953;
  assign n9956 = ~n9954 & n9955;
  assign n9957 = x74 & x95;
  assign n9958 = n9956 & n9957;
  assign n9959 = n9956 | n9957;
  assign n9960 = ~n9958 & n9959;
  assign n14388 = n9781 | n9783;
  assign n14420 = n9960 & n14388;
  assign n14421 = n9781 & n9960;
  assign n14422 = (n14303 & n14420) | (n14303 & n14421) | (n14420 & n14421);
  assign n14423 = n9960 | n14388;
  assign n14424 = n9781 | n9960;
  assign n14425 = (n14303 & n14423) | (n14303 & n14424) | (n14423 & n14424);
  assign n9963 = ~n14422 & n14425;
  assign n9964 = x73 & x96;
  assign n9965 = n9963 & n9964;
  assign n9966 = n9963 | n9964;
  assign n9967 = ~n9965 & n9966;
  assign n14426 = n9788 & n9967;
  assign n14427 = (n9967 & n17080) | (n9967 & n14426) | (n17080 & n14426);
  assign n14428 = n9788 | n9967;
  assign n14429 = n17080 | n14428;
  assign n9970 = ~n14427 & n14429;
  assign n9971 = x72 & x97;
  assign n9972 = n9970 & n9971;
  assign n9973 = n9970 | n9971;
  assign n9974 = ~n9972 & n9973;
  assign n14430 = n9795 & n9974;
  assign n14431 = (n9974 & n14343) | (n9974 & n14430) | (n14343 & n14430);
  assign n14432 = n9795 | n9974;
  assign n14433 = n14343 | n14432;
  assign n9977 = ~n14431 & n14433;
  assign n9978 = x71 & x98;
  assign n9979 = n9977 & n9978;
  assign n9980 = n9977 | n9978;
  assign n9981 = ~n9979 & n9980;
  assign n14434 = n9802 & n9981;
  assign n14435 = (n9981 & n14347) | (n9981 & n14434) | (n14347 & n14434);
  assign n14436 = n9802 | n9981;
  assign n14437 = n14347 | n14436;
  assign n9984 = ~n14435 & n14437;
  assign n9985 = x70 & x99;
  assign n9986 = n9984 & n9985;
  assign n9987 = n9984 | n9985;
  assign n9988 = ~n9986 & n9987;
  assign n14438 = n9809 & n9988;
  assign n14439 = (n9988 & n14351) | (n9988 & n14438) | (n14351 & n14438);
  assign n14440 = n9809 | n9988;
  assign n14441 = n14351 | n14440;
  assign n9991 = ~n14439 & n14441;
  assign n9992 = x69 & x100;
  assign n9993 = n9991 & n9992;
  assign n9994 = n9991 | n9992;
  assign n9995 = ~n9993 & n9994;
  assign n14442 = n9816 & n9995;
  assign n14443 = (n9995 & n14355) | (n9995 & n14442) | (n14355 & n14442);
  assign n14444 = n9816 | n9995;
  assign n14445 = n14355 | n14444;
  assign n9998 = ~n14443 & n14445;
  assign n9999 = x68 & x101;
  assign n10000 = n9998 & n9999;
  assign n10001 = n9998 | n9999;
  assign n10002 = ~n10000 & n10001;
  assign n14446 = n9823 & n10002;
  assign n14447 = (n10002 & n14359) | (n10002 & n14446) | (n14359 & n14446);
  assign n14448 = n9823 | n10002;
  assign n14449 = n14359 | n14448;
  assign n10005 = ~n14447 & n14449;
  assign n10006 = x67 & x102;
  assign n10007 = n10005 & n10006;
  assign n10008 = n10005 | n10006;
  assign n10009 = ~n10007 & n10008;
  assign n14450 = n9830 & n10009;
  assign n14451 = (n10009 & n14363) | (n10009 & n14450) | (n14363 & n14450);
  assign n14452 = n9830 | n10009;
  assign n14453 = n14363 | n14452;
  assign n10012 = ~n14451 & n14453;
  assign n10013 = x66 & x103;
  assign n10014 = n10012 & n10013;
  assign n10015 = n10012 | n10013;
  assign n10016 = ~n10014 & n10015;
  assign n14454 = n9837 & n10016;
  assign n14455 = (n10016 & n14368) | (n10016 & n14454) | (n14368 & n14454);
  assign n14456 = n9837 | n10016;
  assign n14457 = n14368 | n14456;
  assign n10019 = ~n14455 & n14457;
  assign n10020 = x65 & x104;
  assign n10021 = n10019 & n10020;
  assign n10022 = n10019 | n10020;
  assign n10023 = ~n10021 & n10022;
  assign n14386 = n9844 | n9846;
  assign n14458 = n10023 & n14386;
  assign n14459 = n9844 & n10023;
  assign n14460 = (n14298 & n14458) | (n14298 & n14459) | (n14458 & n14459);
  assign n14461 = n10023 | n14386;
  assign n14462 = n9844 | n10023;
  assign n14463 = (n14298 & n14461) | (n14298 & n14462) | (n14461 & n14462);
  assign n10026 = ~n14460 & n14463;
  assign n10027 = x64 & x105;
  assign n10028 = n10026 & n10027;
  assign n10029 = n10026 | n10027;
  assign n10030 = ~n10028 & n10029;
  assign n14384 = n9851 | n9853;
  assign n17122 = n10030 & n14384;
  assign n17123 = n9851 & n10030;
  assign n17124 = (n14296 & n17122) | (n14296 & n17123) | (n17122 & n17123);
  assign n17125 = n10030 | n14384;
  assign n17126 = n9851 | n10030;
  assign n17127 = (n14296 & n17125) | (n14296 & n17126) | (n17125 & n17126);
  assign n10033 = ~n17124 & n17127;
  assign n10034 = x63 & x106;
  assign n10035 = n10033 & n10034;
  assign n10036 = n10033 | n10034;
  assign n10037 = ~n10035 & n10036;
  assign n14382 = n9858 | n9860;
  assign n17128 = n10037 & n14382;
  assign n17129 = n9858 & n10037;
  assign n17130 = (n14294 & n17128) | (n14294 & n17129) | (n17128 & n17129);
  assign n17131 = n10037 | n14382;
  assign n17132 = n9858 | n10037;
  assign n17133 = (n14294 & n17131) | (n14294 & n17132) | (n17131 & n17132);
  assign n10040 = ~n17130 & n17133;
  assign n10041 = x62 & x107;
  assign n10042 = n10040 & n10041;
  assign n10043 = n10040 | n10041;
  assign n10044 = ~n10042 & n10043;
  assign n10045 = n14381 & n10044;
  assign n10046 = n14381 | n10044;
  assign n10047 = ~n10045 & n10046;
  assign n10048 = x61 & x108;
  assign n10049 = n10047 & n10048;
  assign n10050 = n10047 | n10048;
  assign n10051 = ~n10049 & n10050;
  assign n10052 = n14379 & n10051;
  assign n10053 = n14379 | n10051;
  assign n10054 = ~n10052 & n10053;
  assign n10055 = x60 & x109;
  assign n10056 = n10054 & n10055;
  assign n10057 = n10054 | n10055;
  assign n10058 = ~n10056 & n10057;
  assign n10059 = n14377 & n10058;
  assign n10060 = n14377 | n10058;
  assign n10061 = ~n10059 & n10060;
  assign n10062 = x59 & x110;
  assign n10063 = n10061 & n10062;
  assign n10064 = n10061 | n10062;
  assign n10065 = ~n10063 & n10064;
  assign n10066 = n14375 & n10065;
  assign n10067 = n14375 | n10065;
  assign n10068 = ~n10066 & n10067;
  assign n10069 = x58 & x111;
  assign n10070 = n10068 & n10069;
  assign n10071 = n10068 | n10069;
  assign n10072 = ~n10070 & n10071;
  assign n10073 = n14373 & n10072;
  assign n10074 = n14373 | n10072;
  assign n10075 = ~n10073 & n10074;
  assign n14464 = n10070 | n10072;
  assign n14465 = (n10070 & n14373) | (n10070 & n14464) | (n14373 & n14464);
  assign n14466 = n10063 | n10065;
  assign n14467 = (n10063 & n14375) | (n10063 & n14466) | (n14375 & n14466);
  assign n14468 = n10056 | n10058;
  assign n14469 = (n10056 & n14377) | (n10056 & n14468) | (n14377 & n14468);
  assign n14470 = n10049 | n10051;
  assign n14471 = (n10049 & n14379) | (n10049 & n14470) | (n14379 & n14470);
  assign n14383 = (n9858 & n14294) | (n9858 & n14382) | (n14294 & n14382);
  assign n14385 = (n9851 & n14296) | (n9851 & n14384) | (n14296 & n14384);
  assign n14484 = n9944 | n9946;
  assign n17136 = n9767 | n9944;
  assign n17137 = (n9944 & n9946) | (n9944 & n17136) | (n9946 & n17136);
  assign n17138 = (n14329 & n14484) | (n14329 & n17137) | (n14484 & n17137);
  assign n17139 = (n14328 & n14484) | (n14328 & n17137) | (n14484 & n17137);
  assign n17140 = (n16996 & n17138) | (n16996 & n17139) | (n17138 & n17139);
  assign n10098 = x79 & x91;
  assign n14489 = n9925 | n14402;
  assign n17141 = (n9746 & n14402) | (n9746 & n14489) | (n14402 & n14489);
  assign n14491 = n10098 & n17141;
  assign n17844 = n10098 & n17107;
  assign n17845 = n10098 & n14401;
  assign n17846 = (n17047 & n17844) | (n17047 & n17845) | (n17844 & n17845);
  assign n17143 = (n9925 & n10098) | (n9925 & n17846) | (n10098 & n17846);
  assign n17144 = (n14319 & n14491) | (n14319 & n17143) | (n14491 & n17143);
  assign n17145 = (n14318 & n14491) | (n14318 & n17143) | (n14491 & n17143);
  assign n17146 = (n17001 & n17144) | (n17001 & n17145) | (n17144 & n17145);
  assign n14494 = n10098 | n17141;
  assign n17847 = n10098 | n17107;
  assign n17848 = n10098 | n14401;
  assign n17849 = (n17047 & n17847) | (n17047 & n17848) | (n17847 & n17848);
  assign n17148 = n9925 | n17849;
  assign n17149 = (n14319 & n14494) | (n14319 & n17148) | (n14494 & n17148);
  assign n17150 = (n14318 & n14494) | (n14318 & n17148) | (n14494 & n17148);
  assign n17151 = (n17001 & n17149) | (n17001 & n17150) | (n17149 & n17150);
  assign n10101 = ~n17146 & n17151;
  assign n14498 = n9930 & n10101;
  assign n17152 = (n9932 & n10101) | (n9932 & n14498) | (n10101 & n14498);
  assign n14499 = (n17105 & n17152) | (n17105 & n14498) | (n17152 & n14498);
  assign n14501 = n9930 | n10101;
  assign n17153 = n9932 | n14501;
  assign n14502 = (n17105 & n17153) | (n17105 & n14501) | (n17153 & n14501);
  assign n10104 = ~n14499 & n14502;
  assign n10105 = x78 & x92;
  assign n10106 = n10104 & n10105;
  assign n10107 = n10104 | n10105;
  assign n10108 = ~n10106 & n10107;
  assign n14503 = n9937 & n10108;
  assign n17154 = (n10108 & n14411) | (n10108 & n14503) | (n14411 & n14503);
  assign n17155 = (n10108 & n14410) | (n10108 & n14503) | (n14410 & n14503);
  assign n17156 = (n17042 & n17154) | (n17042 & n17155) | (n17154 & n17155);
  assign n14505 = n9937 | n10108;
  assign n17157 = n14411 | n14505;
  assign n17158 = n14410 | n14505;
  assign n17159 = (n17042 & n17157) | (n17042 & n17158) | (n17157 & n17158);
  assign n10111 = ~n17156 & n17159;
  assign n10112 = x77 & x93;
  assign n10113 = n10111 & n10112;
  assign n10114 = n10111 | n10112;
  assign n10115 = ~n10113 & n10114;
  assign n10116 = n17140 & n10115;
  assign n10117 = n17140 | n10115;
  assign n10118 = ~n10116 & n10117;
  assign n10119 = x76 & x94;
  assign n10120 = n10118 & n10119;
  assign n10121 = n10118 | n10119;
  assign n10122 = ~n10120 & n10121;
  assign n14481 = n9951 | n9953;
  assign n14507 = n10122 & n14481;
  assign n14508 = n9951 & n10122;
  assign n14509 = (n17100 & n14507) | (n17100 & n14508) | (n14507 & n14508);
  assign n14510 = n10122 | n14481;
  assign n14511 = n9951 | n10122;
  assign n14512 = (n17100 & n14510) | (n17100 & n14511) | (n14510 & n14511);
  assign n10125 = ~n14509 & n14512;
  assign n10126 = x75 & x95;
  assign n10127 = n10125 & n10126;
  assign n10128 = n10125 | n10126;
  assign n10129 = ~n10127 & n10128;
  assign n14513 = n9958 & n10129;
  assign n17160 = (n10129 & n14421) | (n10129 & n14513) | (n14421 & n14513);
  assign n17161 = (n10129 & n14420) | (n10129 & n14513) | (n14420 & n14513);
  assign n17162 = (n14303 & n17160) | (n14303 & n17161) | (n17160 & n17161);
  assign n14515 = n9958 | n10129;
  assign n17163 = n14421 | n14515;
  assign n17164 = n14420 | n14515;
  assign n17165 = (n14303 & n17163) | (n14303 & n17164) | (n17163 & n17164);
  assign n10132 = ~n17162 & n17165;
  assign n10133 = x74 & x96;
  assign n10134 = n10132 & n10133;
  assign n10135 = n10132 | n10133;
  assign n10136 = ~n10134 & n10135;
  assign n14479 = n9965 | n9967;
  assign n17166 = n10136 & n14479;
  assign n17134 = n9788 | n9965;
  assign n17135 = (n9965 & n9967) | (n9965 & n17134) | (n9967 & n17134);
  assign n17167 = n10136 & n17135;
  assign n17168 = (n17080 & n17166) | (n17080 & n17167) | (n17166 & n17167);
  assign n17169 = n10136 | n14479;
  assign n17170 = n10136 | n17135;
  assign n17171 = (n17080 & n17169) | (n17080 & n17170) | (n17169 & n17170);
  assign n10139 = ~n17168 & n17171;
  assign n10140 = x73 & x97;
  assign n10141 = n10139 & n10140;
  assign n10142 = n10139 | n10140;
  assign n10143 = ~n10141 & n10142;
  assign n14517 = n9972 & n10143;
  assign n17172 = (n10143 & n14430) | (n10143 & n14517) | (n14430 & n14517);
  assign n17173 = (n9974 & n10143) | (n9974 & n14517) | (n10143 & n14517);
  assign n17174 = (n14343 & n17172) | (n14343 & n17173) | (n17172 & n17173);
  assign n14519 = n9972 | n10143;
  assign n17175 = n14430 | n14519;
  assign n17176 = n9974 | n14519;
  assign n17177 = (n14343 & n17175) | (n14343 & n17176) | (n17175 & n17176);
  assign n10146 = ~n17174 & n17177;
  assign n10147 = x72 & x98;
  assign n10148 = n10146 & n10147;
  assign n10149 = n10146 | n10147;
  assign n10150 = ~n10148 & n10149;
  assign n14521 = n9979 & n10150;
  assign n14522 = (n10150 & n14435) | (n10150 & n14521) | (n14435 & n14521);
  assign n14523 = n9979 | n10150;
  assign n14524 = n14435 | n14523;
  assign n10153 = ~n14522 & n14524;
  assign n10154 = x71 & x99;
  assign n10155 = n10153 & n10154;
  assign n10156 = n10153 | n10154;
  assign n10157 = ~n10155 & n10156;
  assign n14525 = n9986 & n10157;
  assign n14526 = (n10157 & n14439) | (n10157 & n14525) | (n14439 & n14525);
  assign n14527 = n9986 | n10157;
  assign n14528 = n14439 | n14527;
  assign n10160 = ~n14526 & n14528;
  assign n10161 = x70 & x100;
  assign n10162 = n10160 & n10161;
  assign n10163 = n10160 | n10161;
  assign n10164 = ~n10162 & n10163;
  assign n14529 = n9993 & n10164;
  assign n14530 = (n10164 & n14443) | (n10164 & n14529) | (n14443 & n14529);
  assign n14531 = n9993 | n10164;
  assign n14532 = n14443 | n14531;
  assign n10167 = ~n14530 & n14532;
  assign n10168 = x69 & x101;
  assign n10169 = n10167 & n10168;
  assign n10170 = n10167 | n10168;
  assign n10171 = ~n10169 & n10170;
  assign n14533 = n10000 & n10171;
  assign n14534 = (n10171 & n14447) | (n10171 & n14533) | (n14447 & n14533);
  assign n14535 = n10000 | n10171;
  assign n14536 = n14447 | n14535;
  assign n10174 = ~n14534 & n14536;
  assign n10175 = x68 & x102;
  assign n10176 = n10174 & n10175;
  assign n10177 = n10174 | n10175;
  assign n10178 = ~n10176 & n10177;
  assign n14537 = n10007 & n10178;
  assign n14538 = (n10178 & n14451) | (n10178 & n14537) | (n14451 & n14537);
  assign n14539 = n10007 | n10178;
  assign n14540 = n14451 | n14539;
  assign n10181 = ~n14538 & n14540;
  assign n10182 = x67 & x103;
  assign n10183 = n10181 & n10182;
  assign n10184 = n10181 | n10182;
  assign n10185 = ~n10183 & n10184;
  assign n14541 = n10014 & n10185;
  assign n14542 = (n10185 & n14455) | (n10185 & n14541) | (n14455 & n14541);
  assign n14543 = n10014 | n10185;
  assign n14544 = n14455 | n14543;
  assign n10188 = ~n14542 & n14544;
  assign n10189 = x66 & x104;
  assign n10190 = n10188 & n10189;
  assign n10191 = n10188 | n10189;
  assign n10192 = ~n10190 & n10191;
  assign n14545 = n10021 & n10192;
  assign n14546 = (n10192 & n14460) | (n10192 & n14545) | (n14460 & n14545);
  assign n14547 = n10021 | n10192;
  assign n14548 = n14460 | n14547;
  assign n10195 = ~n14546 & n14548;
  assign n10196 = x65 & x105;
  assign n10197 = n10195 & n10196;
  assign n10198 = n10195 | n10196;
  assign n10199 = ~n10197 & n10198;
  assign n14476 = n10028 | n10030;
  assign n14549 = n10199 & n14476;
  assign n14550 = n10028 & n10199;
  assign n14551 = (n14385 & n14549) | (n14385 & n14550) | (n14549 & n14550);
  assign n14552 = n10199 | n14476;
  assign n14553 = n10028 | n10199;
  assign n14554 = (n14385 & n14552) | (n14385 & n14553) | (n14552 & n14553);
  assign n10202 = ~n14551 & n14554;
  assign n10203 = x64 & x106;
  assign n10204 = n10202 & n10203;
  assign n10205 = n10202 | n10203;
  assign n10206 = ~n10204 & n10205;
  assign n14474 = n10035 | n10037;
  assign n17178 = n10206 & n14474;
  assign n17179 = n10035 & n10206;
  assign n17180 = (n14383 & n17178) | (n14383 & n17179) | (n17178 & n17179);
  assign n17181 = n10206 | n14474;
  assign n17182 = n10035 | n10206;
  assign n17183 = (n14383 & n17181) | (n14383 & n17182) | (n17181 & n17182);
  assign n10209 = ~n17180 & n17183;
  assign n10210 = x63 & x107;
  assign n10211 = n10209 & n10210;
  assign n10212 = n10209 | n10210;
  assign n10213 = ~n10211 & n10212;
  assign n14472 = n10042 | n10044;
  assign n17184 = n10213 & n14472;
  assign n17185 = n10042 & n10213;
  assign n17186 = (n14381 & n17184) | (n14381 & n17185) | (n17184 & n17185);
  assign n17187 = n10213 | n14472;
  assign n17188 = n10042 | n10213;
  assign n17189 = (n14381 & n17187) | (n14381 & n17188) | (n17187 & n17188);
  assign n10216 = ~n17186 & n17189;
  assign n10217 = x62 & x108;
  assign n10218 = n10216 & n10217;
  assign n10219 = n10216 | n10217;
  assign n10220 = ~n10218 & n10219;
  assign n10221 = n14471 & n10220;
  assign n10222 = n14471 | n10220;
  assign n10223 = ~n10221 & n10222;
  assign n10224 = x61 & x109;
  assign n10225 = n10223 & n10224;
  assign n10226 = n10223 | n10224;
  assign n10227 = ~n10225 & n10226;
  assign n10228 = n14469 & n10227;
  assign n10229 = n14469 | n10227;
  assign n10230 = ~n10228 & n10229;
  assign n10231 = x60 & x110;
  assign n10232 = n10230 & n10231;
  assign n10233 = n10230 | n10231;
  assign n10234 = ~n10232 & n10233;
  assign n10235 = n14467 & n10234;
  assign n10236 = n14467 | n10234;
  assign n10237 = ~n10235 & n10236;
  assign n10238 = x59 & x111;
  assign n10239 = n10237 & n10238;
  assign n10240 = n10237 | n10238;
  assign n10241 = ~n10239 & n10240;
  assign n10242 = n14465 & n10241;
  assign n10243 = n14465 | n10241;
  assign n10244 = ~n10242 & n10243;
  assign n14555 = n10239 | n10241;
  assign n14556 = (n10239 & n14465) | (n10239 & n14555) | (n14465 & n14555);
  assign n14557 = n10232 | n10234;
  assign n14558 = (n10232 & n14467) | (n10232 & n14557) | (n14467 & n14557);
  assign n14559 = n10225 | n10227;
  assign n14560 = (n10225 & n14469) | (n10225 & n14559) | (n14469 & n14559);
  assign n14473 = (n10042 & n14381) | (n10042 & n14472) | (n14381 & n14472);
  assign n14475 = (n10035 & n14383) | (n10035 & n14474) | (n14383 & n14474);
  assign n14480 = (n17080 & n17135) | (n17080 & n14479) | (n17135 & n14479);
  assign n14570 = n10127 | n10129;
  assign n17190 = n9958 | n10127;
  assign n17191 = (n10127 & n10129) | (n10127 & n17190) | (n10129 & n17190);
  assign n17192 = (n14421 & n14570) | (n14421 & n17191) | (n14570 & n17191);
  assign n17193 = (n14420 & n14570) | (n14420 & n17191) | (n14570 & n17191);
  assign n17194 = (n14303 & n17192) | (n14303 & n17193) | (n17192 & n17193);
  assign n14575 = n10106 | n10108;
  assign n17195 = n9937 | n10106;
  assign n17196 = (n10106 & n10108) | (n10106 & n17195) | (n10108 & n17195);
  assign n17197 = (n14411 & n14575) | (n14411 & n17196) | (n14575 & n17196);
  assign n17198 = (n14410 & n14575) | (n14410 & n17196) | (n14575 & n17196);
  assign n17199 = (n17042 & n17197) | (n17042 & n17198) | (n17197 & n17198);
  assign n10266 = x79 & x92;
  assign n14577 = n10266 & n17146;
  assign n17200 = (n10266 & n14577) | (n10266 & n17152) | (n14577 & n17152);
  assign n17850 = (n10101 & n10266) | (n10101 & n14577) | (n10266 & n14577);
  assign n17851 = n10266 & n14577;
  assign n17852 = (n9930 & n17850) | (n9930 & n17851) | (n17850 & n17851);
  assign n17202 = (n17105 & n17200) | (n17105 & n17852) | (n17200 & n17852);
  assign n14579 = n10266 | n17146;
  assign n17203 = n14579 | n17152;
  assign n17853 = n10101 | n14579;
  assign n17854 = (n9930 & n14579) | (n9930 & n17853) | (n14579 & n17853);
  assign n17205 = (n17105 & n17203) | (n17105 & n17854) | (n17203 & n17854);
  assign n10269 = ~n17202 & n17205;
  assign n10270 = n17199 & n10269;
  assign n10271 = n17199 | n10269;
  assign n10272 = ~n10270 & n10271;
  assign n10273 = x78 & x93;
  assign n10274 = n10272 & n10273;
  assign n10275 = n10272 | n10273;
  assign n10276 = ~n10274 & n10275;
  assign n14572 = n10113 | n10115;
  assign n14581 = n10276 & n14572;
  assign n14582 = n10113 & n10276;
  assign n14583 = (n17140 & n14581) | (n17140 & n14582) | (n14581 & n14582);
  assign n14584 = n10276 | n14572;
  assign n14585 = n10113 | n10276;
  assign n14586 = (n17140 & n14584) | (n17140 & n14585) | (n14584 & n14585);
  assign n10279 = ~n14583 & n14586;
  assign n10280 = x77 & x94;
  assign n10281 = n10279 & n10280;
  assign n10282 = n10279 | n10280;
  assign n10283 = ~n10281 & n10282;
  assign n14587 = n10120 & n10283;
  assign n17206 = (n10283 & n14508) | (n10283 & n14587) | (n14508 & n14587);
  assign n17207 = (n10283 & n14507) | (n10283 & n14587) | (n14507 & n14587);
  assign n17208 = (n17100 & n17206) | (n17100 & n17207) | (n17206 & n17207);
  assign n14589 = n10120 | n10283;
  assign n17209 = n14508 | n14589;
  assign n17210 = n14507 | n14589;
  assign n17211 = (n17100 & n17209) | (n17100 & n17210) | (n17209 & n17210);
  assign n10286 = ~n17208 & n17211;
  assign n10287 = x76 & x95;
  assign n10288 = n10286 & n10287;
  assign n10289 = n10286 | n10287;
  assign n10290 = ~n10288 & n10289;
  assign n10291 = n17194 & n10290;
  assign n10292 = n17194 | n10290;
  assign n10293 = ~n10291 & n10292;
  assign n10294 = x75 & x96;
  assign n10295 = n10293 & n10294;
  assign n10296 = n10293 | n10294;
  assign n10297 = ~n10295 & n10296;
  assign n14567 = n10134 | n10136;
  assign n14591 = n10297 & n14567;
  assign n14592 = n10134 & n10297;
  assign n14593 = (n14480 & n14591) | (n14480 & n14592) | (n14591 & n14592);
  assign n14594 = n10297 | n14567;
  assign n14595 = n10134 | n10297;
  assign n14596 = (n14480 & n14594) | (n14480 & n14595) | (n14594 & n14595);
  assign n10300 = ~n14593 & n14596;
  assign n10301 = x74 & x97;
  assign n10302 = n10300 & n10301;
  assign n10303 = n10300 | n10301;
  assign n10304 = ~n10302 & n10303;
  assign n14597 = n10141 & n10304;
  assign n14598 = (n10304 & n17174) | (n10304 & n14597) | (n17174 & n14597);
  assign n14599 = n10141 | n10304;
  assign n14600 = n17174 | n14599;
  assign n10307 = ~n14598 & n14600;
  assign n10308 = x73 & x98;
  assign n10309 = n10307 & n10308;
  assign n10310 = n10307 | n10308;
  assign n10311 = ~n10309 & n10310;
  assign n14601 = n10148 & n10311;
  assign n14602 = (n10311 & n14522) | (n10311 & n14601) | (n14522 & n14601);
  assign n14603 = n10148 | n10311;
  assign n14604 = n14522 | n14603;
  assign n10314 = ~n14602 & n14604;
  assign n10315 = x72 & x99;
  assign n10316 = n10314 & n10315;
  assign n10317 = n10314 | n10315;
  assign n10318 = ~n10316 & n10317;
  assign n14605 = n10155 & n10318;
  assign n14606 = (n10318 & n14526) | (n10318 & n14605) | (n14526 & n14605);
  assign n14607 = n10155 | n10318;
  assign n14608 = n14526 | n14607;
  assign n10321 = ~n14606 & n14608;
  assign n10322 = x71 & x100;
  assign n10323 = n10321 & n10322;
  assign n10324 = n10321 | n10322;
  assign n10325 = ~n10323 & n10324;
  assign n14609 = n10162 & n10325;
  assign n14610 = (n10325 & n14530) | (n10325 & n14609) | (n14530 & n14609);
  assign n14611 = n10162 | n10325;
  assign n14612 = n14530 | n14611;
  assign n10328 = ~n14610 & n14612;
  assign n10329 = x70 & x101;
  assign n10330 = n10328 & n10329;
  assign n10331 = n10328 | n10329;
  assign n10332 = ~n10330 & n10331;
  assign n14613 = n10169 & n10332;
  assign n14614 = (n10332 & n14534) | (n10332 & n14613) | (n14534 & n14613);
  assign n14615 = n10169 | n10332;
  assign n14616 = n14534 | n14615;
  assign n10335 = ~n14614 & n14616;
  assign n10336 = x69 & x102;
  assign n10337 = n10335 & n10336;
  assign n10338 = n10335 | n10336;
  assign n10339 = ~n10337 & n10338;
  assign n14617 = n10176 & n10339;
  assign n14618 = (n10339 & n14538) | (n10339 & n14617) | (n14538 & n14617);
  assign n14619 = n10176 | n10339;
  assign n14620 = n14538 | n14619;
  assign n10342 = ~n14618 & n14620;
  assign n10343 = x68 & x103;
  assign n10344 = n10342 & n10343;
  assign n10345 = n10342 | n10343;
  assign n10346 = ~n10344 & n10345;
  assign n14621 = n10183 & n10346;
  assign n14622 = (n10346 & n14542) | (n10346 & n14621) | (n14542 & n14621);
  assign n14623 = n10183 | n10346;
  assign n14624 = n14542 | n14623;
  assign n10349 = ~n14622 & n14624;
  assign n10350 = x67 & x104;
  assign n10351 = n10349 & n10350;
  assign n10352 = n10349 | n10350;
  assign n10353 = ~n10351 & n10352;
  assign n14625 = n10190 & n10353;
  assign n14626 = (n10353 & n14546) | (n10353 & n14625) | (n14546 & n14625);
  assign n14627 = n10190 | n10353;
  assign n14628 = n14546 | n14627;
  assign n10356 = ~n14626 & n14628;
  assign n10357 = x66 & x105;
  assign n10358 = n10356 & n10357;
  assign n10359 = n10356 | n10357;
  assign n10360 = ~n10358 & n10359;
  assign n14629 = n10197 & n10360;
  assign n14630 = (n10360 & n14551) | (n10360 & n14629) | (n14551 & n14629);
  assign n14631 = n10197 | n10360;
  assign n14632 = n14551 | n14631;
  assign n10363 = ~n14630 & n14632;
  assign n10364 = x65 & x106;
  assign n10365 = n10363 & n10364;
  assign n10366 = n10363 | n10364;
  assign n10367 = ~n10365 & n10366;
  assign n14565 = n10204 | n10206;
  assign n14633 = n10367 & n14565;
  assign n14634 = n10204 & n10367;
  assign n14635 = (n14475 & n14633) | (n14475 & n14634) | (n14633 & n14634);
  assign n14636 = n10367 | n14565;
  assign n14637 = n10204 | n10367;
  assign n14638 = (n14475 & n14636) | (n14475 & n14637) | (n14636 & n14637);
  assign n10370 = ~n14635 & n14638;
  assign n10371 = x64 & x107;
  assign n10372 = n10370 & n10371;
  assign n10373 = n10370 | n10371;
  assign n10374 = ~n10372 & n10373;
  assign n14563 = n10211 | n10213;
  assign n17212 = n10374 & n14563;
  assign n17213 = n10211 & n10374;
  assign n17214 = (n14473 & n17212) | (n14473 & n17213) | (n17212 & n17213);
  assign n17215 = n10374 | n14563;
  assign n17216 = n10211 | n10374;
  assign n17217 = (n14473 & n17215) | (n14473 & n17216) | (n17215 & n17216);
  assign n10377 = ~n17214 & n17217;
  assign n10378 = x63 & x108;
  assign n10379 = n10377 & n10378;
  assign n10380 = n10377 | n10378;
  assign n10381 = ~n10379 & n10380;
  assign n14561 = n10218 | n10220;
  assign n17218 = n10381 & n14561;
  assign n17219 = n10218 & n10381;
  assign n17220 = (n14471 & n17218) | (n14471 & n17219) | (n17218 & n17219);
  assign n17221 = n10381 | n14561;
  assign n17222 = n10218 | n10381;
  assign n17223 = (n14471 & n17221) | (n14471 & n17222) | (n17221 & n17222);
  assign n10384 = ~n17220 & n17223;
  assign n10385 = x62 & x109;
  assign n10386 = n10384 & n10385;
  assign n10387 = n10384 | n10385;
  assign n10388 = ~n10386 & n10387;
  assign n10389 = n14560 & n10388;
  assign n10390 = n14560 | n10388;
  assign n10391 = ~n10389 & n10390;
  assign n10392 = x61 & x110;
  assign n10393 = n10391 & n10392;
  assign n10394 = n10391 | n10392;
  assign n10395 = ~n10393 & n10394;
  assign n10396 = n14558 & n10395;
  assign n10397 = n14558 | n10395;
  assign n10398 = ~n10396 & n10397;
  assign n10399 = x60 & x111;
  assign n10400 = n10398 & n10399;
  assign n10401 = n10398 | n10399;
  assign n10402 = ~n10400 & n10401;
  assign n10403 = n14556 & n10402;
  assign n10404 = n14556 | n10402;
  assign n10405 = ~n10403 & n10404;
  assign n14639 = n10400 | n10402;
  assign n14640 = (n10400 & n14556) | (n10400 & n14639) | (n14556 & n14639);
  assign n14641 = n10393 | n10395;
  assign n14642 = (n10393 & n14558) | (n10393 & n14641) | (n14558 & n14641);
  assign n14562 = (n10218 & n14471) | (n10218 & n14561) | (n14471 & n14561);
  assign n14564 = (n10211 & n14473) | (n10211 & n14563) | (n14473 & n14563);
  assign n14655 = n10281 | n10283;
  assign n17226 = n10120 | n10281;
  assign n17227 = (n10281 & n10283) | (n10281 & n17226) | (n10283 & n17226);
  assign n17228 = (n14508 & n14655) | (n14508 & n17227) | (n14655 & n17227);
  assign n17229 = (n14507 & n14655) | (n14507 & n17227) | (n14655 & n17227);
  assign n17230 = (n17100 & n17228) | (n17100 & n17229) | (n17228 & n17229);
  assign n10426 = x79 & x93;
  assign n17857 = n10426 & n14577;
  assign n17858 = n10266 & n10426;
  assign n17859 = (n17152 & n17857) | (n17152 & n17858) | (n17857 & n17858);
  assign n17855 = n10426 & n17852;
  assign n17856 = (n17105 & n17859) | (n17105 & n17855) | (n17859 & n17855);
  assign n17232 = (n10269 & n10426) | (n10269 & n17856) | (n10426 & n17856);
  assign n17234 = n10426 & n17852;
  assign n17235 = (n17105 & n17859) | (n17105 & n17234) | (n17859 & n17234);
  assign n14661 = (n17199 & n17232) | (n17199 & n17235) | (n17232 & n17235);
  assign n17862 = n10426 | n14577;
  assign n17863 = n10266 | n10426;
  assign n17864 = (n17152 & n17862) | (n17152 & n17863) | (n17862 & n17863);
  assign n17860 = n10426 | n17852;
  assign n17861 = (n17105 & n17864) | (n17105 & n17860) | (n17864 & n17860);
  assign n17237 = n10269 | n17861;
  assign n17239 = n10426 | n17852;
  assign n17240 = (n17105 & n17864) | (n17105 & n17239) | (n17864 & n17239);
  assign n14664 = (n17199 & n17237) | (n17199 & n17240) | (n17237 & n17240);
  assign n10429 = ~n14661 & n14664;
  assign n14665 = n10274 & n10429;
  assign n17241 = (n10429 & n14582) | (n10429 & n14665) | (n14582 & n14665);
  assign n17242 = (n10429 & n14581) | (n10429 & n14665) | (n14581 & n14665);
  assign n17243 = (n17140 & n17241) | (n17140 & n17242) | (n17241 & n17242);
  assign n14667 = n10274 | n10429;
  assign n17244 = n14582 | n14667;
  assign n17245 = n14581 | n14667;
  assign n17246 = (n17140 & n17244) | (n17140 & n17245) | (n17244 & n17245);
  assign n10432 = ~n17243 & n17246;
  assign n10433 = x78 & x94;
  assign n10434 = n10432 & n10433;
  assign n10435 = n10432 | n10433;
  assign n10436 = ~n10434 & n10435;
  assign n10437 = n17230 & n10436;
  assign n10438 = n17230 | n10436;
  assign n10439 = ~n10437 & n10438;
  assign n10440 = x77 & x95;
  assign n10441 = n10439 & n10440;
  assign n10442 = n10439 | n10440;
  assign n10443 = ~n10441 & n10442;
  assign n14652 = n10288 | n10290;
  assign n14669 = n10443 & n14652;
  assign n14670 = n10288 & n10443;
  assign n14671 = (n17194 & n14669) | (n17194 & n14670) | (n14669 & n14670);
  assign n14672 = n10443 | n14652;
  assign n14673 = n10288 | n10443;
  assign n14674 = (n17194 & n14672) | (n17194 & n14673) | (n14672 & n14673);
  assign n10446 = ~n14671 & n14674;
  assign n10447 = x76 & x96;
  assign n10448 = n10446 & n10447;
  assign n10449 = n10446 | n10447;
  assign n10450 = ~n10448 & n10449;
  assign n14675 = n10295 & n10450;
  assign n17247 = (n10450 & n14592) | (n10450 & n14675) | (n14592 & n14675);
  assign n17248 = (n10450 & n14591) | (n10450 & n14675) | (n14591 & n14675);
  assign n17249 = (n14480 & n17247) | (n14480 & n17248) | (n17247 & n17248);
  assign n14677 = n10295 | n10450;
  assign n17250 = n14592 | n14677;
  assign n17251 = n14591 | n14677;
  assign n17252 = (n14480 & n17250) | (n14480 & n17251) | (n17250 & n17251);
  assign n10453 = ~n17249 & n17252;
  assign n10454 = x75 & x97;
  assign n10455 = n10453 & n10454;
  assign n10456 = n10453 | n10454;
  assign n10457 = ~n10455 & n10456;
  assign n14650 = n10302 | n10304;
  assign n17253 = n10457 & n14650;
  assign n17224 = n10141 | n10302;
  assign n17225 = (n10302 & n10304) | (n10302 & n17224) | (n10304 & n17224);
  assign n17254 = n10457 & n17225;
  assign n17255 = (n17174 & n17253) | (n17174 & n17254) | (n17253 & n17254);
  assign n17256 = n10457 | n14650;
  assign n17257 = n10457 | n17225;
  assign n17258 = (n17174 & n17256) | (n17174 & n17257) | (n17256 & n17257);
  assign n10460 = ~n17255 & n17258;
  assign n10461 = x74 & x98;
  assign n10462 = n10460 & n10461;
  assign n10463 = n10460 | n10461;
  assign n10464 = ~n10462 & n10463;
  assign n14679 = n10309 & n10464;
  assign n17259 = (n10464 & n14601) | (n10464 & n14679) | (n14601 & n14679);
  assign n17260 = (n10311 & n10464) | (n10311 & n14679) | (n10464 & n14679);
  assign n17261 = (n14522 & n17259) | (n14522 & n17260) | (n17259 & n17260);
  assign n14681 = n10309 | n10464;
  assign n17262 = n14601 | n14681;
  assign n17263 = n10311 | n14681;
  assign n17264 = (n14522 & n17262) | (n14522 & n17263) | (n17262 & n17263);
  assign n10467 = ~n17261 & n17264;
  assign n10468 = x73 & x99;
  assign n10469 = n10467 & n10468;
  assign n10470 = n10467 | n10468;
  assign n10471 = ~n10469 & n10470;
  assign n14683 = n10316 & n10471;
  assign n14684 = (n10471 & n14606) | (n10471 & n14683) | (n14606 & n14683);
  assign n14685 = n10316 | n10471;
  assign n14686 = n14606 | n14685;
  assign n10474 = ~n14684 & n14686;
  assign n10475 = x72 & x100;
  assign n10476 = n10474 & n10475;
  assign n10477 = n10474 | n10475;
  assign n10478 = ~n10476 & n10477;
  assign n14687 = n10323 & n10478;
  assign n14688 = (n10478 & n14610) | (n10478 & n14687) | (n14610 & n14687);
  assign n14689 = n10323 | n10478;
  assign n14690 = n14610 | n14689;
  assign n10481 = ~n14688 & n14690;
  assign n10482 = x71 & x101;
  assign n10483 = n10481 & n10482;
  assign n10484 = n10481 | n10482;
  assign n10485 = ~n10483 & n10484;
  assign n14691 = n10330 & n10485;
  assign n14692 = (n10485 & n14614) | (n10485 & n14691) | (n14614 & n14691);
  assign n14693 = n10330 | n10485;
  assign n14694 = n14614 | n14693;
  assign n10488 = ~n14692 & n14694;
  assign n10489 = x70 & x102;
  assign n10490 = n10488 & n10489;
  assign n10491 = n10488 | n10489;
  assign n10492 = ~n10490 & n10491;
  assign n14695 = n10337 & n10492;
  assign n14696 = (n10492 & n14618) | (n10492 & n14695) | (n14618 & n14695);
  assign n14697 = n10337 | n10492;
  assign n14698 = n14618 | n14697;
  assign n10495 = ~n14696 & n14698;
  assign n10496 = x69 & x103;
  assign n10497 = n10495 & n10496;
  assign n10498 = n10495 | n10496;
  assign n10499 = ~n10497 & n10498;
  assign n14699 = n10344 & n10499;
  assign n14700 = (n10499 & n14622) | (n10499 & n14699) | (n14622 & n14699);
  assign n14701 = n10344 | n10499;
  assign n14702 = n14622 | n14701;
  assign n10502 = ~n14700 & n14702;
  assign n10503 = x68 & x104;
  assign n10504 = n10502 & n10503;
  assign n10505 = n10502 | n10503;
  assign n10506 = ~n10504 & n10505;
  assign n14703 = n10351 & n10506;
  assign n14704 = (n10506 & n14626) | (n10506 & n14703) | (n14626 & n14703);
  assign n14705 = n10351 | n10506;
  assign n14706 = n14626 | n14705;
  assign n10509 = ~n14704 & n14706;
  assign n10510 = x67 & x105;
  assign n10511 = n10509 & n10510;
  assign n10512 = n10509 | n10510;
  assign n10513 = ~n10511 & n10512;
  assign n14707 = n10358 & n10513;
  assign n14708 = (n10513 & n14630) | (n10513 & n14707) | (n14630 & n14707);
  assign n14709 = n10358 | n10513;
  assign n14710 = n14630 | n14709;
  assign n10516 = ~n14708 & n14710;
  assign n10517 = x66 & x106;
  assign n10518 = n10516 & n10517;
  assign n10519 = n10516 | n10517;
  assign n10520 = ~n10518 & n10519;
  assign n14711 = n10365 & n10520;
  assign n14712 = (n10520 & n14635) | (n10520 & n14711) | (n14635 & n14711);
  assign n14713 = n10365 | n10520;
  assign n14714 = n14635 | n14713;
  assign n10523 = ~n14712 & n14714;
  assign n10524 = x65 & x107;
  assign n10525 = n10523 & n10524;
  assign n10526 = n10523 | n10524;
  assign n10527 = ~n10525 & n10526;
  assign n14647 = n10372 | n10374;
  assign n14715 = n10527 & n14647;
  assign n14716 = n10372 & n10527;
  assign n14717 = (n14564 & n14715) | (n14564 & n14716) | (n14715 & n14716);
  assign n14718 = n10527 | n14647;
  assign n14719 = n10372 | n10527;
  assign n14720 = (n14564 & n14718) | (n14564 & n14719) | (n14718 & n14719);
  assign n10530 = ~n14717 & n14720;
  assign n10531 = x64 & x108;
  assign n10532 = n10530 & n10531;
  assign n10533 = n10530 | n10531;
  assign n10534 = ~n10532 & n10533;
  assign n14645 = n10379 | n10381;
  assign n17265 = n10534 & n14645;
  assign n17266 = n10379 & n10534;
  assign n17267 = (n14562 & n17265) | (n14562 & n17266) | (n17265 & n17266);
  assign n17268 = n10534 | n14645;
  assign n17269 = n10379 | n10534;
  assign n17270 = (n14562 & n17268) | (n14562 & n17269) | (n17268 & n17269);
  assign n10537 = ~n17267 & n17270;
  assign n10538 = x63 & x109;
  assign n10539 = n10537 & n10538;
  assign n10540 = n10537 | n10538;
  assign n10541 = ~n10539 & n10540;
  assign n14643 = n10386 | n10388;
  assign n17271 = n10541 & n14643;
  assign n17272 = n10386 & n10541;
  assign n17273 = (n14560 & n17271) | (n14560 & n17272) | (n17271 & n17272);
  assign n17274 = n10541 | n14643;
  assign n17275 = n10386 | n10541;
  assign n17276 = (n14560 & n17274) | (n14560 & n17275) | (n17274 & n17275);
  assign n10544 = ~n17273 & n17276;
  assign n10545 = x62 & x110;
  assign n10546 = n10544 & n10545;
  assign n10547 = n10544 | n10545;
  assign n10548 = ~n10546 & n10547;
  assign n10549 = n14642 & n10548;
  assign n10550 = n14642 | n10548;
  assign n10551 = ~n10549 & n10550;
  assign n10552 = x61 & x111;
  assign n10553 = n10551 & n10552;
  assign n10554 = n10551 | n10552;
  assign n10555 = ~n10553 & n10554;
  assign n10556 = n14640 & n10555;
  assign n10557 = n14640 | n10555;
  assign n10558 = ~n10556 & n10557;
  assign n14721 = n10553 | n10555;
  assign n14722 = (n10553 & n14640) | (n10553 & n14721) | (n14640 & n14721);
  assign n14644 = (n10386 & n14560) | (n10386 & n14643) | (n14560 & n14643);
  assign n14646 = (n10379 & n14562) | (n10379 & n14645) | (n14562 & n14645);
  assign n14651 = (n17174 & n17225) | (n17174 & n14650) | (n17225 & n14650);
  assign n14732 = n10448 | n10450;
  assign n17277 = n10295 | n10448;
  assign n17278 = (n10448 & n10450) | (n10448 & n17277) | (n10450 & n17277);
  assign n17279 = (n14592 & n14732) | (n14592 & n17278) | (n14732 & n17278);
  assign n17280 = (n14591 & n14732) | (n14591 & n17278) | (n14732 & n17278);
  assign n17281 = (n14480 & n17279) | (n14480 & n17280) | (n17279 & n17280);
  assign n10578 = x79 & x94;
  assign n14737 = n10429 | n14661;
  assign n17282 = (n10274 & n14661) | (n10274 & n14737) | (n14661 & n14737);
  assign n14739 = n10578 & n17282;
  assign n17865 = n10578 & n17232;
  assign n17866 = n10578 & n17235;
  assign n17867 = (n17199 & n17865) | (n17199 & n17866) | (n17865 & n17866);
  assign n17284 = (n10429 & n10578) | (n10429 & n17867) | (n10578 & n17867);
  assign n17285 = (n14582 & n14739) | (n14582 & n17284) | (n14739 & n17284);
  assign n17286 = (n14581 & n14739) | (n14581 & n17284) | (n14739 & n17284);
  assign n17287 = (n17140 & n17285) | (n17140 & n17286) | (n17285 & n17286);
  assign n14742 = n10578 | n17282;
  assign n17868 = n10578 | n17232;
  assign n17869 = n10578 | n17235;
  assign n17870 = (n17199 & n17868) | (n17199 & n17869) | (n17868 & n17869);
  assign n17289 = n10429 | n17870;
  assign n17290 = (n14582 & n14742) | (n14582 & n17289) | (n14742 & n17289);
  assign n17291 = (n14581 & n14742) | (n14581 & n17289) | (n14742 & n17289);
  assign n17292 = (n17140 & n17290) | (n17140 & n17291) | (n17290 & n17291);
  assign n10581 = ~n17287 & n17292;
  assign n14746 = n10434 & n10581;
  assign n17293 = (n10436 & n10581) | (n10436 & n14746) | (n10581 & n14746);
  assign n14747 = (n17230 & n17293) | (n17230 & n14746) | (n17293 & n14746);
  assign n14749 = n10434 | n10581;
  assign n17294 = n10436 | n14749;
  assign n14750 = (n17230 & n17294) | (n17230 & n14749) | (n17294 & n14749);
  assign n10584 = ~n14747 & n14750;
  assign n10585 = x78 & x95;
  assign n10586 = n10584 & n10585;
  assign n10587 = n10584 | n10585;
  assign n10588 = ~n10586 & n10587;
  assign n14751 = n10441 & n10588;
  assign n17295 = (n10588 & n14670) | (n10588 & n14751) | (n14670 & n14751);
  assign n17296 = (n10588 & n14669) | (n10588 & n14751) | (n14669 & n14751);
  assign n17297 = (n17194 & n17295) | (n17194 & n17296) | (n17295 & n17296);
  assign n14753 = n10441 | n10588;
  assign n17298 = n14670 | n14753;
  assign n17299 = n14669 | n14753;
  assign n17300 = (n17194 & n17298) | (n17194 & n17299) | (n17298 & n17299);
  assign n10591 = ~n17297 & n17300;
  assign n10592 = x77 & x96;
  assign n10593 = n10591 & n10592;
  assign n10594 = n10591 | n10592;
  assign n10595 = ~n10593 & n10594;
  assign n10596 = n17281 & n10595;
  assign n10597 = n17281 | n10595;
  assign n10598 = ~n10596 & n10597;
  assign n10599 = x76 & x97;
  assign n10600 = n10598 & n10599;
  assign n10601 = n10598 | n10599;
  assign n10602 = ~n10600 & n10601;
  assign n14729 = n10455 | n10457;
  assign n14755 = n10602 & n14729;
  assign n14756 = n10455 & n10602;
  assign n14757 = (n14651 & n14755) | (n14651 & n14756) | (n14755 & n14756);
  assign n14758 = n10602 | n14729;
  assign n14759 = n10455 | n10602;
  assign n14760 = (n14651 & n14758) | (n14651 & n14759) | (n14758 & n14759);
  assign n10605 = ~n14757 & n14760;
  assign n10606 = x75 & x98;
  assign n10607 = n10605 & n10606;
  assign n10608 = n10605 | n10606;
  assign n10609 = ~n10607 & n10608;
  assign n14761 = n10462 & n10609;
  assign n14762 = (n10609 & n17261) | (n10609 & n14761) | (n17261 & n14761);
  assign n14763 = n10462 | n10609;
  assign n14764 = n17261 | n14763;
  assign n10612 = ~n14762 & n14764;
  assign n10613 = x74 & x99;
  assign n10614 = n10612 & n10613;
  assign n10615 = n10612 | n10613;
  assign n10616 = ~n10614 & n10615;
  assign n14765 = n10469 & n10616;
  assign n14766 = (n10616 & n14684) | (n10616 & n14765) | (n14684 & n14765);
  assign n14767 = n10469 | n10616;
  assign n14768 = n14684 | n14767;
  assign n10619 = ~n14766 & n14768;
  assign n10620 = x73 & x100;
  assign n10621 = n10619 & n10620;
  assign n10622 = n10619 | n10620;
  assign n10623 = ~n10621 & n10622;
  assign n14769 = n10476 & n10623;
  assign n14770 = (n10623 & n14688) | (n10623 & n14769) | (n14688 & n14769);
  assign n14771 = n10476 | n10623;
  assign n14772 = n14688 | n14771;
  assign n10626 = ~n14770 & n14772;
  assign n10627 = x72 & x101;
  assign n10628 = n10626 & n10627;
  assign n10629 = n10626 | n10627;
  assign n10630 = ~n10628 & n10629;
  assign n14773 = n10483 & n10630;
  assign n14774 = (n10630 & n14692) | (n10630 & n14773) | (n14692 & n14773);
  assign n14775 = n10483 | n10630;
  assign n14776 = n14692 | n14775;
  assign n10633 = ~n14774 & n14776;
  assign n10634 = x71 & x102;
  assign n10635 = n10633 & n10634;
  assign n10636 = n10633 | n10634;
  assign n10637 = ~n10635 & n10636;
  assign n14777 = n10490 & n10637;
  assign n14778 = (n10637 & n14696) | (n10637 & n14777) | (n14696 & n14777);
  assign n14779 = n10490 | n10637;
  assign n14780 = n14696 | n14779;
  assign n10640 = ~n14778 & n14780;
  assign n10641 = x70 & x103;
  assign n10642 = n10640 & n10641;
  assign n10643 = n10640 | n10641;
  assign n10644 = ~n10642 & n10643;
  assign n14781 = n10497 & n10644;
  assign n14782 = (n10644 & n14700) | (n10644 & n14781) | (n14700 & n14781);
  assign n14783 = n10497 | n10644;
  assign n14784 = n14700 | n14783;
  assign n10647 = ~n14782 & n14784;
  assign n10648 = x69 & x104;
  assign n10649 = n10647 & n10648;
  assign n10650 = n10647 | n10648;
  assign n10651 = ~n10649 & n10650;
  assign n14785 = n10504 & n10651;
  assign n14786 = (n10651 & n14704) | (n10651 & n14785) | (n14704 & n14785);
  assign n14787 = n10504 | n10651;
  assign n14788 = n14704 | n14787;
  assign n10654 = ~n14786 & n14788;
  assign n10655 = x68 & x105;
  assign n10656 = n10654 & n10655;
  assign n10657 = n10654 | n10655;
  assign n10658 = ~n10656 & n10657;
  assign n14789 = n10511 & n10658;
  assign n14790 = (n10658 & n14708) | (n10658 & n14789) | (n14708 & n14789);
  assign n14791 = n10511 | n10658;
  assign n14792 = n14708 | n14791;
  assign n10661 = ~n14790 & n14792;
  assign n10662 = x67 & x106;
  assign n10663 = n10661 & n10662;
  assign n10664 = n10661 | n10662;
  assign n10665 = ~n10663 & n10664;
  assign n14793 = n10518 & n10665;
  assign n14794 = (n10665 & n14712) | (n10665 & n14793) | (n14712 & n14793);
  assign n14795 = n10518 | n10665;
  assign n14796 = n14712 | n14795;
  assign n10668 = ~n14794 & n14796;
  assign n10669 = x66 & x107;
  assign n10670 = n10668 & n10669;
  assign n10671 = n10668 | n10669;
  assign n10672 = ~n10670 & n10671;
  assign n14797 = n10525 & n10672;
  assign n14798 = (n10672 & n14717) | (n10672 & n14797) | (n14717 & n14797);
  assign n14799 = n10525 | n10672;
  assign n14800 = n14717 | n14799;
  assign n10675 = ~n14798 & n14800;
  assign n10676 = x65 & x108;
  assign n10677 = n10675 & n10676;
  assign n10678 = n10675 | n10676;
  assign n10679 = ~n10677 & n10678;
  assign n14727 = n10532 | n10534;
  assign n14801 = n10679 & n14727;
  assign n14802 = n10532 & n10679;
  assign n14803 = (n14646 & n14801) | (n14646 & n14802) | (n14801 & n14802);
  assign n14804 = n10679 | n14727;
  assign n14805 = n10532 | n10679;
  assign n14806 = (n14646 & n14804) | (n14646 & n14805) | (n14804 & n14805);
  assign n10682 = ~n14803 & n14806;
  assign n10683 = x64 & x109;
  assign n10684 = n10682 & n10683;
  assign n10685 = n10682 | n10683;
  assign n10686 = ~n10684 & n10685;
  assign n14725 = n10539 | n10541;
  assign n17301 = n10686 & n14725;
  assign n17302 = n10539 & n10686;
  assign n17303 = (n14644 & n17301) | (n14644 & n17302) | (n17301 & n17302);
  assign n17304 = n10686 | n14725;
  assign n17305 = n10539 | n10686;
  assign n17306 = (n14644 & n17304) | (n14644 & n17305) | (n17304 & n17305);
  assign n10689 = ~n17303 & n17306;
  assign n10690 = x63 & x110;
  assign n10691 = n10689 & n10690;
  assign n10692 = n10689 | n10690;
  assign n10693 = ~n10691 & n10692;
  assign n14723 = n10546 | n10548;
  assign n17307 = n10693 & n14723;
  assign n17308 = n10546 & n10693;
  assign n17309 = (n14642 & n17307) | (n14642 & n17308) | (n17307 & n17308);
  assign n17310 = n10693 | n14723;
  assign n17311 = n10546 | n10693;
  assign n17312 = (n14642 & n17310) | (n14642 & n17311) | (n17310 & n17311);
  assign n10696 = ~n17309 & n17312;
  assign n10697 = x62 & x111;
  assign n10698 = n10696 & n10697;
  assign n10699 = n10696 | n10697;
  assign n10700 = ~n10698 & n10699;
  assign n10701 = n14722 & n10700;
  assign n10702 = n14722 | n10700;
  assign n10703 = ~n10701 & n10702;
  assign n14724 = (n10546 & n14642) | (n10546 & n14723) | (n14642 & n14723);
  assign n14726 = (n10539 & n14644) | (n10539 & n14725) | (n14644 & n14725);
  assign n14819 = n10586 | n10588;
  assign n17315 = n10441 | n10586;
  assign n17316 = (n10586 & n10588) | (n10586 & n17315) | (n10588 & n17315);
  assign n17317 = (n14670 & n14819) | (n14670 & n17316) | (n14819 & n17316);
  assign n17318 = (n14669 & n14819) | (n14669 & n17316) | (n14819 & n17316);
  assign n17319 = (n17194 & n17317) | (n17194 & n17318) | (n17317 & n17318);
  assign n10722 = x79 & x95;
  assign n14821 = n10722 & n17287;
  assign n17320 = (n10722 & n14821) | (n10722 & n17293) | (n14821 & n17293);
  assign n17871 = (n10581 & n10722) | (n10581 & n14821) | (n10722 & n14821);
  assign n17872 = n10722 & n14821;
  assign n17873 = (n10434 & n17871) | (n10434 & n17872) | (n17871 & n17872);
  assign n17322 = (n17230 & n17320) | (n17230 & n17873) | (n17320 & n17873);
  assign n14823 = n10722 | n17287;
  assign n17323 = n14823 | n17293;
  assign n17874 = n10581 | n14823;
  assign n17875 = (n10434 & n14823) | (n10434 & n17874) | (n14823 & n17874);
  assign n17325 = (n17230 & n17323) | (n17230 & n17875) | (n17323 & n17875);
  assign n10725 = ~n17322 & n17325;
  assign n10726 = n17319 & n10725;
  assign n10727 = n17319 | n10725;
  assign n10728 = ~n10726 & n10727;
  assign n10729 = x78 & x96;
  assign n10730 = n10728 & n10729;
  assign n10731 = n10728 | n10729;
  assign n10732 = ~n10730 & n10731;
  assign n14816 = n10593 | n10595;
  assign n14825 = n10732 & n14816;
  assign n14826 = n10593 & n10732;
  assign n14827 = (n17281 & n14825) | (n17281 & n14826) | (n14825 & n14826);
  assign n14828 = n10732 | n14816;
  assign n14829 = n10593 | n10732;
  assign n14830 = (n17281 & n14828) | (n17281 & n14829) | (n14828 & n14829);
  assign n10735 = ~n14827 & n14830;
  assign n10736 = x77 & x97;
  assign n10737 = n10735 & n10736;
  assign n10738 = n10735 | n10736;
  assign n10739 = ~n10737 & n10738;
  assign n14831 = n10600 & n10739;
  assign n17326 = (n10739 & n14756) | (n10739 & n14831) | (n14756 & n14831);
  assign n17327 = (n10739 & n14755) | (n10739 & n14831) | (n14755 & n14831);
  assign n17328 = (n14651 & n17326) | (n14651 & n17327) | (n17326 & n17327);
  assign n14833 = n10600 | n10739;
  assign n17329 = n14756 | n14833;
  assign n17330 = n14755 | n14833;
  assign n17331 = (n14651 & n17329) | (n14651 & n17330) | (n17329 & n17330);
  assign n10742 = ~n17328 & n17331;
  assign n10743 = x76 & x98;
  assign n10744 = n10742 & n10743;
  assign n10745 = n10742 | n10743;
  assign n10746 = ~n10744 & n10745;
  assign n14814 = n10607 | n10609;
  assign n17332 = n10746 & n14814;
  assign n17313 = n10462 | n10607;
  assign n17314 = (n10607 & n10609) | (n10607 & n17313) | (n10609 & n17313);
  assign n17333 = n10746 & n17314;
  assign n17334 = (n17261 & n17332) | (n17261 & n17333) | (n17332 & n17333);
  assign n17335 = n10746 | n14814;
  assign n17336 = n10746 | n17314;
  assign n17337 = (n17261 & n17335) | (n17261 & n17336) | (n17335 & n17336);
  assign n10749 = ~n17334 & n17337;
  assign n10750 = x75 & x99;
  assign n10751 = n10749 & n10750;
  assign n10752 = n10749 | n10750;
  assign n10753 = ~n10751 & n10752;
  assign n14835 = n10614 & n10753;
  assign n17338 = (n10753 & n14765) | (n10753 & n14835) | (n14765 & n14835);
  assign n17339 = (n10616 & n10753) | (n10616 & n14835) | (n10753 & n14835);
  assign n17340 = (n14684 & n17338) | (n14684 & n17339) | (n17338 & n17339);
  assign n14837 = n10614 | n10753;
  assign n17341 = n14765 | n14837;
  assign n17342 = n10616 | n14837;
  assign n17343 = (n14684 & n17341) | (n14684 & n17342) | (n17341 & n17342);
  assign n10756 = ~n17340 & n17343;
  assign n10757 = x74 & x100;
  assign n10758 = n10756 & n10757;
  assign n10759 = n10756 | n10757;
  assign n10760 = ~n10758 & n10759;
  assign n14839 = n10621 & n10760;
  assign n14840 = (n10760 & n14770) | (n10760 & n14839) | (n14770 & n14839);
  assign n14841 = n10621 | n10760;
  assign n14842 = n14770 | n14841;
  assign n10763 = ~n14840 & n14842;
  assign n10764 = x73 & x101;
  assign n10765 = n10763 & n10764;
  assign n10766 = n10763 | n10764;
  assign n10767 = ~n10765 & n10766;
  assign n14843 = n10628 & n10767;
  assign n14844 = (n10767 & n14774) | (n10767 & n14843) | (n14774 & n14843);
  assign n14845 = n10628 | n10767;
  assign n14846 = n14774 | n14845;
  assign n10770 = ~n14844 & n14846;
  assign n10771 = x72 & x102;
  assign n10772 = n10770 & n10771;
  assign n10773 = n10770 | n10771;
  assign n10774 = ~n10772 & n10773;
  assign n14847 = n10635 & n10774;
  assign n14848 = (n10774 & n14778) | (n10774 & n14847) | (n14778 & n14847);
  assign n14849 = n10635 | n10774;
  assign n14850 = n14778 | n14849;
  assign n10777 = ~n14848 & n14850;
  assign n10778 = x71 & x103;
  assign n10779 = n10777 & n10778;
  assign n10780 = n10777 | n10778;
  assign n10781 = ~n10779 & n10780;
  assign n14851 = n10642 & n10781;
  assign n14852 = (n10781 & n14782) | (n10781 & n14851) | (n14782 & n14851);
  assign n14853 = n10642 | n10781;
  assign n14854 = n14782 | n14853;
  assign n10784 = ~n14852 & n14854;
  assign n10785 = x70 & x104;
  assign n10786 = n10784 & n10785;
  assign n10787 = n10784 | n10785;
  assign n10788 = ~n10786 & n10787;
  assign n14855 = n10649 & n10788;
  assign n14856 = (n10788 & n14786) | (n10788 & n14855) | (n14786 & n14855);
  assign n14857 = n10649 | n10788;
  assign n14858 = n14786 | n14857;
  assign n10791 = ~n14856 & n14858;
  assign n10792 = x69 & x105;
  assign n10793 = n10791 & n10792;
  assign n10794 = n10791 | n10792;
  assign n10795 = ~n10793 & n10794;
  assign n14859 = n10656 & n10795;
  assign n14860 = (n10795 & n14790) | (n10795 & n14859) | (n14790 & n14859);
  assign n14861 = n10656 | n10795;
  assign n14862 = n14790 | n14861;
  assign n10798 = ~n14860 & n14862;
  assign n10799 = x68 & x106;
  assign n10800 = n10798 & n10799;
  assign n10801 = n10798 | n10799;
  assign n10802 = ~n10800 & n10801;
  assign n14863 = n10663 & n10802;
  assign n14864 = (n10802 & n14794) | (n10802 & n14863) | (n14794 & n14863);
  assign n14865 = n10663 | n10802;
  assign n14866 = n14794 | n14865;
  assign n10805 = ~n14864 & n14866;
  assign n10806 = x67 & x107;
  assign n10807 = n10805 & n10806;
  assign n10808 = n10805 | n10806;
  assign n10809 = ~n10807 & n10808;
  assign n14867 = n10670 & n10809;
  assign n14868 = (n10809 & n14798) | (n10809 & n14867) | (n14798 & n14867);
  assign n14869 = n10670 | n10809;
  assign n14870 = n14798 | n14869;
  assign n10812 = ~n14868 & n14870;
  assign n10813 = x66 & x108;
  assign n10814 = n10812 & n10813;
  assign n10815 = n10812 | n10813;
  assign n10816 = ~n10814 & n10815;
  assign n14871 = n10677 & n10816;
  assign n14872 = (n10816 & n14803) | (n10816 & n14871) | (n14803 & n14871);
  assign n14873 = n10677 | n10816;
  assign n14874 = n14803 | n14873;
  assign n10819 = ~n14872 & n14874;
  assign n10820 = x65 & x109;
  assign n10821 = n10819 & n10820;
  assign n10822 = n10819 | n10820;
  assign n10823 = ~n10821 & n10822;
  assign n14811 = n10684 | n10686;
  assign n14875 = n10823 & n14811;
  assign n14876 = n10684 & n10823;
  assign n14877 = (n14726 & n14875) | (n14726 & n14876) | (n14875 & n14876);
  assign n14878 = n10823 | n14811;
  assign n14879 = n10684 | n10823;
  assign n14880 = (n14726 & n14878) | (n14726 & n14879) | (n14878 & n14879);
  assign n10826 = ~n14877 & n14880;
  assign n10827 = x64 & x110;
  assign n10828 = n10826 & n10827;
  assign n10829 = n10826 | n10827;
  assign n10830 = ~n10828 & n10829;
  assign n14809 = n10691 | n10693;
  assign n17344 = n10830 & n14809;
  assign n17345 = n10691 & n10830;
  assign n17346 = (n14724 & n17344) | (n14724 & n17345) | (n17344 & n17345);
  assign n17347 = n10830 | n14809;
  assign n17348 = n10691 | n10830;
  assign n17349 = (n14724 & n17347) | (n14724 & n17348) | (n17347 & n17348);
  assign n10833 = ~n17346 & n17349;
  assign n10834 = x63 & x111;
  assign n10835 = n10833 & n10834;
  assign n10836 = n10833 | n10834;
  assign n10837 = ~n10835 & n10836;
  assign n14807 = n10698 | n10700;
  assign n17350 = n10837 & n14807;
  assign n17351 = n10698 & n10837;
  assign n17352 = (n14722 & n17350) | (n14722 & n17351) | (n17350 & n17351);
  assign n17353 = n10837 | n14807;
  assign n17354 = n10698 | n10837;
  assign n17355 = (n14722 & n17353) | (n14722 & n17354) | (n17353 & n17354);
  assign n10840 = ~n17352 & n17355;
  assign n14808 = (n10698 & n14722) | (n10698 & n14807) | (n14722 & n14807);
  assign n14810 = (n10691 & n14724) | (n10691 & n14809) | (n14724 & n14809);
  assign n14815 = (n17261 & n17314) | (n17261 & n14814) | (n17314 & n14814);
  assign n14888 = n10737 | n10739;
  assign n17356 = n10600 | n10737;
  assign n17357 = (n10737 & n10739) | (n10737 & n17356) | (n10739 & n17356);
  assign n17358 = (n14756 & n14888) | (n14756 & n17357) | (n14888 & n17357);
  assign n17359 = (n14755 & n14888) | (n14755 & n17357) | (n14888 & n17357);
  assign n17360 = (n14651 & n17358) | (n14651 & n17359) | (n17358 & n17359);
  assign n10858 = x79 & x96;
  assign n17878 = n10858 & n14821;
  assign n17879 = n10722 & n10858;
  assign n17880 = (n17293 & n17878) | (n17293 & n17879) | (n17878 & n17879);
  assign n17876 = n10858 & n17873;
  assign n17877 = (n17230 & n17880) | (n17230 & n17876) | (n17880 & n17876);
  assign n17362 = (n10725 & n10858) | (n10725 & n17877) | (n10858 & n17877);
  assign n17364 = n10858 & n17873;
  assign n17365 = (n17230 & n17880) | (n17230 & n17364) | (n17880 & n17364);
  assign n14894 = (n17319 & n17362) | (n17319 & n17365) | (n17362 & n17365);
  assign n17883 = n10858 | n14821;
  assign n17884 = n10722 | n10858;
  assign n17885 = (n17293 & n17883) | (n17293 & n17884) | (n17883 & n17884);
  assign n17881 = n10858 | n17873;
  assign n17882 = (n17230 & n17885) | (n17230 & n17881) | (n17885 & n17881);
  assign n17367 = n10725 | n17882;
  assign n17369 = n10858 | n17873;
  assign n17370 = (n17230 & n17885) | (n17230 & n17369) | (n17885 & n17369);
  assign n14897 = (n17319 & n17367) | (n17319 & n17370) | (n17367 & n17370);
  assign n10861 = ~n14894 & n14897;
  assign n14898 = n10730 & n10861;
  assign n17371 = (n10861 & n14826) | (n10861 & n14898) | (n14826 & n14898);
  assign n17372 = (n10861 & n14825) | (n10861 & n14898) | (n14825 & n14898);
  assign n17373 = (n17281 & n17371) | (n17281 & n17372) | (n17371 & n17372);
  assign n14900 = n10730 | n10861;
  assign n17374 = n14826 | n14900;
  assign n17375 = n14825 | n14900;
  assign n17376 = (n17281 & n17374) | (n17281 & n17375) | (n17374 & n17375);
  assign n10864 = ~n17373 & n17376;
  assign n10865 = x78 & x97;
  assign n10866 = n10864 & n10865;
  assign n10867 = n10864 | n10865;
  assign n10868 = ~n10866 & n10867;
  assign n10869 = n17360 & n10868;
  assign n10870 = n17360 | n10868;
  assign n10871 = ~n10869 & n10870;
  assign n10872 = x77 & x98;
  assign n10873 = n10871 & n10872;
  assign n10874 = n10871 | n10872;
  assign n10875 = ~n10873 & n10874;
  assign n14885 = n10744 | n10746;
  assign n14902 = n10875 & n14885;
  assign n14903 = n10744 & n10875;
  assign n14904 = (n14815 & n14902) | (n14815 & n14903) | (n14902 & n14903);
  assign n14905 = n10875 | n14885;
  assign n14906 = n10744 | n10875;
  assign n14907 = (n14815 & n14905) | (n14815 & n14906) | (n14905 & n14906);
  assign n10878 = ~n14904 & n14907;
  assign n10879 = x76 & x99;
  assign n10880 = n10878 & n10879;
  assign n10881 = n10878 | n10879;
  assign n10882 = ~n10880 & n10881;
  assign n14908 = n10751 & n10882;
  assign n14909 = (n10882 & n17340) | (n10882 & n14908) | (n17340 & n14908);
  assign n14910 = n10751 | n10882;
  assign n14911 = n17340 | n14910;
  assign n10885 = ~n14909 & n14911;
  assign n10886 = x75 & x100;
  assign n10887 = n10885 & n10886;
  assign n10888 = n10885 | n10886;
  assign n10889 = ~n10887 & n10888;
  assign n14912 = n10758 & n10889;
  assign n14913 = (n10889 & n14840) | (n10889 & n14912) | (n14840 & n14912);
  assign n14914 = n10758 | n10889;
  assign n14915 = n14840 | n14914;
  assign n10892 = ~n14913 & n14915;
  assign n10893 = x74 & x101;
  assign n10894 = n10892 & n10893;
  assign n10895 = n10892 | n10893;
  assign n10896 = ~n10894 & n10895;
  assign n14916 = n10765 & n10896;
  assign n14917 = (n10896 & n14844) | (n10896 & n14916) | (n14844 & n14916);
  assign n14918 = n10765 | n10896;
  assign n14919 = n14844 | n14918;
  assign n10899 = ~n14917 & n14919;
  assign n10900 = x73 & x102;
  assign n10901 = n10899 & n10900;
  assign n10902 = n10899 | n10900;
  assign n10903 = ~n10901 & n10902;
  assign n14920 = n10772 & n10903;
  assign n14921 = (n10903 & n14848) | (n10903 & n14920) | (n14848 & n14920);
  assign n14922 = n10772 | n10903;
  assign n14923 = n14848 | n14922;
  assign n10906 = ~n14921 & n14923;
  assign n10907 = x72 & x103;
  assign n10908 = n10906 & n10907;
  assign n10909 = n10906 | n10907;
  assign n10910 = ~n10908 & n10909;
  assign n14924 = n10779 & n10910;
  assign n14925 = (n10910 & n14852) | (n10910 & n14924) | (n14852 & n14924);
  assign n14926 = n10779 | n10910;
  assign n14927 = n14852 | n14926;
  assign n10913 = ~n14925 & n14927;
  assign n10914 = x71 & x104;
  assign n10915 = n10913 & n10914;
  assign n10916 = n10913 | n10914;
  assign n10917 = ~n10915 & n10916;
  assign n14928 = n10786 & n10917;
  assign n14929 = (n10917 & n14856) | (n10917 & n14928) | (n14856 & n14928);
  assign n14930 = n10786 | n10917;
  assign n14931 = n14856 | n14930;
  assign n10920 = ~n14929 & n14931;
  assign n10921 = x70 & x105;
  assign n10922 = n10920 & n10921;
  assign n10923 = n10920 | n10921;
  assign n10924 = ~n10922 & n10923;
  assign n14932 = n10793 & n10924;
  assign n14933 = (n10924 & n14860) | (n10924 & n14932) | (n14860 & n14932);
  assign n14934 = n10793 | n10924;
  assign n14935 = n14860 | n14934;
  assign n10927 = ~n14933 & n14935;
  assign n10928 = x69 & x106;
  assign n10929 = n10927 & n10928;
  assign n10930 = n10927 | n10928;
  assign n10931 = ~n10929 & n10930;
  assign n14936 = n10800 & n10931;
  assign n14937 = (n10931 & n14864) | (n10931 & n14936) | (n14864 & n14936);
  assign n14938 = n10800 | n10931;
  assign n14939 = n14864 | n14938;
  assign n10934 = ~n14937 & n14939;
  assign n10935 = x68 & x107;
  assign n10936 = n10934 & n10935;
  assign n10937 = n10934 | n10935;
  assign n10938 = ~n10936 & n10937;
  assign n14940 = n10807 & n10938;
  assign n14941 = (n10938 & n14868) | (n10938 & n14940) | (n14868 & n14940);
  assign n14942 = n10807 | n10938;
  assign n14943 = n14868 | n14942;
  assign n10941 = ~n14941 & n14943;
  assign n10942 = x67 & x108;
  assign n10943 = n10941 & n10942;
  assign n10944 = n10941 | n10942;
  assign n10945 = ~n10943 & n10944;
  assign n14944 = n10814 & n10945;
  assign n14945 = (n10945 & n14872) | (n10945 & n14944) | (n14872 & n14944);
  assign n14946 = n10814 | n10945;
  assign n14947 = n14872 | n14946;
  assign n10948 = ~n14945 & n14947;
  assign n10949 = x66 & x109;
  assign n10950 = n10948 & n10949;
  assign n10951 = n10948 | n10949;
  assign n10952 = ~n10950 & n10951;
  assign n14948 = n10821 & n10952;
  assign n14949 = (n10952 & n14877) | (n10952 & n14948) | (n14877 & n14948);
  assign n14950 = n10821 | n10952;
  assign n14951 = n14877 | n14950;
  assign n10955 = ~n14949 & n14951;
  assign n10956 = x65 & x110;
  assign n10957 = n10955 & n10956;
  assign n10958 = n10955 | n10956;
  assign n10959 = ~n10957 & n10958;
  assign n14883 = n10828 | n10830;
  assign n14952 = n10959 & n14883;
  assign n14953 = n10828 & n10959;
  assign n14954 = (n14810 & n14952) | (n14810 & n14953) | (n14952 & n14953);
  assign n14955 = n10959 | n14883;
  assign n14956 = n10828 | n10959;
  assign n14957 = (n14810 & n14955) | (n14810 & n14956) | (n14955 & n14956);
  assign n10962 = ~n14954 & n14957;
  assign n10963 = x64 & x111;
  assign n10964 = n10962 & n10963;
  assign n10965 = n10962 | n10963;
  assign n10966 = ~n10964 & n10965;
  assign n14881 = n10835 | n10837;
  assign n17377 = n10966 & n14881;
  assign n17378 = n10835 & n10966;
  assign n17379 = (n14808 & n17377) | (n14808 & n17378) | (n17377 & n17378);
  assign n17380 = n10966 | n14881;
  assign n17381 = n10835 | n10966;
  assign n17382 = (n14808 & n17380) | (n14808 & n17381) | (n17380 & n17381);
  assign n10969 = ~n17379 & n17382;
  assign n14882 = (n10835 & n14808) | (n10835 & n14881) | (n14808 & n14881);
  assign n10986 = x79 & x97;
  assign n14966 = n10861 | n14894;
  assign n17385 = (n10730 & n14894) | (n10730 & n14966) | (n14894 & n14966);
  assign n14968 = n10986 & n17385;
  assign n17886 = n10986 & n17362;
  assign n17887 = n10986 & n17365;
  assign n17888 = (n17319 & n17886) | (n17319 & n17887) | (n17886 & n17887);
  assign n17387 = (n10861 & n10986) | (n10861 & n17888) | (n10986 & n17888);
  assign n17388 = (n14826 & n14968) | (n14826 & n17387) | (n14968 & n17387);
  assign n17389 = (n14825 & n14968) | (n14825 & n17387) | (n14968 & n17387);
  assign n17390 = (n17281 & n17388) | (n17281 & n17389) | (n17388 & n17389);
  assign n14971 = n10986 | n17385;
  assign n17889 = n10986 | n17362;
  assign n17890 = n10986 | n17365;
  assign n17891 = (n17319 & n17889) | (n17319 & n17890) | (n17889 & n17890);
  assign n17392 = n10861 | n17891;
  assign n17393 = (n14826 & n14971) | (n14826 & n17392) | (n14971 & n17392);
  assign n17394 = (n14825 & n14971) | (n14825 & n17392) | (n14971 & n17392);
  assign n17395 = (n17281 & n17393) | (n17281 & n17394) | (n17393 & n17394);
  assign n10989 = ~n17390 & n17395;
  assign n14975 = n10866 & n10989;
  assign n17396 = (n10868 & n10989) | (n10868 & n14975) | (n10989 & n14975);
  assign n14976 = (n17360 & n17396) | (n17360 & n14975) | (n17396 & n14975);
  assign n14978 = n10866 | n10989;
  assign n17397 = n10868 | n14978;
  assign n14979 = (n17360 & n17397) | (n17360 & n14978) | (n17397 & n14978);
  assign n10992 = ~n14976 & n14979;
  assign n10993 = x78 & x98;
  assign n10994 = n10992 & n10993;
  assign n10995 = n10992 | n10993;
  assign n10996 = ~n10994 & n10995;
  assign n14980 = n10873 & n10996;
  assign n17398 = (n10996 & n14903) | (n10996 & n14980) | (n14903 & n14980);
  assign n17399 = (n10996 & n14902) | (n10996 & n14980) | (n14902 & n14980);
  assign n17400 = (n14815 & n17398) | (n14815 & n17399) | (n17398 & n17399);
  assign n14982 = n10873 | n10996;
  assign n17401 = n14903 | n14982;
  assign n17402 = n14902 | n14982;
  assign n17403 = (n14815 & n17401) | (n14815 & n17402) | (n17401 & n17402);
  assign n10999 = ~n17400 & n17403;
  assign n11000 = x77 & x99;
  assign n11001 = n10999 & n11000;
  assign n11002 = n10999 | n11000;
  assign n11003 = ~n11001 & n11002;
  assign n14961 = n10880 | n10882;
  assign n17404 = n11003 & n14961;
  assign n17383 = n10751 | n10880;
  assign n17384 = (n10880 & n10882) | (n10880 & n17383) | (n10882 & n17383);
  assign n17405 = n11003 & n17384;
  assign n17406 = (n17340 & n17404) | (n17340 & n17405) | (n17404 & n17405);
  assign n17407 = n11003 | n14961;
  assign n17408 = n11003 | n17384;
  assign n17409 = (n17340 & n17407) | (n17340 & n17408) | (n17407 & n17408);
  assign n11006 = ~n17406 & n17409;
  assign n11007 = x76 & x100;
  assign n11008 = n11006 & n11007;
  assign n11009 = n11006 | n11007;
  assign n11010 = ~n11008 & n11009;
  assign n14984 = n10887 & n11010;
  assign n17410 = (n11010 & n14912) | (n11010 & n14984) | (n14912 & n14984);
  assign n17411 = (n10889 & n11010) | (n10889 & n14984) | (n11010 & n14984);
  assign n17412 = (n14840 & n17410) | (n14840 & n17411) | (n17410 & n17411);
  assign n14986 = n10887 | n11010;
  assign n17413 = n14912 | n14986;
  assign n17414 = n10889 | n14986;
  assign n17415 = (n14840 & n17413) | (n14840 & n17414) | (n17413 & n17414);
  assign n11013 = ~n17412 & n17415;
  assign n11014 = x75 & x101;
  assign n11015 = n11013 & n11014;
  assign n11016 = n11013 | n11014;
  assign n11017 = ~n11015 & n11016;
  assign n14988 = n10894 & n11017;
  assign n14989 = (n11017 & n14917) | (n11017 & n14988) | (n14917 & n14988);
  assign n14990 = n10894 | n11017;
  assign n14991 = n14917 | n14990;
  assign n11020 = ~n14989 & n14991;
  assign n11021 = x74 & x102;
  assign n11022 = n11020 & n11021;
  assign n11023 = n11020 | n11021;
  assign n11024 = ~n11022 & n11023;
  assign n14992 = n10901 & n11024;
  assign n14993 = (n11024 & n14921) | (n11024 & n14992) | (n14921 & n14992);
  assign n14994 = n10901 | n11024;
  assign n14995 = n14921 | n14994;
  assign n11027 = ~n14993 & n14995;
  assign n11028 = x73 & x103;
  assign n11029 = n11027 & n11028;
  assign n11030 = n11027 | n11028;
  assign n11031 = ~n11029 & n11030;
  assign n14996 = n10908 & n11031;
  assign n14997 = (n11031 & n14925) | (n11031 & n14996) | (n14925 & n14996);
  assign n14998 = n10908 | n11031;
  assign n14999 = n14925 | n14998;
  assign n11034 = ~n14997 & n14999;
  assign n11035 = x72 & x104;
  assign n11036 = n11034 & n11035;
  assign n11037 = n11034 | n11035;
  assign n11038 = ~n11036 & n11037;
  assign n15000 = n10915 & n11038;
  assign n15001 = (n11038 & n14929) | (n11038 & n15000) | (n14929 & n15000);
  assign n15002 = n10915 | n11038;
  assign n15003 = n14929 | n15002;
  assign n11041 = ~n15001 & n15003;
  assign n11042 = x71 & x105;
  assign n11043 = n11041 & n11042;
  assign n11044 = n11041 | n11042;
  assign n11045 = ~n11043 & n11044;
  assign n15004 = n10922 & n11045;
  assign n15005 = (n11045 & n14933) | (n11045 & n15004) | (n14933 & n15004);
  assign n15006 = n10922 | n11045;
  assign n15007 = n14933 | n15006;
  assign n11048 = ~n15005 & n15007;
  assign n11049 = x70 & x106;
  assign n11050 = n11048 & n11049;
  assign n11051 = n11048 | n11049;
  assign n11052 = ~n11050 & n11051;
  assign n15008 = n10929 & n11052;
  assign n15009 = (n11052 & n14937) | (n11052 & n15008) | (n14937 & n15008);
  assign n15010 = n10929 | n11052;
  assign n15011 = n14937 | n15010;
  assign n11055 = ~n15009 & n15011;
  assign n11056 = x69 & x107;
  assign n11057 = n11055 & n11056;
  assign n11058 = n11055 | n11056;
  assign n11059 = ~n11057 & n11058;
  assign n15012 = n10936 & n11059;
  assign n15013 = (n11059 & n14941) | (n11059 & n15012) | (n14941 & n15012);
  assign n15014 = n10936 | n11059;
  assign n15015 = n14941 | n15014;
  assign n11062 = ~n15013 & n15015;
  assign n11063 = x68 & x108;
  assign n11064 = n11062 & n11063;
  assign n11065 = n11062 | n11063;
  assign n11066 = ~n11064 & n11065;
  assign n15016 = n10943 & n11066;
  assign n15017 = (n11066 & n14945) | (n11066 & n15016) | (n14945 & n15016);
  assign n15018 = n10943 | n11066;
  assign n15019 = n14945 | n15018;
  assign n11069 = ~n15017 & n15019;
  assign n11070 = x67 & x109;
  assign n11071 = n11069 & n11070;
  assign n11072 = n11069 | n11070;
  assign n11073 = ~n11071 & n11072;
  assign n15020 = n10950 & n11073;
  assign n15021 = (n11073 & n14949) | (n11073 & n15020) | (n14949 & n15020);
  assign n15022 = n10950 | n11073;
  assign n15023 = n14949 | n15022;
  assign n11076 = ~n15021 & n15023;
  assign n11077 = x66 & x110;
  assign n11078 = n11076 & n11077;
  assign n11079 = n11076 | n11077;
  assign n11080 = ~n11078 & n11079;
  assign n15024 = n10957 & n11080;
  assign n15025 = (n11080 & n14954) | (n11080 & n15024) | (n14954 & n15024);
  assign n15026 = n10957 | n11080;
  assign n15027 = n14954 | n15026;
  assign n11083 = ~n15025 & n15027;
  assign n11084 = x65 & x111;
  assign n11085 = n11083 & n11084;
  assign n11086 = n11083 | n11084;
  assign n11087 = ~n11085 & n11086;
  assign n14958 = n10964 | n10966;
  assign n15028 = n11087 & n14958;
  assign n15029 = n10964 & n11087;
  assign n15030 = (n14882 & n15028) | (n14882 & n15029) | (n15028 & n15029);
  assign n15031 = n11087 | n14958;
  assign n15032 = n10964 | n11087;
  assign n15033 = (n14882 & n15031) | (n14882 & n15032) | (n15031 & n15032);
  assign n11090 = ~n15030 & n15033;
  assign n14962 = (n17340 & n17384) | (n17340 & n14961) | (n17384 & n14961);
  assign n15037 = n10994 | n10996;
  assign n17416 = n10873 | n10994;
  assign n17417 = (n10994 & n10996) | (n10994 & n17416) | (n10996 & n17416);
  assign n17418 = (n14903 & n15037) | (n14903 & n17417) | (n15037 & n17417);
  assign n17419 = (n14902 & n15037) | (n14902 & n17417) | (n15037 & n17417);
  assign n17420 = (n14815 & n17418) | (n14815 & n17419) | (n17418 & n17419);
  assign n11106 = x79 & x98;
  assign n15039 = n11106 & n17390;
  assign n17421 = (n11106 & n15039) | (n11106 & n17396) | (n15039 & n17396);
  assign n17892 = (n10989 & n11106) | (n10989 & n15039) | (n11106 & n15039);
  assign n17893 = n11106 & n15039;
  assign n17894 = (n10866 & n17892) | (n10866 & n17893) | (n17892 & n17893);
  assign n17423 = (n17360 & n17421) | (n17360 & n17894) | (n17421 & n17894);
  assign n15041 = n11106 | n17390;
  assign n17424 = n15041 | n17396;
  assign n17895 = n10989 | n15041;
  assign n17896 = (n10866 & n15041) | (n10866 & n17895) | (n15041 & n17895);
  assign n17426 = (n17360 & n17424) | (n17360 & n17896) | (n17424 & n17896);
  assign n11109 = ~n17423 & n17426;
  assign n11110 = n17420 & n11109;
  assign n11111 = n17420 | n11109;
  assign n11112 = ~n11110 & n11111;
  assign n11113 = x78 & x99;
  assign n11114 = n11112 & n11113;
  assign n11115 = n11112 | n11113;
  assign n11116 = ~n11114 & n11115;
  assign n15034 = n11001 | n11003;
  assign n15043 = n11116 & n15034;
  assign n15044 = n11001 & n11116;
  assign n15045 = (n14962 & n15043) | (n14962 & n15044) | (n15043 & n15044);
  assign n15046 = n11116 | n15034;
  assign n15047 = n11001 | n11116;
  assign n15048 = (n14962 & n15046) | (n14962 & n15047) | (n15046 & n15047);
  assign n11119 = ~n15045 & n15048;
  assign n11120 = x77 & x100;
  assign n11121 = n11119 & n11120;
  assign n11122 = n11119 | n11120;
  assign n11123 = ~n11121 & n11122;
  assign n15049 = n11008 & n11123;
  assign n15050 = (n11123 & n17412) | (n11123 & n15049) | (n17412 & n15049);
  assign n15051 = n11008 | n11123;
  assign n15052 = n17412 | n15051;
  assign n11126 = ~n15050 & n15052;
  assign n11127 = x76 & x101;
  assign n11128 = n11126 & n11127;
  assign n11129 = n11126 | n11127;
  assign n11130 = ~n11128 & n11129;
  assign n15053 = n11015 & n11130;
  assign n15054 = (n11130 & n14989) | (n11130 & n15053) | (n14989 & n15053);
  assign n15055 = n11015 | n11130;
  assign n15056 = n14989 | n15055;
  assign n11133 = ~n15054 & n15056;
  assign n11134 = x75 & x102;
  assign n11135 = n11133 & n11134;
  assign n11136 = n11133 | n11134;
  assign n11137 = ~n11135 & n11136;
  assign n15057 = n11022 & n11137;
  assign n15058 = (n11137 & n14993) | (n11137 & n15057) | (n14993 & n15057);
  assign n15059 = n11022 | n11137;
  assign n15060 = n14993 | n15059;
  assign n11140 = ~n15058 & n15060;
  assign n11141 = x74 & x103;
  assign n11142 = n11140 & n11141;
  assign n11143 = n11140 | n11141;
  assign n11144 = ~n11142 & n11143;
  assign n15061 = n11029 & n11144;
  assign n15062 = (n11144 & n14997) | (n11144 & n15061) | (n14997 & n15061);
  assign n15063 = n11029 | n11144;
  assign n15064 = n14997 | n15063;
  assign n11147 = ~n15062 & n15064;
  assign n11148 = x73 & x104;
  assign n11149 = n11147 & n11148;
  assign n11150 = n11147 | n11148;
  assign n11151 = ~n11149 & n11150;
  assign n15065 = n11036 & n11151;
  assign n15066 = (n11151 & n15001) | (n11151 & n15065) | (n15001 & n15065);
  assign n15067 = n11036 | n11151;
  assign n15068 = n15001 | n15067;
  assign n11154 = ~n15066 & n15068;
  assign n11155 = x72 & x105;
  assign n11156 = n11154 & n11155;
  assign n11157 = n11154 | n11155;
  assign n11158 = ~n11156 & n11157;
  assign n15069 = n11043 & n11158;
  assign n15070 = (n11158 & n15005) | (n11158 & n15069) | (n15005 & n15069);
  assign n15071 = n11043 | n11158;
  assign n15072 = n15005 | n15071;
  assign n11161 = ~n15070 & n15072;
  assign n11162 = x71 & x106;
  assign n11163 = n11161 & n11162;
  assign n11164 = n11161 | n11162;
  assign n11165 = ~n11163 & n11164;
  assign n15073 = n11050 & n11165;
  assign n15074 = (n11165 & n15009) | (n11165 & n15073) | (n15009 & n15073);
  assign n15075 = n11050 | n11165;
  assign n15076 = n15009 | n15075;
  assign n11168 = ~n15074 & n15076;
  assign n11169 = x70 & x107;
  assign n11170 = n11168 & n11169;
  assign n11171 = n11168 | n11169;
  assign n11172 = ~n11170 & n11171;
  assign n15077 = n11057 & n11172;
  assign n15078 = (n11172 & n15013) | (n11172 & n15077) | (n15013 & n15077);
  assign n15079 = n11057 | n11172;
  assign n15080 = n15013 | n15079;
  assign n11175 = ~n15078 & n15080;
  assign n11176 = x69 & x108;
  assign n11177 = n11175 & n11176;
  assign n11178 = n11175 | n11176;
  assign n11179 = ~n11177 & n11178;
  assign n15081 = n11064 & n11179;
  assign n15082 = (n11179 & n15017) | (n11179 & n15081) | (n15017 & n15081);
  assign n15083 = n11064 | n11179;
  assign n15084 = n15017 | n15083;
  assign n11182 = ~n15082 & n15084;
  assign n11183 = x68 & x109;
  assign n11184 = n11182 & n11183;
  assign n11185 = n11182 | n11183;
  assign n11186 = ~n11184 & n11185;
  assign n15085 = n11071 & n11186;
  assign n15086 = (n11186 & n15021) | (n11186 & n15085) | (n15021 & n15085);
  assign n15087 = n11071 | n11186;
  assign n15088 = n15021 | n15087;
  assign n11189 = ~n15086 & n15088;
  assign n11190 = x67 & x110;
  assign n11191 = n11189 & n11190;
  assign n11192 = n11189 | n11190;
  assign n11193 = ~n11191 & n11192;
  assign n15089 = n11078 & n11193;
  assign n15090 = (n11193 & n15025) | (n11193 & n15089) | (n15025 & n15089);
  assign n15091 = n11078 | n11193;
  assign n15092 = n15025 | n15091;
  assign n11196 = ~n15090 & n15092;
  assign n11197 = x66 & x111;
  assign n11198 = n11196 & n11197;
  assign n11199 = n11196 | n11197;
  assign n11200 = ~n11198 & n11199;
  assign n15093 = n11085 & n11200;
  assign n15094 = (n11200 & n15030) | (n11200 & n15093) | (n15030 & n15093);
  assign n15095 = n11085 | n11200;
  assign n15096 = n15030 | n15095;
  assign n11203 = ~n15094 & n15096;
  assign n11218 = x79 & x99;
  assign n17899 = n11218 & n15039;
  assign n17900 = n11106 & n11218;
  assign n17901 = (n17396 & n17899) | (n17396 & n17900) | (n17899 & n17900);
  assign n17897 = n11218 & n17894;
  assign n17898 = (n17360 & n17901) | (n17360 & n17897) | (n17901 & n17897);
  assign n17430 = (n11109 & n11218) | (n11109 & n17898) | (n11218 & n17898);
  assign n17432 = n11218 & n17894;
  assign n17433 = (n17360 & n17901) | (n17360 & n17432) | (n17901 & n17432);
  assign n15104 = (n17420 & n17430) | (n17420 & n17433) | (n17430 & n17433);
  assign n17904 = n11218 | n15039;
  assign n17905 = n11106 | n11218;
  assign n17906 = (n17396 & n17904) | (n17396 & n17905) | (n17904 & n17905);
  assign n17902 = n11218 | n17894;
  assign n17903 = (n17360 & n17906) | (n17360 & n17902) | (n17906 & n17902);
  assign n17435 = n11109 | n17903;
  assign n17437 = n11218 | n17894;
  assign n17438 = (n17360 & n17906) | (n17360 & n17437) | (n17906 & n17437);
  assign n15107 = (n17420 & n17435) | (n17420 & n17438) | (n17435 & n17438);
  assign n11221 = ~n15104 & n15107;
  assign n15108 = n11114 & n11221;
  assign n17439 = (n11221 & n15044) | (n11221 & n15108) | (n15044 & n15108);
  assign n17440 = (n11221 & n15043) | (n11221 & n15108) | (n15043 & n15108);
  assign n17441 = (n14962 & n17439) | (n14962 & n17440) | (n17439 & n17440);
  assign n15110 = n11114 | n11221;
  assign n17442 = n15044 | n15110;
  assign n17443 = n15043 | n15110;
  assign n17444 = (n14962 & n17442) | (n14962 & n17443) | (n17442 & n17443);
  assign n11224 = ~n17441 & n17444;
  assign n11225 = x78 & x100;
  assign n11226 = n11224 & n11225;
  assign n11227 = n11224 | n11225;
  assign n11228 = ~n11226 & n11227;
  assign n15098 = n11121 | n11123;
  assign n17445 = n11228 & n15098;
  assign n17427 = n11008 | n11121;
  assign n17428 = (n11121 & n11123) | (n11121 & n17427) | (n11123 & n17427);
  assign n17446 = n11228 & n17428;
  assign n17447 = (n17412 & n17445) | (n17412 & n17446) | (n17445 & n17446);
  assign n17448 = n11228 | n15098;
  assign n17449 = n11228 | n17428;
  assign n17450 = (n17412 & n17448) | (n17412 & n17449) | (n17448 & n17449);
  assign n11231 = ~n17447 & n17450;
  assign n11232 = x77 & x101;
  assign n11233 = n11231 & n11232;
  assign n11234 = n11231 | n11232;
  assign n11235 = ~n11233 & n11234;
  assign n15112 = n11128 & n11235;
  assign n17451 = (n11235 & n15053) | (n11235 & n15112) | (n15053 & n15112);
  assign n17452 = (n11130 & n11235) | (n11130 & n15112) | (n11235 & n15112);
  assign n17453 = (n14989 & n17451) | (n14989 & n17452) | (n17451 & n17452);
  assign n15114 = n11128 | n11235;
  assign n17454 = n15053 | n15114;
  assign n17455 = n11130 | n15114;
  assign n17456 = (n14989 & n17454) | (n14989 & n17455) | (n17454 & n17455);
  assign n11238 = ~n17453 & n17456;
  assign n11239 = x76 & x102;
  assign n11240 = n11238 & n11239;
  assign n11241 = n11238 | n11239;
  assign n11242 = ~n11240 & n11241;
  assign n15116 = n11135 & n11242;
  assign n15117 = (n11242 & n15058) | (n11242 & n15116) | (n15058 & n15116);
  assign n15118 = n11135 | n11242;
  assign n15119 = n15058 | n15118;
  assign n11245 = ~n15117 & n15119;
  assign n11246 = x75 & x103;
  assign n11247 = n11245 & n11246;
  assign n11248 = n11245 | n11246;
  assign n11249 = ~n11247 & n11248;
  assign n15120 = n11142 & n11249;
  assign n15121 = (n11249 & n15062) | (n11249 & n15120) | (n15062 & n15120);
  assign n15122 = n11142 | n11249;
  assign n15123 = n15062 | n15122;
  assign n11252 = ~n15121 & n15123;
  assign n11253 = x74 & x104;
  assign n11254 = n11252 & n11253;
  assign n11255 = n11252 | n11253;
  assign n11256 = ~n11254 & n11255;
  assign n15124 = n11149 & n11256;
  assign n15125 = (n11256 & n15066) | (n11256 & n15124) | (n15066 & n15124);
  assign n15126 = n11149 | n11256;
  assign n15127 = n15066 | n15126;
  assign n11259 = ~n15125 & n15127;
  assign n11260 = x73 & x105;
  assign n11261 = n11259 & n11260;
  assign n11262 = n11259 | n11260;
  assign n11263 = ~n11261 & n11262;
  assign n15128 = n11156 & n11263;
  assign n15129 = (n11263 & n15070) | (n11263 & n15128) | (n15070 & n15128);
  assign n15130 = n11156 | n11263;
  assign n15131 = n15070 | n15130;
  assign n11266 = ~n15129 & n15131;
  assign n11267 = x72 & x106;
  assign n11268 = n11266 & n11267;
  assign n11269 = n11266 | n11267;
  assign n11270 = ~n11268 & n11269;
  assign n15132 = n11163 & n11270;
  assign n15133 = (n11270 & n15074) | (n11270 & n15132) | (n15074 & n15132);
  assign n15134 = n11163 | n11270;
  assign n15135 = n15074 | n15134;
  assign n11273 = ~n15133 & n15135;
  assign n11274 = x71 & x107;
  assign n11275 = n11273 & n11274;
  assign n11276 = n11273 | n11274;
  assign n11277 = ~n11275 & n11276;
  assign n15136 = n11170 & n11277;
  assign n15137 = (n11277 & n15078) | (n11277 & n15136) | (n15078 & n15136);
  assign n15138 = n11170 | n11277;
  assign n15139 = n15078 | n15138;
  assign n11280 = ~n15137 & n15139;
  assign n11281 = x70 & x108;
  assign n11282 = n11280 & n11281;
  assign n11283 = n11280 | n11281;
  assign n11284 = ~n11282 & n11283;
  assign n15140 = n11177 & n11284;
  assign n15141 = (n11284 & n15082) | (n11284 & n15140) | (n15082 & n15140);
  assign n15142 = n11177 | n11284;
  assign n15143 = n15082 | n15142;
  assign n11287 = ~n15141 & n15143;
  assign n11288 = x69 & x109;
  assign n11289 = n11287 & n11288;
  assign n11290 = n11287 | n11288;
  assign n11291 = ~n11289 & n11290;
  assign n15144 = n11184 & n11291;
  assign n15145 = (n11291 & n15086) | (n11291 & n15144) | (n15086 & n15144);
  assign n15146 = n11184 | n11291;
  assign n15147 = n15086 | n15146;
  assign n11294 = ~n15145 & n15147;
  assign n11295 = x68 & x110;
  assign n11296 = n11294 & n11295;
  assign n11297 = n11294 | n11295;
  assign n11298 = ~n11296 & n11297;
  assign n15148 = n11191 & n11298;
  assign n15149 = (n11298 & n15090) | (n11298 & n15148) | (n15090 & n15148);
  assign n15150 = n11191 | n11298;
  assign n15151 = n15090 | n15150;
  assign n11301 = ~n15149 & n15151;
  assign n11302 = x67 & x111;
  assign n11303 = n11301 & n11302;
  assign n11304 = n11301 | n11302;
  assign n11305 = ~n11303 & n11304;
  assign n15152 = n11198 & n11305;
  assign n15153 = (n11305 & n15094) | (n11305 & n15152) | (n15094 & n15152);
  assign n15154 = n11198 | n11305;
  assign n15155 = n15094 | n15154;
  assign n11308 = ~n15153 & n15155;
  assign n11322 = x79 & x100;
  assign n15159 = n11221 | n15104;
  assign n17457 = (n11114 & n15104) | (n11114 & n15159) | (n15104 & n15159);
  assign n15161 = n11322 & n17457;
  assign n17907 = n11322 & n17430;
  assign n17908 = n11322 & n17433;
  assign n17909 = (n17420 & n17907) | (n17420 & n17908) | (n17907 & n17908);
  assign n17459 = (n11221 & n11322) | (n11221 & n17909) | (n11322 & n17909);
  assign n17460 = (n15044 & n15161) | (n15044 & n17459) | (n15161 & n17459);
  assign n17461 = (n15043 & n15161) | (n15043 & n17459) | (n15161 & n17459);
  assign n17462 = (n14962 & n17460) | (n14962 & n17461) | (n17460 & n17461);
  assign n15164 = n11322 | n17457;
  assign n17910 = n11322 | n17430;
  assign n17911 = n11322 | n17433;
  assign n17912 = (n17420 & n17910) | (n17420 & n17911) | (n17910 & n17911);
  assign n17464 = n11221 | n17912;
  assign n17465 = (n15044 & n15164) | (n15044 & n17464) | (n15164 & n17464);
  assign n17466 = (n15043 & n15164) | (n15043 & n17464) | (n15164 & n17464);
  assign n17467 = (n14962 & n17465) | (n14962 & n17466) | (n17465 & n17466);
  assign n11325 = ~n17462 & n17467;
  assign n15168 = n11226 & n11325;
  assign n17468 = (n11228 & n11325) | (n11228 & n15168) | (n11325 & n15168);
  assign n17469 = (n15098 & n15168) | (n15098 & n17468) | (n15168 & n17468);
  assign n17470 = (n15168 & n17428) | (n15168 & n17468) | (n17428 & n17468);
  assign n17471 = (n17412 & n17469) | (n17412 & n17470) | (n17469 & n17470);
  assign n15171 = n11226 | n11325;
  assign n17472 = n11228 | n15171;
  assign n17473 = (n15098 & n15171) | (n15098 & n17472) | (n15171 & n17472);
  assign n17474 = (n15171 & n17428) | (n15171 & n17472) | (n17428 & n17472);
  assign n17475 = (n17412 & n17473) | (n17412 & n17474) | (n17473 & n17474);
  assign n11328 = ~n17471 & n17475;
  assign n11329 = x78 & x101;
  assign n11330 = n11328 & n11329;
  assign n11331 = n11328 | n11329;
  assign n11332 = ~n11330 & n11331;
  assign n15173 = n11233 & n11332;
  assign n15174 = (n11332 & n17453) | (n11332 & n15173) | (n17453 & n15173);
  assign n15175 = n11233 | n11332;
  assign n15176 = n17453 | n15175;
  assign n11335 = ~n15174 & n15176;
  assign n11336 = x77 & x102;
  assign n11337 = n11335 & n11336;
  assign n11338 = n11335 | n11336;
  assign n11339 = ~n11337 & n11338;
  assign n15177 = n11240 & n11339;
  assign n15178 = (n11339 & n15117) | (n11339 & n15177) | (n15117 & n15177);
  assign n15179 = n11240 | n11339;
  assign n15180 = n15117 | n15179;
  assign n11342 = ~n15178 & n15180;
  assign n11343 = x76 & x103;
  assign n11344 = n11342 & n11343;
  assign n11345 = n11342 | n11343;
  assign n11346 = ~n11344 & n11345;
  assign n15181 = n11247 & n11346;
  assign n15182 = (n11346 & n15121) | (n11346 & n15181) | (n15121 & n15181);
  assign n15183 = n11247 | n11346;
  assign n15184 = n15121 | n15183;
  assign n11349 = ~n15182 & n15184;
  assign n11350 = x75 & x104;
  assign n11351 = n11349 & n11350;
  assign n11352 = n11349 | n11350;
  assign n11353 = ~n11351 & n11352;
  assign n15185 = n11254 & n11353;
  assign n15186 = (n11353 & n15125) | (n11353 & n15185) | (n15125 & n15185);
  assign n15187 = n11254 | n11353;
  assign n15188 = n15125 | n15187;
  assign n11356 = ~n15186 & n15188;
  assign n11357 = x74 & x105;
  assign n11358 = n11356 & n11357;
  assign n11359 = n11356 | n11357;
  assign n11360 = ~n11358 & n11359;
  assign n15189 = n11261 & n11360;
  assign n15190 = (n11360 & n15129) | (n11360 & n15189) | (n15129 & n15189);
  assign n15191 = n11261 | n11360;
  assign n15192 = n15129 | n15191;
  assign n11363 = ~n15190 & n15192;
  assign n11364 = x73 & x106;
  assign n11365 = n11363 & n11364;
  assign n11366 = n11363 | n11364;
  assign n11367 = ~n11365 & n11366;
  assign n15193 = n11268 & n11367;
  assign n15194 = (n11367 & n15133) | (n11367 & n15193) | (n15133 & n15193);
  assign n15195 = n11268 | n11367;
  assign n15196 = n15133 | n15195;
  assign n11370 = ~n15194 & n15196;
  assign n11371 = x72 & x107;
  assign n11372 = n11370 & n11371;
  assign n11373 = n11370 | n11371;
  assign n11374 = ~n11372 & n11373;
  assign n15197 = n11275 & n11374;
  assign n15198 = (n11374 & n15137) | (n11374 & n15197) | (n15137 & n15197);
  assign n15199 = n11275 | n11374;
  assign n15200 = n15137 | n15199;
  assign n11377 = ~n15198 & n15200;
  assign n11378 = x71 & x108;
  assign n11379 = n11377 & n11378;
  assign n11380 = n11377 | n11378;
  assign n11381 = ~n11379 & n11380;
  assign n15201 = n11282 & n11381;
  assign n15202 = (n11381 & n15141) | (n11381 & n15201) | (n15141 & n15201);
  assign n15203 = n11282 | n11381;
  assign n15204 = n15141 | n15203;
  assign n11384 = ~n15202 & n15204;
  assign n11385 = x70 & x109;
  assign n11386 = n11384 & n11385;
  assign n11387 = n11384 | n11385;
  assign n11388 = ~n11386 & n11387;
  assign n15205 = n11289 & n11388;
  assign n15206 = (n11388 & n15145) | (n11388 & n15205) | (n15145 & n15205);
  assign n15207 = n11289 | n11388;
  assign n15208 = n15145 | n15207;
  assign n11391 = ~n15206 & n15208;
  assign n11392 = x69 & x110;
  assign n11393 = n11391 & n11392;
  assign n11394 = n11391 | n11392;
  assign n11395 = ~n11393 & n11394;
  assign n15209 = n11296 & n11395;
  assign n15210 = (n11395 & n15149) | (n11395 & n15209) | (n15149 & n15209);
  assign n15211 = n11296 | n11395;
  assign n15212 = n15149 | n15211;
  assign n11398 = ~n15210 & n15212;
  assign n11399 = x68 & x111;
  assign n11400 = n11398 & n11399;
  assign n11401 = n11398 | n11399;
  assign n11402 = ~n11400 & n11401;
  assign n15213 = n11303 & n11402;
  assign n15214 = (n11402 & n15153) | (n11402 & n15213) | (n15153 & n15213);
  assign n15215 = n11303 | n11402;
  assign n15216 = n15153 | n15215;
  assign n11405 = ~n15214 & n15216;
  assign n11418 = x79 & x101;
  assign n15220 = n11418 & n17462;
  assign n15221 = (n11418 & n17471) | (n11418 & n15220) | (n17471 & n15220);
  assign n15222 = n11418 | n17462;
  assign n15223 = n17471 | n15222;
  assign n11421 = ~n15221 & n15223;
  assign n17913 = n11330 & n11421;
  assign n17914 = (n11332 & n11421) | (n11332 & n17913) | (n11421 & n17913);
  assign n17476 = n11233 | n11330;
  assign n17477 = (n11330 & n11332) | (n11330 & n17476) | (n11332 & n17476);
  assign n17479 = n11421 & n17477;
  assign n17480 = (n17453 & n17914) | (n17453 & n17479) | (n17914 & n17479);
  assign n17915 = n11330 | n11421;
  assign n17916 = n11332 | n17915;
  assign n17482 = n11421 | n17477;
  assign n17483 = (n17453 & n17916) | (n17453 & n17482) | (n17916 & n17482);
  assign n11424 = ~n17480 & n17483;
  assign n11425 = x78 & x102;
  assign n11426 = n11424 & n11425;
  assign n11427 = n11424 | n11425;
  assign n11428 = ~n11426 & n11427;
  assign n15224 = n11337 & n11428;
  assign n17484 = (n11428 & n15177) | (n11428 & n15224) | (n15177 & n15224);
  assign n17485 = (n11339 & n11428) | (n11339 & n15224) | (n11428 & n15224);
  assign n17486 = (n15117 & n17484) | (n15117 & n17485) | (n17484 & n17485);
  assign n15226 = n11337 | n11428;
  assign n17487 = n15177 | n15226;
  assign n17488 = n11339 | n15226;
  assign n17489 = (n15117 & n17487) | (n15117 & n17488) | (n17487 & n17488);
  assign n11431 = ~n17486 & n17489;
  assign n11432 = x77 & x103;
  assign n11433 = n11431 & n11432;
  assign n11434 = n11431 | n11432;
  assign n11435 = ~n11433 & n11434;
  assign n15228 = n11344 & n11435;
  assign n15229 = (n11435 & n15182) | (n11435 & n15228) | (n15182 & n15228);
  assign n15230 = n11344 | n11435;
  assign n15231 = n15182 | n15230;
  assign n11438 = ~n15229 & n15231;
  assign n11439 = x76 & x104;
  assign n11440 = n11438 & n11439;
  assign n11441 = n11438 | n11439;
  assign n11442 = ~n11440 & n11441;
  assign n15232 = n11351 & n11442;
  assign n15233 = (n11442 & n15186) | (n11442 & n15232) | (n15186 & n15232);
  assign n15234 = n11351 | n11442;
  assign n15235 = n15186 | n15234;
  assign n11445 = ~n15233 & n15235;
  assign n11446 = x75 & x105;
  assign n11447 = n11445 & n11446;
  assign n11448 = n11445 | n11446;
  assign n11449 = ~n11447 & n11448;
  assign n15236 = n11358 & n11449;
  assign n15237 = (n11449 & n15190) | (n11449 & n15236) | (n15190 & n15236);
  assign n15238 = n11358 | n11449;
  assign n15239 = n15190 | n15238;
  assign n11452 = ~n15237 & n15239;
  assign n11453 = x74 & x106;
  assign n11454 = n11452 & n11453;
  assign n11455 = n11452 | n11453;
  assign n11456 = ~n11454 & n11455;
  assign n15240 = n11365 & n11456;
  assign n15241 = (n11456 & n15194) | (n11456 & n15240) | (n15194 & n15240);
  assign n15242 = n11365 | n11456;
  assign n15243 = n15194 | n15242;
  assign n11459 = ~n15241 & n15243;
  assign n11460 = x73 & x107;
  assign n11461 = n11459 & n11460;
  assign n11462 = n11459 | n11460;
  assign n11463 = ~n11461 & n11462;
  assign n15244 = n11372 & n11463;
  assign n15245 = (n11463 & n15198) | (n11463 & n15244) | (n15198 & n15244);
  assign n15246 = n11372 | n11463;
  assign n15247 = n15198 | n15246;
  assign n11466 = ~n15245 & n15247;
  assign n11467 = x72 & x108;
  assign n11468 = n11466 & n11467;
  assign n11469 = n11466 | n11467;
  assign n11470 = ~n11468 & n11469;
  assign n15248 = n11379 & n11470;
  assign n15249 = (n11470 & n15202) | (n11470 & n15248) | (n15202 & n15248);
  assign n15250 = n11379 | n11470;
  assign n15251 = n15202 | n15250;
  assign n11473 = ~n15249 & n15251;
  assign n11474 = x71 & x109;
  assign n11475 = n11473 & n11474;
  assign n11476 = n11473 | n11474;
  assign n11477 = ~n11475 & n11476;
  assign n15252 = n11386 & n11477;
  assign n15253 = (n11477 & n15206) | (n11477 & n15252) | (n15206 & n15252);
  assign n15254 = n11386 | n11477;
  assign n15255 = n15206 | n15254;
  assign n11480 = ~n15253 & n15255;
  assign n11481 = x70 & x110;
  assign n11482 = n11480 & n11481;
  assign n11483 = n11480 | n11481;
  assign n11484 = ~n11482 & n11483;
  assign n15256 = n11393 & n11484;
  assign n15257 = (n11484 & n15210) | (n11484 & n15256) | (n15210 & n15256);
  assign n15258 = n11393 | n11484;
  assign n15259 = n15210 | n15258;
  assign n11487 = ~n15257 & n15259;
  assign n11488 = x69 & x111;
  assign n11489 = n11487 & n11488;
  assign n11490 = n11487 | n11488;
  assign n11491 = ~n11489 & n11490;
  assign n15260 = n11400 & n11491;
  assign n15261 = (n11491 & n15214) | (n11491 & n15260) | (n15214 & n15260);
  assign n15262 = n11400 | n11491;
  assign n15263 = n15214 | n15262;
  assign n11494 = ~n15261 & n15263;
  assign n15218 = n11330 | n11332;
  assign n11506 = x79 & x102;
  assign n17492 = n11418 & n11506;
  assign n17917 = n17462 & n17492;
  assign n17493 = (n17471 & n17917) | (n17471 & n17492) | (n17917 & n17492);
  assign n17490 = (n11421 & n11506) | (n11421 & n17493) | (n11506 & n17493);
  assign n17494 = (n15218 & n17490) | (n15218 & n17493) | (n17490 & n17493);
  assign n17495 = (n17477 & n17490) | (n17477 & n17493) | (n17490 & n17493);
  assign n17496 = (n17453 & n17494) | (n17453 & n17495) | (n17494 & n17495);
  assign n17499 = n11418 | n11506;
  assign n17918 = (n11506 & n17462) | (n11506 & n17499) | (n17462 & n17499);
  assign n17500 = (n17471 & n17918) | (n17471 & n17499) | (n17918 & n17499);
  assign n17497 = n11421 | n17500;
  assign n17501 = (n15218 & n17497) | (n15218 & n17500) | (n17497 & n17500);
  assign n17502 = (n17477 & n17497) | (n17477 & n17500) | (n17497 & n17500);
  assign n17503 = (n17453 & n17501) | (n17453 & n17502) | (n17501 & n17502);
  assign n11509 = ~n17496 & n17503;
  assign n15272 = n11426 & n11509;
  assign n15273 = (n11509 & n17486) | (n11509 & n15272) | (n17486 & n15272);
  assign n15274 = n11426 | n11509;
  assign n15275 = n17486 | n15274;
  assign n11512 = ~n15273 & n15275;
  assign n11513 = x78 & x103;
  assign n11514 = n11512 & n11513;
  assign n11515 = n11512 | n11513;
  assign n11516 = ~n11514 & n11515;
  assign n15276 = n11433 & n11516;
  assign n15277 = (n11516 & n15229) | (n11516 & n15276) | (n15229 & n15276);
  assign n15278 = n11433 | n11516;
  assign n15279 = n15229 | n15278;
  assign n11519 = ~n15277 & n15279;
  assign n11520 = x77 & x104;
  assign n11521 = n11519 & n11520;
  assign n11522 = n11519 | n11520;
  assign n11523 = ~n11521 & n11522;
  assign n15280 = n11440 & n11523;
  assign n15281 = (n11523 & n15233) | (n11523 & n15280) | (n15233 & n15280);
  assign n15282 = n11440 | n11523;
  assign n15283 = n15233 | n15282;
  assign n11526 = ~n15281 & n15283;
  assign n11527 = x76 & x105;
  assign n11528 = n11526 & n11527;
  assign n11529 = n11526 | n11527;
  assign n11530 = ~n11528 & n11529;
  assign n15284 = n11447 & n11530;
  assign n15285 = (n11530 & n15237) | (n11530 & n15284) | (n15237 & n15284);
  assign n15286 = n11447 | n11530;
  assign n15287 = n15237 | n15286;
  assign n11533 = ~n15285 & n15287;
  assign n11534 = x75 & x106;
  assign n11535 = n11533 & n11534;
  assign n11536 = n11533 | n11534;
  assign n11537 = ~n11535 & n11536;
  assign n15288 = n11454 & n11537;
  assign n15289 = (n11537 & n15241) | (n11537 & n15288) | (n15241 & n15288);
  assign n15290 = n11454 | n11537;
  assign n15291 = n15241 | n15290;
  assign n11540 = ~n15289 & n15291;
  assign n11541 = x74 & x107;
  assign n11542 = n11540 & n11541;
  assign n11543 = n11540 | n11541;
  assign n11544 = ~n11542 & n11543;
  assign n15292 = n11461 & n11544;
  assign n15293 = (n11544 & n15245) | (n11544 & n15292) | (n15245 & n15292);
  assign n15294 = n11461 | n11544;
  assign n15295 = n15245 | n15294;
  assign n11547 = ~n15293 & n15295;
  assign n11548 = x73 & x108;
  assign n11549 = n11547 & n11548;
  assign n11550 = n11547 | n11548;
  assign n11551 = ~n11549 & n11550;
  assign n15296 = n11468 & n11551;
  assign n15297 = (n11551 & n15249) | (n11551 & n15296) | (n15249 & n15296);
  assign n15298 = n11468 | n11551;
  assign n15299 = n15249 | n15298;
  assign n11554 = ~n15297 & n15299;
  assign n11555 = x72 & x109;
  assign n11556 = n11554 & n11555;
  assign n11557 = n11554 | n11555;
  assign n11558 = ~n11556 & n11557;
  assign n15300 = n11475 & n11558;
  assign n15301 = (n11558 & n15253) | (n11558 & n15300) | (n15253 & n15300);
  assign n15302 = n11475 | n11558;
  assign n15303 = n15253 | n15302;
  assign n11561 = ~n15301 & n15303;
  assign n11562 = x71 & x110;
  assign n11563 = n11561 & n11562;
  assign n11564 = n11561 | n11562;
  assign n11565 = ~n11563 & n11564;
  assign n15304 = n11482 & n11565;
  assign n15305 = (n11565 & n15257) | (n11565 & n15304) | (n15257 & n15304);
  assign n15306 = n11482 | n11565;
  assign n15307 = n15257 | n15306;
  assign n11568 = ~n15305 & n15307;
  assign n11569 = x70 & x111;
  assign n11570 = n11568 & n11569;
  assign n11571 = n11568 | n11569;
  assign n11572 = ~n11570 & n11571;
  assign n15308 = n11489 & n11572;
  assign n15309 = (n11572 & n15261) | (n11572 & n15308) | (n15261 & n15308);
  assign n15310 = n11489 | n11572;
  assign n15311 = n15261 | n15310;
  assign n11575 = ~n15309 & n15311;
  assign n11586 = x79 & x103;
  assign n17504 = n11509 | n17496;
  assign n17505 = (n11426 & n17496) | (n11426 & n17504) | (n17496 & n17504);
  assign n15315 = n11586 & n17505;
  assign n17919 = n11586 & n17495;
  assign n17920 = n11586 & n17494;
  assign n17921 = (n17453 & n17919) | (n17453 & n17920) | (n17919 & n17920);
  assign n17507 = (n11509 & n11586) | (n11509 & n17921) | (n11586 & n17921);
  assign n15317 = (n17486 & n15315) | (n17486 & n17507) | (n15315 & n17507);
  assign n15318 = n11586 | n17505;
  assign n17922 = n11586 | n17495;
  assign n17923 = n11586 | n17494;
  assign n17924 = (n17453 & n17922) | (n17453 & n17923) | (n17922 & n17923);
  assign n17509 = n11509 | n17924;
  assign n15320 = (n17486 & n15318) | (n17486 & n17509) | (n15318 & n17509);
  assign n11589 = ~n15317 & n15320;
  assign n15321 = n11514 & n11589;
  assign n17510 = (n11589 & n15276) | (n11589 & n15321) | (n15276 & n15321);
  assign n17511 = (n11516 & n11589) | (n11516 & n15321) | (n11589 & n15321);
  assign n17512 = (n15229 & n17510) | (n15229 & n17511) | (n17510 & n17511);
  assign n15323 = n11514 | n11589;
  assign n17513 = n15276 | n15323;
  assign n17514 = n11516 | n15323;
  assign n17515 = (n15229 & n17513) | (n15229 & n17514) | (n17513 & n17514);
  assign n11592 = ~n17512 & n17515;
  assign n11593 = x78 & x104;
  assign n11594 = n11592 & n11593;
  assign n11595 = n11592 | n11593;
  assign n11596 = ~n11594 & n11595;
  assign n15325 = n11521 & n11596;
  assign n15326 = (n11596 & n15281) | (n11596 & n15325) | (n15281 & n15325);
  assign n15327 = n11521 | n11596;
  assign n15328 = n15281 | n15327;
  assign n11599 = ~n15326 & n15328;
  assign n11600 = x77 & x105;
  assign n11601 = n11599 & n11600;
  assign n11602 = n11599 | n11600;
  assign n11603 = ~n11601 & n11602;
  assign n15329 = n11528 & n11603;
  assign n15330 = (n11603 & n15285) | (n11603 & n15329) | (n15285 & n15329);
  assign n15331 = n11528 | n11603;
  assign n15332 = n15285 | n15331;
  assign n11606 = ~n15330 & n15332;
  assign n11607 = x76 & x106;
  assign n11608 = n11606 & n11607;
  assign n11609 = n11606 | n11607;
  assign n11610 = ~n11608 & n11609;
  assign n15333 = n11535 & n11610;
  assign n15334 = (n11610 & n15289) | (n11610 & n15333) | (n15289 & n15333);
  assign n15335 = n11535 | n11610;
  assign n15336 = n15289 | n15335;
  assign n11613 = ~n15334 & n15336;
  assign n11614 = x75 & x107;
  assign n11615 = n11613 & n11614;
  assign n11616 = n11613 | n11614;
  assign n11617 = ~n11615 & n11616;
  assign n15337 = n11542 & n11617;
  assign n15338 = (n11617 & n15293) | (n11617 & n15337) | (n15293 & n15337);
  assign n15339 = n11542 | n11617;
  assign n15340 = n15293 | n15339;
  assign n11620 = ~n15338 & n15340;
  assign n11621 = x74 & x108;
  assign n11622 = n11620 & n11621;
  assign n11623 = n11620 | n11621;
  assign n11624 = ~n11622 & n11623;
  assign n15341 = n11549 & n11624;
  assign n15342 = (n11624 & n15297) | (n11624 & n15341) | (n15297 & n15341);
  assign n15343 = n11549 | n11624;
  assign n15344 = n15297 | n15343;
  assign n11627 = ~n15342 & n15344;
  assign n11628 = x73 & x109;
  assign n11629 = n11627 & n11628;
  assign n11630 = n11627 | n11628;
  assign n11631 = ~n11629 & n11630;
  assign n15345 = n11556 & n11631;
  assign n15346 = (n11631 & n15301) | (n11631 & n15345) | (n15301 & n15345);
  assign n15347 = n11556 | n11631;
  assign n15348 = n15301 | n15347;
  assign n11634 = ~n15346 & n15348;
  assign n11635 = x72 & x110;
  assign n11636 = n11634 & n11635;
  assign n11637 = n11634 | n11635;
  assign n11638 = ~n11636 & n11637;
  assign n15349 = n11563 & n11638;
  assign n15350 = (n11638 & n15305) | (n11638 & n15349) | (n15305 & n15349);
  assign n15351 = n11563 | n11638;
  assign n15352 = n15305 | n15351;
  assign n11641 = ~n15350 & n15352;
  assign n11642 = x71 & x111;
  assign n11643 = n11641 & n11642;
  assign n11644 = n11641 | n11642;
  assign n11645 = ~n11643 & n11644;
  assign n15353 = n11570 & n11645;
  assign n15354 = (n11645 & n15309) | (n11645 & n15353) | (n15309 & n15353);
  assign n15355 = n11570 | n11645;
  assign n15356 = n15309 | n15355;
  assign n11648 = ~n15354 & n15356;
  assign n11658 = x79 & x104;
  assign n15358 = n11589 | n15317;
  assign n17516 = (n11514 & n15317) | (n11514 & n15358) | (n15317 & n15358);
  assign n15360 = n11658 & n17516;
  assign n17925 = n11658 & n15315;
  assign n17926 = n11658 & n17507;
  assign n17927 = (n17486 & n17925) | (n17486 & n17926) | (n17925 & n17926);
  assign n17518 = (n11589 & n11658) | (n11589 & n17927) | (n11658 & n17927);
  assign n17519 = (n15276 & n15360) | (n15276 & n17518) | (n15360 & n17518);
  assign n17520 = (n11516 & n15360) | (n11516 & n17518) | (n15360 & n17518);
  assign n17521 = (n15229 & n17519) | (n15229 & n17520) | (n17519 & n17520);
  assign n15363 = n11658 | n17516;
  assign n17928 = n11658 | n15315;
  assign n17929 = n11658 | n17507;
  assign n17930 = (n17486 & n17928) | (n17486 & n17929) | (n17928 & n17929);
  assign n17523 = n11589 | n17930;
  assign n17524 = (n15276 & n15363) | (n15276 & n17523) | (n15363 & n17523);
  assign n17525 = (n11516 & n15363) | (n11516 & n17523) | (n15363 & n17523);
  assign n17526 = (n15229 & n17524) | (n15229 & n17525) | (n17524 & n17525);
  assign n11661 = ~n17521 & n17526;
  assign n15366 = n11594 & n11661;
  assign n17527 = (n11661 & n15325) | (n11661 & n15366) | (n15325 & n15366);
  assign n17528 = (n11596 & n11661) | (n11596 & n15366) | (n11661 & n15366);
  assign n17529 = (n15281 & n17527) | (n15281 & n17528) | (n17527 & n17528);
  assign n15368 = n11594 | n11661;
  assign n17530 = n15325 | n15368;
  assign n17531 = n11596 | n15368;
  assign n17532 = (n15281 & n17530) | (n15281 & n17531) | (n17530 & n17531);
  assign n11664 = ~n17529 & n17532;
  assign n11665 = x78 & x105;
  assign n11666 = n11664 & n11665;
  assign n11667 = n11664 | n11665;
  assign n11668 = ~n11666 & n11667;
  assign n15370 = n11601 & n11668;
  assign n15371 = (n11668 & n15330) | (n11668 & n15370) | (n15330 & n15370);
  assign n15372 = n11601 | n11668;
  assign n15373 = n15330 | n15372;
  assign n11671 = ~n15371 & n15373;
  assign n11672 = x77 & x106;
  assign n11673 = n11671 & n11672;
  assign n11674 = n11671 | n11672;
  assign n11675 = ~n11673 & n11674;
  assign n15374 = n11608 & n11675;
  assign n15375 = (n11675 & n15334) | (n11675 & n15374) | (n15334 & n15374);
  assign n15376 = n11608 | n11675;
  assign n15377 = n15334 | n15376;
  assign n11678 = ~n15375 & n15377;
  assign n11679 = x76 & x107;
  assign n11680 = n11678 & n11679;
  assign n11681 = n11678 | n11679;
  assign n11682 = ~n11680 & n11681;
  assign n15378 = n11615 & n11682;
  assign n15379 = (n11682 & n15338) | (n11682 & n15378) | (n15338 & n15378);
  assign n15380 = n11615 | n11682;
  assign n15381 = n15338 | n15380;
  assign n11685 = ~n15379 & n15381;
  assign n11686 = x75 & x108;
  assign n11687 = n11685 & n11686;
  assign n11688 = n11685 | n11686;
  assign n11689 = ~n11687 & n11688;
  assign n15382 = n11622 & n11689;
  assign n15383 = (n11689 & n15342) | (n11689 & n15382) | (n15342 & n15382);
  assign n15384 = n11622 | n11689;
  assign n15385 = n15342 | n15384;
  assign n11692 = ~n15383 & n15385;
  assign n11693 = x74 & x109;
  assign n11694 = n11692 & n11693;
  assign n11695 = n11692 | n11693;
  assign n11696 = ~n11694 & n11695;
  assign n15386 = n11629 & n11696;
  assign n15387 = (n11696 & n15346) | (n11696 & n15386) | (n15346 & n15386);
  assign n15388 = n11629 | n11696;
  assign n15389 = n15346 | n15388;
  assign n11699 = ~n15387 & n15389;
  assign n11700 = x73 & x110;
  assign n11701 = n11699 & n11700;
  assign n11702 = n11699 | n11700;
  assign n11703 = ~n11701 & n11702;
  assign n15390 = n11636 & n11703;
  assign n15391 = (n11703 & n15350) | (n11703 & n15390) | (n15350 & n15390);
  assign n15392 = n11636 | n11703;
  assign n15393 = n15350 | n15392;
  assign n11706 = ~n15391 & n15393;
  assign n11707 = x72 & x111;
  assign n11708 = n11706 & n11707;
  assign n11709 = n11706 | n11707;
  assign n11710 = ~n11708 & n11709;
  assign n15394 = n11643 & n11710;
  assign n15395 = (n11710 & n15354) | (n11710 & n15394) | (n15354 & n15394);
  assign n15396 = n11643 | n11710;
  assign n15397 = n15354 | n15396;
  assign n11713 = ~n15395 & n15397;
  assign n11722 = x79 & x105;
  assign n17533 = n11661 | n17521;
  assign n17534 = (n11594 & n17521) | (n11594 & n17533) | (n17521 & n17533);
  assign n15401 = n11722 & n17534;
  assign n17535 = n11722 & n17521;
  assign n17536 = (n11661 & n11722) | (n11661 & n17535) | (n11722 & n17535);
  assign n17537 = (n15325 & n15401) | (n15325 & n17536) | (n15401 & n17536);
  assign n17538 = (n11596 & n15401) | (n11596 & n17536) | (n15401 & n17536);
  assign n17539 = (n15281 & n17537) | (n15281 & n17538) | (n17537 & n17538);
  assign n15404 = n11722 | n17534;
  assign n17540 = n11722 | n17521;
  assign n17541 = n11661 | n17540;
  assign n17542 = (n15325 & n15404) | (n15325 & n17541) | (n15404 & n17541);
  assign n17543 = (n11596 & n15404) | (n11596 & n17541) | (n15404 & n17541);
  assign n17544 = (n15281 & n17542) | (n15281 & n17543) | (n17542 & n17543);
  assign n11725 = ~n17539 & n17544;
  assign n15407 = n11666 & n11725;
  assign n17545 = (n11725 & n15370) | (n11725 & n15407) | (n15370 & n15407);
  assign n17546 = (n11668 & n11725) | (n11668 & n15407) | (n11725 & n15407);
  assign n17547 = (n15330 & n17545) | (n15330 & n17546) | (n17545 & n17546);
  assign n15409 = n11666 | n11725;
  assign n17548 = n15370 | n15409;
  assign n17549 = n11668 | n15409;
  assign n17550 = (n15330 & n17548) | (n15330 & n17549) | (n17548 & n17549);
  assign n11728 = ~n17547 & n17550;
  assign n11729 = x78 & x106;
  assign n11730 = n11728 & n11729;
  assign n11731 = n11728 | n11729;
  assign n11732 = ~n11730 & n11731;
  assign n15411 = n11673 & n11732;
  assign n15412 = (n11732 & n15375) | (n11732 & n15411) | (n15375 & n15411);
  assign n15413 = n11673 | n11732;
  assign n15414 = n15375 | n15413;
  assign n11735 = ~n15412 & n15414;
  assign n11736 = x77 & x107;
  assign n11737 = n11735 & n11736;
  assign n11738 = n11735 | n11736;
  assign n11739 = ~n11737 & n11738;
  assign n15415 = n11680 & n11739;
  assign n15416 = (n11739 & n15379) | (n11739 & n15415) | (n15379 & n15415);
  assign n15417 = n11680 | n11739;
  assign n15418 = n15379 | n15417;
  assign n11742 = ~n15416 & n15418;
  assign n11743 = x76 & x108;
  assign n11744 = n11742 & n11743;
  assign n11745 = n11742 | n11743;
  assign n11746 = ~n11744 & n11745;
  assign n15419 = n11687 & n11746;
  assign n15420 = (n11746 & n15383) | (n11746 & n15419) | (n15383 & n15419);
  assign n15421 = n11687 | n11746;
  assign n15422 = n15383 | n15421;
  assign n11749 = ~n15420 & n15422;
  assign n11750 = x75 & x109;
  assign n11751 = n11749 & n11750;
  assign n11752 = n11749 | n11750;
  assign n11753 = ~n11751 & n11752;
  assign n15423 = n11694 & n11753;
  assign n15424 = (n11753 & n15387) | (n11753 & n15423) | (n15387 & n15423);
  assign n15425 = n11694 | n11753;
  assign n15426 = n15387 | n15425;
  assign n11756 = ~n15424 & n15426;
  assign n11757 = x74 & x110;
  assign n11758 = n11756 & n11757;
  assign n11759 = n11756 | n11757;
  assign n11760 = ~n11758 & n11759;
  assign n15427 = n11701 & n11760;
  assign n15428 = (n11760 & n15391) | (n11760 & n15427) | (n15391 & n15427);
  assign n15429 = n11701 | n11760;
  assign n15430 = n15391 | n15429;
  assign n11763 = ~n15428 & n15430;
  assign n11764 = x73 & x111;
  assign n11765 = n11763 & n11764;
  assign n11766 = n11763 | n11764;
  assign n11767 = ~n11765 & n11766;
  assign n15431 = n11708 & n11767;
  assign n15432 = (n11767 & n15395) | (n11767 & n15431) | (n15395 & n15431);
  assign n15433 = n11708 | n11767;
  assign n15434 = n15395 | n15433;
  assign n11770 = ~n15432 & n15434;
  assign n11778 = x79 & x106;
  assign n17551 = n11725 | n17539;
  assign n17552 = (n11666 & n17539) | (n11666 & n17551) | (n17539 & n17551);
  assign n15438 = n11778 & n17552;
  assign n17553 = n11778 & n17539;
  assign n17554 = (n11725 & n11778) | (n11725 & n17553) | (n11778 & n17553);
  assign n17555 = (n15370 & n15438) | (n15370 & n17554) | (n15438 & n17554);
  assign n17556 = (n11668 & n15438) | (n11668 & n17554) | (n15438 & n17554);
  assign n17557 = (n15330 & n17555) | (n15330 & n17556) | (n17555 & n17556);
  assign n15441 = n11778 | n17552;
  assign n17558 = n11778 | n17539;
  assign n17559 = n11725 | n17558;
  assign n17560 = (n15370 & n15441) | (n15370 & n17559) | (n15441 & n17559);
  assign n17561 = (n11668 & n15441) | (n11668 & n17559) | (n15441 & n17559);
  assign n17562 = (n15330 & n17560) | (n15330 & n17561) | (n17560 & n17561);
  assign n11781 = ~n17557 & n17562;
  assign n15444 = n11730 & n11781;
  assign n17563 = (n11781 & n15411) | (n11781 & n15444) | (n15411 & n15444);
  assign n17564 = (n11732 & n11781) | (n11732 & n15444) | (n11781 & n15444);
  assign n17565 = (n15375 & n17563) | (n15375 & n17564) | (n17563 & n17564);
  assign n15446 = n11730 | n11781;
  assign n17566 = n15411 | n15446;
  assign n17567 = n11732 | n15446;
  assign n17568 = (n15375 & n17566) | (n15375 & n17567) | (n17566 & n17567);
  assign n11784 = ~n17565 & n17568;
  assign n11785 = x78 & x107;
  assign n11786 = n11784 & n11785;
  assign n11787 = n11784 | n11785;
  assign n11788 = ~n11786 & n11787;
  assign n15448 = n11737 & n11788;
  assign n15449 = (n11788 & n15416) | (n11788 & n15448) | (n15416 & n15448);
  assign n15450 = n11737 | n11788;
  assign n15451 = n15416 | n15450;
  assign n11791 = ~n15449 & n15451;
  assign n11792 = x77 & x108;
  assign n11793 = n11791 & n11792;
  assign n11794 = n11791 | n11792;
  assign n11795 = ~n11793 & n11794;
  assign n15452 = n11744 & n11795;
  assign n15453 = (n11795 & n15420) | (n11795 & n15452) | (n15420 & n15452);
  assign n15454 = n11744 | n11795;
  assign n15455 = n15420 | n15454;
  assign n11798 = ~n15453 & n15455;
  assign n11799 = x76 & x109;
  assign n11800 = n11798 & n11799;
  assign n11801 = n11798 | n11799;
  assign n11802 = ~n11800 & n11801;
  assign n15456 = n11751 & n11802;
  assign n15457 = (n11802 & n15424) | (n11802 & n15456) | (n15424 & n15456);
  assign n15458 = n11751 | n11802;
  assign n15459 = n15424 | n15458;
  assign n11805 = ~n15457 & n15459;
  assign n11806 = x75 & x110;
  assign n11807 = n11805 & n11806;
  assign n11808 = n11805 | n11806;
  assign n11809 = ~n11807 & n11808;
  assign n15460 = n11758 & n11809;
  assign n15461 = (n11809 & n15428) | (n11809 & n15460) | (n15428 & n15460);
  assign n15462 = n11758 | n11809;
  assign n15463 = n15428 | n15462;
  assign n11812 = ~n15461 & n15463;
  assign n11813 = x74 & x111;
  assign n11814 = n11812 & n11813;
  assign n11815 = n11812 | n11813;
  assign n11816 = ~n11814 & n11815;
  assign n15464 = n11765 & n11816;
  assign n15465 = (n11816 & n15432) | (n11816 & n15464) | (n15432 & n15464);
  assign n15466 = n11765 | n11816;
  assign n15467 = n15432 | n15466;
  assign n11819 = ~n15465 & n15467;
  assign n11826 = x79 & x107;
  assign n17569 = n11781 | n17557;
  assign n17570 = (n11730 & n17557) | (n11730 & n17569) | (n17557 & n17569);
  assign n15471 = n11826 & n17570;
  assign n17571 = n11826 & n17557;
  assign n17572 = (n11781 & n11826) | (n11781 & n17571) | (n11826 & n17571);
  assign n17573 = (n15411 & n15471) | (n15411 & n17572) | (n15471 & n17572);
  assign n17574 = (n11732 & n15471) | (n11732 & n17572) | (n15471 & n17572);
  assign n17575 = (n15375 & n17573) | (n15375 & n17574) | (n17573 & n17574);
  assign n15474 = n11826 | n17570;
  assign n17576 = n11826 | n17557;
  assign n17577 = n11781 | n17576;
  assign n17578 = (n15411 & n15474) | (n15411 & n17577) | (n15474 & n17577);
  assign n17579 = (n11732 & n15474) | (n11732 & n17577) | (n15474 & n17577);
  assign n17580 = (n15375 & n17578) | (n15375 & n17579) | (n17578 & n17579);
  assign n11829 = ~n17575 & n17580;
  assign n15477 = n11786 & n11829;
  assign n17581 = (n11829 & n15448) | (n11829 & n15477) | (n15448 & n15477);
  assign n17582 = (n11788 & n11829) | (n11788 & n15477) | (n11829 & n15477);
  assign n17583 = (n15416 & n17581) | (n15416 & n17582) | (n17581 & n17582);
  assign n15479 = n11786 | n11829;
  assign n17584 = n15448 | n15479;
  assign n17585 = n11788 | n15479;
  assign n17586 = (n15416 & n17584) | (n15416 & n17585) | (n17584 & n17585);
  assign n11832 = ~n17583 & n17586;
  assign n11833 = x78 & x108;
  assign n11834 = n11832 & n11833;
  assign n11835 = n11832 | n11833;
  assign n11836 = ~n11834 & n11835;
  assign n15481 = n11793 & n11836;
  assign n15482 = (n11836 & n15453) | (n11836 & n15481) | (n15453 & n15481);
  assign n15483 = n11793 | n11836;
  assign n15484 = n15453 | n15483;
  assign n11839 = ~n15482 & n15484;
  assign n11840 = x77 & x109;
  assign n11841 = n11839 & n11840;
  assign n11842 = n11839 | n11840;
  assign n11843 = ~n11841 & n11842;
  assign n15485 = n11800 & n11843;
  assign n15486 = (n11843 & n15457) | (n11843 & n15485) | (n15457 & n15485);
  assign n15487 = n11800 | n11843;
  assign n15488 = n15457 | n15487;
  assign n11846 = ~n15486 & n15488;
  assign n11847 = x76 & x110;
  assign n11848 = n11846 & n11847;
  assign n11849 = n11846 | n11847;
  assign n11850 = ~n11848 & n11849;
  assign n15489 = n11807 & n11850;
  assign n15490 = (n11850 & n15461) | (n11850 & n15489) | (n15461 & n15489);
  assign n15491 = n11807 | n11850;
  assign n15492 = n15461 | n15491;
  assign n11853 = ~n15490 & n15492;
  assign n11854 = x75 & x111;
  assign n11855 = n11853 & n11854;
  assign n11856 = n11853 | n11854;
  assign n11857 = ~n11855 & n11856;
  assign n15493 = n11814 & n11857;
  assign n15494 = (n11857 & n15465) | (n11857 & n15493) | (n15465 & n15493);
  assign n15495 = n11814 | n11857;
  assign n15496 = n15465 | n15495;
  assign n11860 = ~n15494 & n15496;
  assign n11866 = x79 & x108;
  assign n17587 = n11829 | n17575;
  assign n17588 = (n11786 & n17575) | (n11786 & n17587) | (n17575 & n17587);
  assign n15500 = n11866 & n17588;
  assign n17589 = n11866 & n17575;
  assign n17590 = (n11829 & n11866) | (n11829 & n17589) | (n11866 & n17589);
  assign n17591 = (n15448 & n15500) | (n15448 & n17590) | (n15500 & n17590);
  assign n17592 = (n11788 & n15500) | (n11788 & n17590) | (n15500 & n17590);
  assign n17593 = (n15416 & n17591) | (n15416 & n17592) | (n17591 & n17592);
  assign n15503 = n11866 | n17588;
  assign n17594 = n11866 | n17575;
  assign n17595 = n11829 | n17594;
  assign n17596 = (n15448 & n15503) | (n15448 & n17595) | (n15503 & n17595);
  assign n17597 = (n11788 & n15503) | (n11788 & n17595) | (n15503 & n17595);
  assign n17598 = (n15416 & n17596) | (n15416 & n17597) | (n17596 & n17597);
  assign n11869 = ~n17593 & n17598;
  assign n15506 = n11834 & n11869;
  assign n17599 = (n11869 & n15481) | (n11869 & n15506) | (n15481 & n15506);
  assign n17600 = (n11836 & n11869) | (n11836 & n15506) | (n11869 & n15506);
  assign n17601 = (n15453 & n17599) | (n15453 & n17600) | (n17599 & n17600);
  assign n15508 = n11834 | n11869;
  assign n17602 = n15481 | n15508;
  assign n17603 = n11836 | n15508;
  assign n17604 = (n15453 & n17602) | (n15453 & n17603) | (n17602 & n17603);
  assign n11872 = ~n17601 & n17604;
  assign n11873 = x78 & x109;
  assign n11874 = n11872 & n11873;
  assign n11875 = n11872 | n11873;
  assign n11876 = ~n11874 & n11875;
  assign n15510 = n11841 & n11876;
  assign n15511 = (n11876 & n15486) | (n11876 & n15510) | (n15486 & n15510);
  assign n15512 = n11841 | n11876;
  assign n15513 = n15486 | n15512;
  assign n11879 = ~n15511 & n15513;
  assign n11880 = x77 & x110;
  assign n11881 = n11879 & n11880;
  assign n11882 = n11879 | n11880;
  assign n11883 = ~n11881 & n11882;
  assign n15514 = n11848 & n11883;
  assign n15515 = (n11883 & n15490) | (n11883 & n15514) | (n15490 & n15514);
  assign n15516 = n11848 | n11883;
  assign n15517 = n15490 | n15516;
  assign n11886 = ~n15515 & n15517;
  assign n11887 = x76 & x111;
  assign n11888 = n11886 & n11887;
  assign n11889 = n11886 | n11887;
  assign n11890 = ~n11888 & n11889;
  assign n15518 = n11855 & n11890;
  assign n15519 = (n11890 & n15494) | (n11890 & n15518) | (n15494 & n15518);
  assign n15520 = n11855 | n11890;
  assign n15521 = n15494 | n15520;
  assign n11893 = ~n15519 & n15521;
  assign n11898 = x79 & x109;
  assign n17605 = n11869 | n17593;
  assign n17606 = (n11834 & n17593) | (n11834 & n17605) | (n17593 & n17605);
  assign n15525 = n11898 & n17606;
  assign n17607 = n11898 & n17593;
  assign n17608 = (n11869 & n11898) | (n11869 & n17607) | (n11898 & n17607);
  assign n17609 = (n15481 & n15525) | (n15481 & n17608) | (n15525 & n17608);
  assign n17610 = (n11836 & n15525) | (n11836 & n17608) | (n15525 & n17608);
  assign n17611 = (n15453 & n17609) | (n15453 & n17610) | (n17609 & n17610);
  assign n15528 = n11898 | n17606;
  assign n17612 = n11898 | n17593;
  assign n17613 = n11869 | n17612;
  assign n17614 = (n15481 & n15528) | (n15481 & n17613) | (n15528 & n17613);
  assign n17615 = (n11836 & n15528) | (n11836 & n17613) | (n15528 & n17613);
  assign n17616 = (n15453 & n17614) | (n15453 & n17615) | (n17614 & n17615);
  assign n11901 = ~n17611 & n17616;
  assign n15531 = n11874 & n11901;
  assign n17617 = (n11901 & n15510) | (n11901 & n15531) | (n15510 & n15531);
  assign n17618 = (n11876 & n11901) | (n11876 & n15531) | (n11901 & n15531);
  assign n17619 = (n15486 & n17617) | (n15486 & n17618) | (n17617 & n17618);
  assign n15533 = n11874 | n11901;
  assign n17620 = n15510 | n15533;
  assign n17621 = n11876 | n15533;
  assign n17622 = (n15486 & n17620) | (n15486 & n17621) | (n17620 & n17621);
  assign n11904 = ~n17619 & n17622;
  assign n11905 = x78 & x110;
  assign n11906 = n11904 & n11905;
  assign n11907 = n11904 | n11905;
  assign n11908 = ~n11906 & n11907;
  assign n15535 = n11881 & n11908;
  assign n15536 = (n11908 & n15515) | (n11908 & n15535) | (n15515 & n15535);
  assign n15537 = n11881 | n11908;
  assign n15538 = n15515 | n15537;
  assign n11911 = ~n15536 & n15538;
  assign n11912 = x77 & x111;
  assign n11913 = n11911 & n11912;
  assign n11914 = n11911 | n11912;
  assign n11915 = ~n11913 & n11914;
  assign n15539 = n11888 & n11915;
  assign n15540 = (n11915 & n15519) | (n11915 & n15539) | (n15519 & n15539);
  assign n15541 = n11888 | n11915;
  assign n15542 = n15519 | n15541;
  assign n11918 = ~n15540 & n15542;
  assign n11922 = x79 & x110;
  assign n17623 = n11901 | n17611;
  assign n17624 = (n11874 & n17611) | (n11874 & n17623) | (n17611 & n17623);
  assign n15546 = n11922 & n17624;
  assign n17625 = n11922 & n17611;
  assign n17626 = (n11901 & n11922) | (n11901 & n17625) | (n11922 & n17625);
  assign n17627 = (n15510 & n15546) | (n15510 & n17626) | (n15546 & n17626);
  assign n17628 = (n11876 & n15546) | (n11876 & n17626) | (n15546 & n17626);
  assign n17629 = (n15486 & n17627) | (n15486 & n17628) | (n17627 & n17628);
  assign n15549 = n11922 | n17624;
  assign n17630 = n11922 | n17611;
  assign n17631 = n11901 | n17630;
  assign n17632 = (n15510 & n15549) | (n15510 & n17631) | (n15549 & n17631);
  assign n17633 = (n11876 & n15549) | (n11876 & n17631) | (n15549 & n17631);
  assign n17634 = (n15486 & n17632) | (n15486 & n17633) | (n17632 & n17633);
  assign n11925 = ~n17629 & n17634;
  assign n15552 = n11906 & n11925;
  assign n17635 = (n11925 & n15535) | (n11925 & n15552) | (n15535 & n15552);
  assign n17636 = (n11908 & n11925) | (n11908 & n15552) | (n11925 & n15552);
  assign n17637 = (n15515 & n17635) | (n15515 & n17636) | (n17635 & n17636);
  assign n15554 = n11906 | n11925;
  assign n17638 = n15535 | n15554;
  assign n17639 = n11908 | n15554;
  assign n17640 = (n15515 & n17638) | (n15515 & n17639) | (n17638 & n17639);
  assign n11928 = ~n17637 & n17640;
  assign n11929 = x78 & x111;
  assign n11930 = n11928 & n11929;
  assign n11931 = n11928 | n11929;
  assign n11932 = ~n11930 & n11931;
  assign n15556 = n11913 & n11932;
  assign n15557 = (n11932 & n15540) | (n11932 & n15556) | (n15540 & n15556);
  assign n15558 = n11913 | n11932;
  assign n15559 = n15540 | n15558;
  assign n11935 = ~n15557 & n15559;
  assign n11938 = x79 & x111;
  assign n17641 = n11925 | n17629;
  assign n17642 = (n11906 & n17629) | (n11906 & n17641) | (n17629 & n17641);
  assign n15563 = n11938 & n17642;
  assign n17643 = n11938 & n17629;
  assign n17644 = (n11925 & n11938) | (n11925 & n17643) | (n11938 & n17643);
  assign n17645 = (n15535 & n15563) | (n15535 & n17644) | (n15563 & n17644);
  assign n17646 = (n11908 & n15563) | (n11908 & n17644) | (n15563 & n17644);
  assign n17647 = (n15515 & n17645) | (n15515 & n17646) | (n17645 & n17646);
  assign n15566 = n11938 | n17642;
  assign n17648 = n11938 | n17629;
  assign n17649 = n11925 | n17648;
  assign n17650 = (n15535 & n15566) | (n15535 & n17649) | (n15566 & n17649);
  assign n17651 = (n11908 & n15566) | (n11908 & n17649) | (n15566 & n17649);
  assign n17652 = (n15515 & n17650) | (n15515 & n17651) | (n17650 & n17651);
  assign n11941 = ~n17647 & n17652;
  assign n15569 = n11930 & n11941;
  assign n17653 = (n11941 & n15556) | (n11941 & n15569) | (n15556 & n15569);
  assign n17654 = (n11932 & n11941) | (n11932 & n15569) | (n11941 & n15569);
  assign n17655 = (n15540 & n17653) | (n15540 & n17654) | (n17653 & n17654);
  assign n15571 = n11930 | n11941;
  assign n17656 = n15556 | n15571;
  assign n17657 = n11932 | n15571;
  assign n17658 = (n15540 & n17656) | (n15540 & n17657) | (n17656 & n17657);
  assign n11944 = ~n17655 & n17658;
  assign n15574 = n11941 | n17647;
  assign n17659 = n11941 | n17647;
  assign n17660 = (n11930 & n17647) | (n11930 & n17659) | (n17647 & n17659);
  assign n17661 = (n15556 & n15574) | (n15556 & n17660) | (n15574 & n17660);
  assign n17662 = (n11932 & n15574) | (n11932 & n17660) | (n15574 & n17660);
  assign n17663 = (n15540 & n17661) | (n15540 & n17662) | (n17661 & n17662);
  assign y0 = n17;
  assign y1 = n22;
  assign y2 = n34;
  assign y3 = n54;
  assign y4 = n82;
  assign y5 = n118;
  assign y6 = n162;
  assign y7 = n214;
  assign y8 = n266;
  assign y9 = n314;
  assign y10 = n355;
  assign y11 = n388;
  assign y12 = n413;
  assign y13 = n430;
  assign y14 = n439;
  assign y15 = n723;
  assign y16 = n799;
  assign y17 = n804;
  assign y18 = n816;
  assign y19 = n836;
  assign y20 = n864;
  assign y21 = n900;
  assign y22 = n944;
  assign y23 = n996;
  assign y24 = n1056;
  assign y25 = n1124;
  assign y26 = n1200;
  assign y27 = n1284;
  assign y28 = n1376;
  assign y29 = n1476;
  assign y30 = n1584;
  assign y31 = n1700;
  assign y32 = n1816;
  assign y33 = n1928;
  assign y34 = n2033;
  assign y35 = n2130;
  assign y36 = n2219;
  assign y37 = n2300;
  assign y38 = n2373;
  assign y39 = n2438;
  assign y40 = n2495;
  assign y41 = n2544;
  assign y42 = n2585;
  assign y43 = n2618;
  assign y44 = n2643;
  assign y45 = n2660;
  assign y46 = n2669;
  assign y47 = n3894;
  assign y48 = n4106;
  assign y49 = n4111;
  assign y50 = n4123;
  assign y51 = n4143;
  assign y52 = n4171;
  assign y53 = n4207;
  assign y54 = n4251;
  assign y55 = n4303;
  assign y56 = n4363;
  assign y57 = n4431;
  assign y58 = n4507;
  assign y59 = n4591;
  assign y60 = n4683;
  assign y61 = n4783;
  assign y62 = n4891;
  assign y63 = n5007;
  assign y64 = n5131;
  assign y65 = n5263;
  assign y66 = n5403;
  assign y67 = n5551;
  assign y68 = n5707;
  assign y69 = n5871;
  assign y70 = n6043;
  assign y71 = n6223;
  assign y72 = n6411;
  assign y73 = n6607;
  assign y74 = n6811;
  assign y75 = n7023;
  assign y76 = n7243;
  assign y77 = n7471;
  assign y78 = n7707;
  assign y79 = n7951;
  assign y80 = n8195;
  assign y81 = n8435;
  assign y82 = n8668;
  assign y83 = n8893;
  assign y84 = n9110;
  assign y85 = n9319;
  assign y86 = n9520;
  assign y87 = n9713;
  assign y88 = n9898;
  assign y89 = n10075;
  assign y90 = n10244;
  assign y91 = n10405;
  assign y92 = n10558;
  assign y93 = n10703;
  assign y94 = n10840;
  assign y95 = n10969;
  assign y96 = n11090;
  assign y97 = n11203;
  assign y98 = n11308;
  assign y99 = n11405;
  assign y100 = n11494;
  assign y101 = n11575;
  assign y102 = n11648;
  assign y103 = n11713;
  assign y104 = n11770;
  assign y105 = n11819;
  assign y106 = n11860;
  assign y107 = n11893;
  assign y108 = n11918;
  assign y109 = n11935;
  assign y110 = n11944;
  assign y111 = n17663;
endmodule

