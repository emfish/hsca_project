module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159, y160, y161, y162, y163, y164, y165, y166, y167, y168, y169, y170, y171, y172, y173, y174, y175);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159, y160, y161, y162, y163, y164, y165, y166, y167, y168, y169, y170, y171, y172, y173, y174, y175;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934;
  assign n17 = x0 & x8;
  assign n18 = x1 & x8;
  assign n19 = x0 & x9;
  assign n20 = n18 & n19;
  assign n21 = n18 | n19;
  assign n22 = ~n20 & n21;
  assign n23 = x2 & x8;
  assign n24 = x1 & x9;
  assign n25 = n23 & n24;
  assign n26 = n23 | n24;
  assign n27 = ~n25 & n26;
  assign n28 = n20 & n27;
  assign n29 = n20 | n27;
  assign n30 = ~n28 & n29;
  assign n31 = x0 & x10;
  assign n32 = n30 & n31;
  assign n33 = n30 | n31;
  assign n34 = ~n32 & n33;
  assign n441 = n20 | n25;
  assign n442 = (n25 & n27) | (n25 & n441) | (n27 & n441);
  assign n36 = x3 & x8;
  assign n37 = x2 & x9;
  assign n38 = n36 & n37;
  assign n39 = n36 | n37;
  assign n40 = ~n38 & n39;
  assign n41 = n442 & n40;
  assign n42 = n442 | n40;
  assign n43 = ~n41 & n42;
  assign n44 = x1 & x10;
  assign n45 = n43 & n44;
  assign n46 = n43 | n44;
  assign n47 = ~n45 & n46;
  assign n48 = n32 & n47;
  assign n49 = n32 | n47;
  assign n50 = ~n48 & n49;
  assign n51 = x0 & x11;
  assign n52 = n50 & n51;
  assign n53 = n50 | n51;
  assign n54 = ~n52 & n53;
  assign n443 = n32 | n45;
  assign n444 = (n45 & n47) | (n45 & n443) | (n47 & n443);
  assign n445 = n38 | n40;
  assign n446 = (n38 & n442) | (n38 & n445) | (n442 & n445);
  assign n57 = x4 & x8;
  assign n58 = x3 & x9;
  assign n59 = n57 & n58;
  assign n60 = n57 | n58;
  assign n61 = ~n59 & n60;
  assign n62 = n446 & n61;
  assign n63 = n446 | n61;
  assign n64 = ~n62 & n63;
  assign n65 = x2 & x10;
  assign n66 = n64 & n65;
  assign n67 = n64 | n65;
  assign n68 = ~n66 & n67;
  assign n69 = n444 & n68;
  assign n70 = n444 | n68;
  assign n71 = ~n69 & n70;
  assign n72 = x1 & x11;
  assign n73 = n71 & n72;
  assign n74 = n71 | n72;
  assign n75 = ~n73 & n74;
  assign n76 = n52 & n75;
  assign n77 = n52 | n75;
  assign n78 = ~n76 & n77;
  assign n79 = x0 & x12;
  assign n80 = n78 & n79;
  assign n81 = n78 | n79;
  assign n82 = ~n80 & n81;
  assign n447 = n52 | n73;
  assign n448 = (n73 & n75) | (n73 & n447) | (n75 & n447);
  assign n86 = x5 & x8;
  assign n87 = x4 & x9;
  assign n88 = n86 & n87;
  assign n89 = n86 | n87;
  assign n90 = ~n88 & n89;
  assign n449 = n59 | n61;
  assign n451 = n90 & n449;
  assign n452 = n59 & n90;
  assign n453 = (n446 & n451) | (n446 & n452) | (n451 & n452);
  assign n454 = n90 | n449;
  assign n455 = n59 | n90;
  assign n456 = (n446 & n454) | (n446 & n455) | (n454 & n455);
  assign n93 = ~n453 & n456;
  assign n94 = x3 & x10;
  assign n95 = n93 & n94;
  assign n96 = n93 | n94;
  assign n97 = ~n95 & n96;
  assign n457 = n66 & n97;
  assign n458 = (n69 & n97) | (n69 & n457) | (n97 & n457);
  assign n459 = n66 | n97;
  assign n460 = n69 | n459;
  assign n100 = ~n458 & n460;
  assign n101 = x2 & x11;
  assign n102 = n100 & n101;
  assign n103 = n100 | n101;
  assign n104 = ~n102 & n103;
  assign n105 = n448 & n104;
  assign n106 = n448 | n104;
  assign n107 = ~n105 & n106;
  assign n108 = x1 & x12;
  assign n109 = n107 & n108;
  assign n110 = n107 | n108;
  assign n111 = ~n109 & n110;
  assign n112 = n80 & n111;
  assign n113 = n80 | n111;
  assign n114 = ~n112 & n113;
  assign n115 = x0 & x13;
  assign n116 = n114 & n115;
  assign n117 = n114 | n115;
  assign n118 = ~n116 & n117;
  assign n461 = n80 | n109;
  assign n462 = (n109 & n111) | (n109 & n461) | (n111 & n461);
  assign n120 = n102 | n105;
  assign n123 = x6 & x8;
  assign n124 = x5 & x9;
  assign n125 = n123 & n124;
  assign n126 = n123 | n124;
  assign n127 = ~n125 & n126;
  assign n463 = n88 & n127;
  assign n464 = (n127 & n453) | (n127 & n463) | (n453 & n463);
  assign n465 = n88 | n127;
  assign n466 = n453 | n465;
  assign n130 = ~n464 & n466;
  assign n131 = x4 & x10;
  assign n132 = n130 & n131;
  assign n133 = n130 | n131;
  assign n134 = ~n132 & n133;
  assign n467 = n95 & n134;
  assign n468 = (n134 & n458) | (n134 & n467) | (n458 & n467);
  assign n469 = n95 | n134;
  assign n470 = n458 | n469;
  assign n137 = ~n468 & n470;
  assign n138 = x3 & x11;
  assign n139 = n137 & n138;
  assign n140 = n137 | n138;
  assign n141 = ~n139 & n140;
  assign n142 = n120 & n141;
  assign n143 = n120 | n141;
  assign n144 = ~n142 & n143;
  assign n145 = x2 & x12;
  assign n146 = n144 & n145;
  assign n147 = n144 | n145;
  assign n148 = ~n146 & n147;
  assign n149 = n462 & n148;
  assign n150 = n462 | n148;
  assign n151 = ~n149 & n150;
  assign n152 = x1 & x13;
  assign n153 = n151 & n152;
  assign n154 = n151 | n152;
  assign n155 = ~n153 & n154;
  assign n156 = n116 & n155;
  assign n157 = n116 | n155;
  assign n158 = ~n156 & n157;
  assign n159 = x0 & x14;
  assign n160 = n158 & n159;
  assign n161 = n158 | n159;
  assign n162 = ~n160 & n161;
  assign n724 = n115 | n152;
  assign n725 = (n114 & n152) | (n114 & n724) | (n152 & n724);
  assign n598 = (n116 & n151) | (n116 & n725) | (n151 & n725);
  assign n472 = (n153 & n155) | (n153 & n598) | (n155 & n598);
  assign n473 = n146 | n462;
  assign n474 = (n146 & n148) | (n146 & n473) | (n148 & n473);
  assign n475 = n139 | n141;
  assign n476 = (n120 & n139) | (n120 & n475) | (n139 & n475);
  assign n168 = x7 & x8;
  assign n169 = x6 & x9;
  assign n170 = n168 & n169;
  assign n171 = n168 | n169;
  assign n172 = ~n170 & n171;
  assign n599 = n88 | n125;
  assign n600 = (n125 & n127) | (n125 & n599) | (n127 & n599);
  assign n480 = n172 & n600;
  assign n478 = n125 | n127;
  assign n481 = n172 & n478;
  assign n482 = (n453 & n480) | (n453 & n481) | (n480 & n481);
  assign n483 = n172 | n600;
  assign n484 = n172 | n478;
  assign n485 = (n453 & n483) | (n453 & n484) | (n483 & n484);
  assign n175 = ~n482 & n485;
  assign n176 = x5 & x10;
  assign n177 = n175 & n176;
  assign n178 = n175 | n176;
  assign n179 = ~n177 & n178;
  assign n486 = n132 & n179;
  assign n487 = (n179 & n468) | (n179 & n486) | (n468 & n486);
  assign n488 = n132 | n179;
  assign n489 = n468 | n488;
  assign n182 = ~n487 & n489;
  assign n183 = x4 & x11;
  assign n184 = n182 & n183;
  assign n185 = n182 | n183;
  assign n186 = ~n184 & n185;
  assign n187 = n476 & n186;
  assign n188 = n476 | n186;
  assign n189 = ~n187 & n188;
  assign n190 = x3 & x12;
  assign n191 = n189 & n190;
  assign n192 = n189 | n190;
  assign n193 = ~n191 & n192;
  assign n194 = n474 & n193;
  assign n195 = n474 | n193;
  assign n196 = ~n194 & n195;
  assign n197 = x2 & x13;
  assign n198 = n196 & n197;
  assign n199 = n196 | n197;
  assign n200 = ~n198 & n199;
  assign n201 = n472 & n200;
  assign n202 = n472 | n200;
  assign n203 = ~n201 & n202;
  assign n204 = x1 & x14;
  assign n205 = n203 & n204;
  assign n206 = n203 | n204;
  assign n207 = ~n205 & n206;
  assign n208 = n160 & n207;
  assign n209 = n160 | n207;
  assign n210 = ~n208 & n209;
  assign n211 = x0 & x15;
  assign n212 = n210 & n211;
  assign n213 = n210 | n211;
  assign n214 = ~n212 & n213;
  assign n490 = n160 | n205;
  assign n491 = (n205 & n207) | (n205 & n490) | (n207 & n490);
  assign n216 = n198 | n201;
  assign n217 = n191 | n194;
  assign n492 = n184 | n186;
  assign n493 = (n184 & n476) | (n184 & n492) | (n476 & n492);
  assign n221 = x7 & x9;
  assign n497 = n170 & n221;
  assign n726 = (n172 & n221) | (n172 & n497) | (n221 & n497);
  assign n728 = (n478 & n726) | (n478 & n497) | (n726 & n497);
  assign n729 = (n600 & n726) | (n600 & n497) | (n726 & n497);
  assign n605 = (n453 & n728) | (n453 & n729) | (n728 & n729);
  assign n499 = n170 | n221;
  assign n730 = n172 | n499;
  assign n731 = (n478 & n499) | (n478 & n730) | (n499 & n730);
  assign n732 = (n499 & n600) | (n499 & n730) | (n600 & n730);
  assign n608 = (n453 & n731) | (n453 & n732) | (n731 & n732);
  assign n224 = ~n605 & n608;
  assign n225 = x6 & x10;
  assign n226 = n224 & n225;
  assign n227 = n224 | n225;
  assign n228 = ~n226 & n227;
  assign n495 = n177 | n179;
  assign n609 = n228 & n495;
  assign n601 = n132 | n177;
  assign n602 = (n177 & n179) | (n177 & n601) | (n179 & n601);
  assign n610 = n228 & n602;
  assign n611 = (n468 & n609) | (n468 & n610) | (n609 & n610);
  assign n612 = n228 | n495;
  assign n613 = n228 | n602;
  assign n614 = (n468 & n612) | (n468 & n613) | (n612 & n613);
  assign n231 = ~n611 & n614;
  assign n232 = x5 & x11;
  assign n233 = n231 & n232;
  assign n234 = n231 | n232;
  assign n235 = ~n233 & n234;
  assign n236 = n493 & n235;
  assign n237 = n493 | n235;
  assign n238 = ~n236 & n237;
  assign n239 = x4 & x12;
  assign n240 = n238 & n239;
  assign n241 = n238 | n239;
  assign n242 = ~n240 & n241;
  assign n243 = n217 & n242;
  assign n244 = n217 | n242;
  assign n245 = ~n243 & n244;
  assign n246 = x3 & x13;
  assign n247 = n245 & n246;
  assign n248 = n245 | n246;
  assign n249 = ~n247 & n248;
  assign n250 = n216 & n249;
  assign n251 = n216 | n249;
  assign n252 = ~n250 & n251;
  assign n253 = x2 & x14;
  assign n254 = n252 & n253;
  assign n255 = n252 | n253;
  assign n256 = ~n254 & n255;
  assign n257 = n491 & n256;
  assign n258 = n491 | n256;
  assign n259 = ~n257 & n258;
  assign n260 = x1 & x15;
  assign n261 = n259 & n260;
  assign n262 = n259 | n260;
  assign n263 = ~n261 & n262;
  assign n264 = n212 & n263;
  assign n265 = n212 | n263;
  assign n266 = ~n264 & n265;
  assign n733 = n211 | n260;
  assign n734 = (n210 & n260) | (n210 & n733) | (n260 & n733);
  assign n616 = (n212 & n259) | (n212 & n734) | (n259 & n734);
  assign n502 = (n261 & n263) | (n261 & n616) | (n263 & n616);
  assign n503 = n254 | n491;
  assign n504 = (n254 & n256) | (n254 & n503) | (n256 & n503);
  assign n269 = n247 | n250;
  assign n505 = n240 | n242;
  assign n506 = (n217 & n240) | (n217 & n505) | (n240 & n505);
  assign n273 = x7 & x10;
  assign n512 = n221 & n273;
  assign n617 = n170 & n512;
  assign n735 = (n172 & n512) | (n172 & n617) | (n512 & n617);
  assign n736 = n512 & n617;
  assign n737 = (n478 & n735) | (n478 & n736) | (n735 & n736);
  assign n738 = (n600 & n735) | (n600 & n736) | (n735 & n736);
  assign n620 = (n453 & n737) | (n453 & n738) | (n737 & n738);
  assign n515 = n221 | n273;
  assign n621 = (n170 & n273) | (n170 & n515) | (n273 & n515);
  assign n739 = (n172 & n515) | (n172 & n621) | (n515 & n621);
  assign n740 = n515 & n621;
  assign n741 = (n478 & n739) | (n478 & n740) | (n739 & n740);
  assign n742 = (n600 & n739) | (n600 & n740) | (n739 & n740);
  assign n624 = (n453 & n741) | (n453 & n742) | (n741 & n742);
  assign n276 = ~n620 & n624;
  assign n518 = n226 & n276;
  assign n625 = (n228 & n276) | (n228 & n518) | (n276 & n518);
  assign n626 = (n495 & n518) | (n495 & n625) | (n518 & n625);
  assign n627 = (n518 & n602) | (n518 & n625) | (n602 & n625);
  assign n628 = (n468 & n626) | (n468 & n627) | (n626 & n627);
  assign n521 = n226 | n276;
  assign n629 = n228 | n521;
  assign n630 = (n495 & n521) | (n495 & n629) | (n521 & n629);
  assign n631 = (n521 & n602) | (n521 & n629) | (n602 & n629);
  assign n632 = (n468 & n630) | (n468 & n631) | (n630 & n631);
  assign n279 = ~n628 & n632;
  assign n280 = x6 & x11;
  assign n281 = n279 & n280;
  assign n282 = n279 | n280;
  assign n283 = ~n281 & n282;
  assign n507 = n233 | n235;
  assign n633 = n283 & n507;
  assign n634 = n233 & n283;
  assign n635 = (n493 & n633) | (n493 & n634) | (n633 & n634);
  assign n636 = n283 | n507;
  assign n637 = n233 | n283;
  assign n638 = (n493 & n636) | (n493 & n637) | (n636 & n637);
  assign n286 = ~n635 & n638;
  assign n287 = x5 & x12;
  assign n288 = n286 & n287;
  assign n289 = n286 | n287;
  assign n290 = ~n288 & n289;
  assign n291 = n506 & n290;
  assign n292 = n506 | n290;
  assign n293 = ~n291 & n292;
  assign n294 = x4 & x13;
  assign n295 = n293 & n294;
  assign n296 = n293 | n294;
  assign n297 = ~n295 & n296;
  assign n298 = n269 & n297;
  assign n299 = n269 | n297;
  assign n300 = ~n298 & n299;
  assign n301 = x3 & x14;
  assign n302 = n300 & n301;
  assign n303 = n300 | n301;
  assign n304 = ~n302 & n303;
  assign n305 = n504 & n304;
  assign n306 = n504 | n304;
  assign n307 = ~n305 & n306;
  assign n308 = x2 & x15;
  assign n309 = n307 & n308;
  assign n310 = n307 | n308;
  assign n311 = ~n309 & n310;
  assign n312 = n502 & n311;
  assign n313 = n502 | n311;
  assign n314 = ~n312 & n313;
  assign n523 = n309 | n502;
  assign n524 = (n309 & n311) | (n309 & n523) | (n311 & n523);
  assign n525 = n302 | n504;
  assign n526 = (n302 & n304) | (n302 & n525) | (n304 & n525);
  assign n527 = n295 | n297;
  assign n528 = (n269 & n295) | (n269 & n527) | (n295 & n527);
  assign n321 = x7 & x11;
  assign n743 = n321 & n738;
  assign n744 = n321 & n737;
  assign n745 = (n453 & n743) | (n453 & n744) | (n743 & n744);
  assign n534 = (n321 & n628) | (n321 & n745) | (n628 & n745);
  assign n746 = n321 | n738;
  assign n747 = n321 | n737;
  assign n748 = (n453 & n746) | (n453 & n747) | (n746 & n747);
  assign n536 = n628 | n748;
  assign n324 = ~n534 & n536;
  assign n538 = n281 & n324;
  assign n639 = (n283 & n324) | (n283 & n538) | (n324 & n538);
  assign n640 = (n507 & n538) | (n507 & n639) | (n538 & n639);
  assign n641 = (n233 & n538) | (n233 & n639) | (n538 & n639);
  assign n642 = (n493 & n640) | (n493 & n641) | (n640 & n641);
  assign n541 = n281 | n324;
  assign n643 = n283 | n541;
  assign n644 = (n507 & n541) | (n507 & n643) | (n541 & n643);
  assign n645 = (n233 & n541) | (n233 & n643) | (n541 & n643);
  assign n646 = (n493 & n644) | (n493 & n645) | (n644 & n645);
  assign n327 = ~n642 & n646;
  assign n328 = x6 & x12;
  assign n329 = n327 & n328;
  assign n330 = n327 | n328;
  assign n331 = ~n329 & n330;
  assign n529 = n288 | n290;
  assign n647 = n331 & n529;
  assign n648 = n288 & n331;
  assign n649 = (n506 & n647) | (n506 & n648) | (n647 & n648);
  assign n650 = n331 | n529;
  assign n651 = n288 | n331;
  assign n652 = (n506 & n650) | (n506 & n651) | (n650 & n651);
  assign n334 = ~n649 & n652;
  assign n335 = x5 & x13;
  assign n336 = n334 & n335;
  assign n337 = n334 | n335;
  assign n338 = ~n336 & n337;
  assign n339 = n528 & n338;
  assign n340 = n528 | n338;
  assign n341 = ~n339 & n340;
  assign n342 = x4 & x14;
  assign n343 = n341 & n342;
  assign n344 = n341 | n342;
  assign n345 = ~n343 & n344;
  assign n346 = n526 & n345;
  assign n347 = n526 | n345;
  assign n348 = ~n346 & n347;
  assign n349 = x3 & x15;
  assign n350 = n348 & n349;
  assign n351 = n348 | n349;
  assign n352 = ~n350 & n351;
  assign n353 = n524 & n352;
  assign n354 = n524 | n352;
  assign n355 = ~n353 & n354;
  assign n356 = n350 | n353;
  assign n361 = x7 & x12;
  assign n653 = n361 & n745;
  assign n654 = n321 & n361;
  assign n655 = (n628 & n653) | (n628 & n654) | (n653 & n654);
  assign n548 = (n361 & n642) | (n361 & n655) | (n642 & n655);
  assign n656 = n361 | n745;
  assign n657 = n321 | n361;
  assign n658 = (n628 & n656) | (n628 & n657) | (n656 & n657);
  assign n550 = n642 | n658;
  assign n364 = ~n548 & n550;
  assign n552 = n329 & n364;
  assign n659 = (n331 & n364) | (n331 & n552) | (n364 & n552);
  assign n660 = (n529 & n552) | (n529 & n659) | (n552 & n659);
  assign n661 = (n288 & n552) | (n288 & n659) | (n552 & n659);
  assign n662 = (n506 & n660) | (n506 & n661) | (n660 & n661);
  assign n555 = n329 | n364;
  assign n663 = n331 | n555;
  assign n664 = (n529 & n555) | (n529 & n663) | (n555 & n663);
  assign n665 = (n288 & n555) | (n288 & n663) | (n555 & n663);
  assign n666 = (n506 & n664) | (n506 & n665) | (n664 & n665);
  assign n367 = ~n662 & n666;
  assign n368 = x6 & x13;
  assign n369 = n367 & n368;
  assign n370 = n367 | n368;
  assign n371 = ~n369 & n370;
  assign n543 = n336 | n338;
  assign n667 = n371 & n543;
  assign n668 = n336 & n371;
  assign n669 = (n528 & n667) | (n528 & n668) | (n667 & n668);
  assign n670 = n371 | n543;
  assign n671 = n336 | n371;
  assign n672 = (n528 & n670) | (n528 & n671) | (n670 & n671);
  assign n374 = ~n669 & n672;
  assign n375 = x5 & x14;
  assign n376 = n374 & n375;
  assign n377 = n374 | n375;
  assign n378 = ~n376 & n377;
  assign n673 = n343 & n378;
  assign n674 = (n346 & n378) | (n346 & n673) | (n378 & n673);
  assign n675 = n343 | n378;
  assign n676 = n346 | n675;
  assign n381 = ~n674 & n676;
  assign n382 = x4 & x15;
  assign n383 = n381 & n382;
  assign n384 = n381 | n382;
  assign n385 = ~n383 & n384;
  assign n386 = n356 & n385;
  assign n387 = n356 | n385;
  assign n388 = ~n386 & n387;
  assign n677 = n383 | n385;
  assign n678 = (n356 & n383) | (n356 & n677) | (n383 & n677);
  assign n357 = n343 | n346;
  assign n393 = x7 & x13;
  assign n680 = n361 & n393;
  assign n767 = n680 & n745;
  assign n750 = n393 & n654;
  assign n751 = (n628 & n767) | (n628 & n750) | (n767 & n750);
  assign n681 = (n642 & n751) | (n642 & n680) | (n751 & n680);
  assign n562 = (n393 & n662) | (n393 & n681) | (n662 & n681);
  assign n683 = n361 | n393;
  assign n768 = (n393 & n683) | (n393 & n745) | (n683 & n745);
  assign n753 = n393 | n654;
  assign n754 = (n628 & n768) | (n628 & n753) | (n768 & n753);
  assign n684 = (n642 & n754) | (n642 & n683) | (n754 & n683);
  assign n564 = n662 | n684;
  assign n396 = ~n562 & n564;
  assign n566 = n369 & n396;
  assign n685 = (n371 & n396) | (n371 & n566) | (n396 & n566);
  assign n686 = (n543 & n566) | (n543 & n685) | (n566 & n685);
  assign n687 = (n336 & n566) | (n336 & n685) | (n566 & n685);
  assign n688 = (n528 & n686) | (n528 & n687) | (n686 & n687);
  assign n569 = n369 | n396;
  assign n689 = n371 | n569;
  assign n690 = (n543 & n569) | (n543 & n689) | (n569 & n689);
  assign n691 = (n336 & n569) | (n336 & n689) | (n569 & n689);
  assign n692 = (n528 & n690) | (n528 & n691) | (n690 & n691);
  assign n399 = ~n688 & n692;
  assign n400 = x6 & x14;
  assign n401 = n399 & n400;
  assign n402 = n399 | n400;
  assign n403 = ~n401 & n402;
  assign n557 = n376 | n378;
  assign n693 = n403 & n557;
  assign n694 = n376 & n403;
  assign n695 = (n357 & n693) | (n357 & n694) | (n693 & n694);
  assign n696 = n403 | n557;
  assign n697 = n376 | n403;
  assign n698 = (n357 & n696) | (n357 & n697) | (n696 & n697);
  assign n406 = ~n695 & n698;
  assign n407 = x5 & x15;
  assign n408 = n406 & n407;
  assign n409 = n406 | n407;
  assign n410 = ~n408 & n409;
  assign n411 = n678 & n410;
  assign n412 = n678 | n410;
  assign n413 = ~n411 & n412;
  assign n571 = n408 | n410;
  assign n572 = (n678 & n408) | (n678 & n571) | (n408 & n571);
  assign n417 = x7 & x14;
  assign n756 = n417 & n680;
  assign n781 = n745 & n756;
  assign n700 = n393 & n417;
  assign n782 = n654 & n700;
  assign n771 = (n628 & n781) | (n628 & n782) | (n781 & n782);
  assign n757 = (n642 & n771) | (n642 & n756) | (n771 & n756);
  assign n701 = (n662 & n757) | (n662 & n700) | (n757 & n700);
  assign n576 = (n417 & n688) | (n417 & n701) | (n688 & n701);
  assign n759 = n417 | n680;
  assign n783 = (n417 & n745) | (n417 & n759) | (n745 & n759);
  assign n703 = n393 | n417;
  assign n784 = (n417 & n654) | (n417 & n703) | (n654 & n703);
  assign n774 = (n628 & n783) | (n628 & n784) | (n783 & n784);
  assign n760 = (n642 & n774) | (n642 & n759) | (n774 & n759);
  assign n704 = (n662 & n760) | (n662 & n703) | (n760 & n703);
  assign n578 = n688 | n704;
  assign n420 = ~n576 & n578;
  assign n580 = n401 & n420;
  assign n705 = (n403 & n420) | (n403 & n580) | (n420 & n580);
  assign n706 = (n557 & n580) | (n557 & n705) | (n580 & n705);
  assign n707 = (n376 & n580) | (n376 & n705) | (n580 & n705);
  assign n708 = (n357 & n706) | (n357 & n707) | (n706 & n707);
  assign n583 = n401 | n420;
  assign n709 = n403 | n583;
  assign n710 = (n557 & n583) | (n557 & n709) | (n583 & n709);
  assign n711 = (n376 & n583) | (n376 & n709) | (n583 & n709);
  assign n712 = (n357 & n710) | (n357 & n711) | (n710 & n711);
  assign n423 = ~n708 & n712;
  assign n424 = x6 & x15;
  assign n425 = n423 & n424;
  assign n426 = n423 | n424;
  assign n427 = ~n425 & n426;
  assign n428 = n572 & n427;
  assign n429 = n572 | n427;
  assign n430 = ~n428 & n429;
  assign n433 = x7 & x15;
  assign n714 = n417 & n433;
  assign n788 = n680 & n714;
  assign n793 = n745 & n788;
  assign n786 = n433 & n782;
  assign n787 = (n628 & n793) | (n628 & n786) | (n793 & n786);
  assign n777 = (n642 & n787) | (n642 & n788) | (n787 & n788);
  assign n762 = n433 & n700;
  assign n763 = (n662 & n777) | (n662 & n762) | (n777 & n762);
  assign n715 = (n688 & n763) | (n688 & n714) | (n763 & n714);
  assign n588 = (n433 & n708) | (n433 & n715) | (n708 & n715);
  assign n717 = n417 | n433;
  assign n792 = (n433 & n680) | (n433 & n717) | (n680 & n717);
  assign n794 = (n433 & n745) | (n433 & n792) | (n745 & n792);
  assign n790 = n433 | n782;
  assign n791 = (n628 & n794) | (n628 & n790) | (n794 & n790);
  assign n780 = (n642 & n791) | (n642 & n792) | (n791 & n792);
  assign n765 = n433 | n700;
  assign n766 = (n662 & n780) | (n662 & n765) | (n780 & n765);
  assign n718 = (n688 & n766) | (n688 & n717) | (n766 & n717);
  assign n590 = n708 | n718;
  assign n436 = ~n588 & n590;
  assign n592 = n425 & n436;
  assign n719 = (n427 & n436) | (n427 & n592) | (n436 & n592);
  assign n593 = (n572 & n719) | (n572 & n592) | (n719 & n592);
  assign n595 = n425 | n436;
  assign n720 = n427 | n595;
  assign n596 = (n572 & n720) | (n572 & n595) | (n720 & n595);
  assign n439 = ~n593 & n596;
  assign n721 = n588 | n719;
  assign n722 = n588 | n592;
  assign n723 = (n572 & n721) | (n572 & n722) | (n721 & n722);
  assign n827 = x16 & x32;
  assign n828 = x17 & x32;
  assign n829 = x16 & x33;
  assign n830 = n828 & n829;
  assign n831 = n828 | n829;
  assign n832 = ~n830 & n831;
  assign n833 = x18 & x32;
  assign n834 = x17 & x33;
  assign n835 = n833 & n834;
  assign n836 = n833 | n834;
  assign n837 = ~n835 & n836;
  assign n838 = n830 & n837;
  assign n839 = n830 | n837;
  assign n840 = ~n838 & n839;
  assign n841 = x16 & x34;
  assign n842 = n840 & n841;
  assign n843 = n840 | n841;
  assign n844 = ~n842 & n843;
  assign n2699 = n830 | n835;
  assign n2700 = (n835 & n837) | (n835 & n2699) | (n837 & n2699);
  assign n846 = x19 & x32;
  assign n847 = x18 & x33;
  assign n848 = n846 & n847;
  assign n849 = n846 | n847;
  assign n850 = ~n848 & n849;
  assign n851 = n2700 & n850;
  assign n852 = n2700 | n850;
  assign n853 = ~n851 & n852;
  assign n854 = x17 & x34;
  assign n855 = n853 & n854;
  assign n856 = n853 | n854;
  assign n857 = ~n855 & n856;
  assign n858 = n842 & n857;
  assign n859 = n842 | n857;
  assign n860 = ~n858 & n859;
  assign n861 = x16 & x35;
  assign n862 = n860 & n861;
  assign n863 = n860 | n861;
  assign n864 = ~n862 & n863;
  assign n2701 = n842 | n855;
  assign n2702 = (n855 & n857) | (n855 & n2701) | (n857 & n2701);
  assign n2703 = n848 | n850;
  assign n2704 = (n848 & n2700) | (n848 & n2703) | (n2700 & n2703);
  assign n867 = x20 & x32;
  assign n868 = x19 & x33;
  assign n869 = n867 & n868;
  assign n870 = n867 | n868;
  assign n871 = ~n869 & n870;
  assign n872 = n2704 & n871;
  assign n873 = n2704 | n871;
  assign n874 = ~n872 & n873;
  assign n875 = x18 & x34;
  assign n876 = n874 & n875;
  assign n877 = n874 | n875;
  assign n878 = ~n876 & n877;
  assign n879 = n2702 & n878;
  assign n880 = n2702 | n878;
  assign n881 = ~n879 & n880;
  assign n882 = x17 & x35;
  assign n883 = n881 & n882;
  assign n884 = n881 | n882;
  assign n885 = ~n883 & n884;
  assign n886 = n862 & n885;
  assign n887 = n862 | n885;
  assign n888 = ~n886 & n887;
  assign n889 = x16 & x36;
  assign n890 = n888 & n889;
  assign n891 = n888 | n889;
  assign n892 = ~n890 & n891;
  assign n2705 = n862 | n883;
  assign n2706 = (n883 & n885) | (n883 & n2705) | (n885 & n2705);
  assign n896 = x21 & x32;
  assign n897 = x20 & x33;
  assign n898 = n896 & n897;
  assign n899 = n896 | n897;
  assign n900 = ~n898 & n899;
  assign n2707 = n869 | n871;
  assign n2709 = n900 & n2707;
  assign n2710 = n869 & n900;
  assign n2711 = (n2704 & n2709) | (n2704 & n2710) | (n2709 & n2710);
  assign n2712 = n900 | n2707;
  assign n2713 = n869 | n900;
  assign n2714 = (n2704 & n2712) | (n2704 & n2713) | (n2712 & n2713);
  assign n903 = ~n2711 & n2714;
  assign n904 = x19 & x34;
  assign n905 = n903 & n904;
  assign n906 = n903 | n904;
  assign n907 = ~n905 & n906;
  assign n2715 = n876 & n907;
  assign n2716 = (n879 & n907) | (n879 & n2715) | (n907 & n2715);
  assign n2717 = n876 | n907;
  assign n2718 = n879 | n2717;
  assign n910 = ~n2716 & n2718;
  assign n911 = x18 & x35;
  assign n912 = n910 & n911;
  assign n913 = n910 | n911;
  assign n914 = ~n912 & n913;
  assign n915 = n2706 & n914;
  assign n916 = n2706 | n914;
  assign n917 = ~n915 & n916;
  assign n918 = x17 & x36;
  assign n919 = n917 & n918;
  assign n920 = n917 | n918;
  assign n921 = ~n919 & n920;
  assign n922 = n890 & n921;
  assign n923 = n890 | n921;
  assign n924 = ~n922 & n923;
  assign n925 = x16 & x37;
  assign n926 = n924 & n925;
  assign n927 = n924 | n925;
  assign n928 = ~n926 & n927;
  assign n2719 = n890 | n919;
  assign n2720 = (n919 & n921) | (n919 & n2719) | (n921 & n2719);
  assign n930 = n912 | n915;
  assign n933 = x22 & x32;
  assign n934 = x21 & x33;
  assign n935 = n933 & n934;
  assign n936 = n933 | n934;
  assign n937 = ~n935 & n936;
  assign n2721 = n898 & n937;
  assign n2722 = (n937 & n2711) | (n937 & n2721) | (n2711 & n2721);
  assign n2723 = n898 | n937;
  assign n2724 = n2711 | n2723;
  assign n940 = ~n2722 & n2724;
  assign n941 = x20 & x34;
  assign n942 = n940 & n941;
  assign n943 = n940 | n941;
  assign n944 = ~n942 & n943;
  assign n2725 = n905 & n944;
  assign n2726 = (n944 & n2716) | (n944 & n2725) | (n2716 & n2725);
  assign n2727 = n905 | n944;
  assign n2728 = n2716 | n2727;
  assign n947 = ~n2726 & n2728;
  assign n948 = x19 & x35;
  assign n949 = n947 & n948;
  assign n950 = n947 | n948;
  assign n951 = ~n949 & n950;
  assign n952 = n930 & n951;
  assign n953 = n930 | n951;
  assign n954 = ~n952 & n953;
  assign n955 = x18 & x36;
  assign n956 = n954 & n955;
  assign n957 = n954 | n955;
  assign n958 = ~n956 & n957;
  assign n959 = n2720 & n958;
  assign n960 = n2720 | n958;
  assign n961 = ~n959 & n960;
  assign n962 = x17 & x37;
  assign n963 = n961 & n962;
  assign n964 = n961 | n962;
  assign n965 = ~n963 & n964;
  assign n966 = n926 & n965;
  assign n967 = n926 | n965;
  assign n968 = ~n966 & n967;
  assign n969 = x16 & x38;
  assign n970 = n968 & n969;
  assign n971 = n968 | n969;
  assign n972 = ~n970 & n971;
  assign n3897 = n925 | n962;
  assign n3898 = (n924 & n962) | (n924 & n3897) | (n962 & n3897);
  assign n3444 = (n926 & n961) | (n926 & n3898) | (n961 & n3898);
  assign n2730 = (n963 & n965) | (n963 & n3444) | (n965 & n3444);
  assign n2731 = n956 | n2720;
  assign n2732 = (n956 & n958) | (n956 & n2731) | (n958 & n2731);
  assign n2733 = n949 | n951;
  assign n2734 = (n930 & n949) | (n930 & n2733) | (n949 & n2733);
  assign n978 = x23 & x32;
  assign n979 = x22 & x33;
  assign n980 = n978 & n979;
  assign n981 = n978 | n979;
  assign n982 = ~n980 & n981;
  assign n3445 = n898 | n935;
  assign n3446 = (n935 & n937) | (n935 & n3445) | (n937 & n3445);
  assign n2738 = n982 & n3446;
  assign n2736 = n935 | n937;
  assign n2739 = n982 & n2736;
  assign n2740 = (n2711 & n2738) | (n2711 & n2739) | (n2738 & n2739);
  assign n2741 = n982 | n3446;
  assign n2742 = n982 | n2736;
  assign n2743 = (n2711 & n2741) | (n2711 & n2742) | (n2741 & n2742);
  assign n985 = ~n2740 & n2743;
  assign n986 = x21 & x34;
  assign n987 = n985 & n986;
  assign n988 = n985 | n986;
  assign n989 = ~n987 & n988;
  assign n2744 = n942 & n989;
  assign n2745 = (n989 & n2726) | (n989 & n2744) | (n2726 & n2744);
  assign n2746 = n942 | n989;
  assign n2747 = n2726 | n2746;
  assign n992 = ~n2745 & n2747;
  assign n993 = x20 & x35;
  assign n994 = n992 & n993;
  assign n995 = n992 | n993;
  assign n996 = ~n994 & n995;
  assign n997 = n2734 & n996;
  assign n998 = n2734 | n996;
  assign n999 = ~n997 & n998;
  assign n1000 = x19 & x36;
  assign n1001 = n999 & n1000;
  assign n1002 = n999 | n1000;
  assign n1003 = ~n1001 & n1002;
  assign n1004 = n2732 & n1003;
  assign n1005 = n2732 | n1003;
  assign n1006 = ~n1004 & n1005;
  assign n1007 = x18 & x37;
  assign n1008 = n1006 & n1007;
  assign n1009 = n1006 | n1007;
  assign n1010 = ~n1008 & n1009;
  assign n1011 = n2730 & n1010;
  assign n1012 = n2730 | n1010;
  assign n1013 = ~n1011 & n1012;
  assign n1014 = x17 & x38;
  assign n1015 = n1013 & n1014;
  assign n1016 = n1013 | n1014;
  assign n1017 = ~n1015 & n1016;
  assign n1018 = n970 & n1017;
  assign n1019 = n970 | n1017;
  assign n1020 = ~n1018 & n1019;
  assign n1021 = x16 & x39;
  assign n1022 = n1020 & n1021;
  assign n1023 = n1020 | n1021;
  assign n1024 = ~n1022 & n1023;
  assign n2748 = n970 | n1015;
  assign n2749 = (n1015 & n1017) | (n1015 & n2748) | (n1017 & n2748);
  assign n1026 = n1008 | n1011;
  assign n1027 = n1001 | n1004;
  assign n2750 = n994 | n996;
  assign n2751 = (n994 & n2734) | (n994 & n2750) | (n2734 & n2750);
  assign n1031 = x24 & x32;
  assign n1032 = x23 & x33;
  assign n1033 = n1031 & n1032;
  assign n1034 = n1031 | n1032;
  assign n1035 = ~n1033 & n1034;
  assign n2755 = n980 & n1035;
  assign n3449 = (n1035 & n2739) | (n1035 & n2755) | (n2739 & n2755);
  assign n3450 = (n1035 & n2738) | (n1035 & n2755) | (n2738 & n2755);
  assign n3451 = (n2711 & n3449) | (n2711 & n3450) | (n3449 & n3450);
  assign n2757 = n980 | n1035;
  assign n3452 = n2739 | n2757;
  assign n3453 = n2738 | n2757;
  assign n3454 = (n2711 & n3452) | (n2711 & n3453) | (n3452 & n3453);
  assign n1038 = ~n3451 & n3454;
  assign n1039 = x22 & x34;
  assign n1040 = n1038 & n1039;
  assign n1041 = n1038 | n1039;
  assign n1042 = ~n1040 & n1041;
  assign n2753 = n987 | n989;
  assign n3455 = n1042 & n2753;
  assign n3447 = n942 | n987;
  assign n3448 = (n987 & n989) | (n987 & n3447) | (n989 & n3447);
  assign n3456 = n1042 & n3448;
  assign n3457 = (n2726 & n3455) | (n2726 & n3456) | (n3455 & n3456);
  assign n3458 = n1042 | n2753;
  assign n3459 = n1042 | n3448;
  assign n3460 = (n2726 & n3458) | (n2726 & n3459) | (n3458 & n3459);
  assign n1045 = ~n3457 & n3460;
  assign n1046 = x21 & x35;
  assign n1047 = n1045 & n1046;
  assign n1048 = n1045 | n1046;
  assign n1049 = ~n1047 & n1048;
  assign n1050 = n2751 & n1049;
  assign n1051 = n2751 | n1049;
  assign n1052 = ~n1050 & n1051;
  assign n1053 = x20 & x36;
  assign n1054 = n1052 & n1053;
  assign n1055 = n1052 | n1053;
  assign n1056 = ~n1054 & n1055;
  assign n1057 = n1027 & n1056;
  assign n1058 = n1027 | n1056;
  assign n1059 = ~n1057 & n1058;
  assign n1060 = x19 & x37;
  assign n1061 = n1059 & n1060;
  assign n1062 = n1059 | n1060;
  assign n1063 = ~n1061 & n1062;
  assign n1064 = n1026 & n1063;
  assign n1065 = n1026 | n1063;
  assign n1066 = ~n1064 & n1065;
  assign n1067 = x18 & x38;
  assign n1068 = n1066 & n1067;
  assign n1069 = n1066 | n1067;
  assign n1070 = ~n1068 & n1069;
  assign n1071 = n2749 & n1070;
  assign n1072 = n2749 | n1070;
  assign n1073 = ~n1071 & n1072;
  assign n1074 = x17 & x39;
  assign n1075 = n1073 & n1074;
  assign n1076 = n1073 | n1074;
  assign n1077 = ~n1075 & n1076;
  assign n1078 = n1022 & n1077;
  assign n1079 = n1022 | n1077;
  assign n1080 = ~n1078 & n1079;
  assign n1081 = x16 & x40;
  assign n1082 = n1080 & n1081;
  assign n1083 = n1080 | n1081;
  assign n1084 = ~n1082 & n1083;
  assign n3899 = n1021 | n1074;
  assign n3900 = (n1020 & n1074) | (n1020 & n3899) | (n1074 & n3899);
  assign n3462 = (n1022 & n1073) | (n1022 & n3900) | (n1073 & n3900);
  assign n2760 = (n1075 & n1077) | (n1075 & n3462) | (n1077 & n3462);
  assign n2761 = n1068 | n2749;
  assign n2762 = (n1068 & n1070) | (n1068 & n2761) | (n1070 & n2761);
  assign n1087 = n1061 | n1064;
  assign n2763 = n1054 | n1056;
  assign n2764 = (n1027 & n1054) | (n1027 & n2763) | (n1054 & n2763);
  assign n2754 = (n2726 & n3448) | (n2726 & n2753) | (n3448 & n2753);
  assign n1092 = x25 & x32;
  assign n1093 = x24 & x33;
  assign n1094 = n1092 & n1093;
  assign n1095 = n1092 | n1093;
  assign n1096 = ~n1094 & n1095;
  assign n3463 = n980 | n1033;
  assign n3464 = (n1033 & n1035) | (n1033 & n3463) | (n1035 & n3463);
  assign n2772 = n1096 & n3464;
  assign n2770 = n1033 | n1035;
  assign n2773 = n1096 & n2770;
  assign n3465 = (n2739 & n2772) | (n2739 & n2773) | (n2772 & n2773);
  assign n3466 = (n2738 & n2772) | (n2738 & n2773) | (n2772 & n2773);
  assign n3467 = (n2711 & n3465) | (n2711 & n3466) | (n3465 & n3466);
  assign n2775 = n1096 | n3464;
  assign n2776 = n1096 | n2770;
  assign n3468 = (n2739 & n2775) | (n2739 & n2776) | (n2775 & n2776);
  assign n3469 = (n2738 & n2775) | (n2738 & n2776) | (n2775 & n2776);
  assign n3470 = (n2711 & n3468) | (n2711 & n3469) | (n3468 & n3469);
  assign n1099 = ~n3467 & n3470;
  assign n1100 = x23 & x34;
  assign n1101 = n1099 & n1100;
  assign n1102 = n1099 | n1100;
  assign n1103 = ~n1101 & n1102;
  assign n2767 = n1040 | n1042;
  assign n2778 = n1103 & n2767;
  assign n2779 = n1040 & n1103;
  assign n2780 = (n2754 & n2778) | (n2754 & n2779) | (n2778 & n2779);
  assign n2781 = n1103 | n2767;
  assign n2782 = n1040 | n1103;
  assign n2783 = (n2754 & n2781) | (n2754 & n2782) | (n2781 & n2782);
  assign n1106 = ~n2780 & n2783;
  assign n1107 = x22 & x35;
  assign n1108 = n1106 & n1107;
  assign n1109 = n1106 | n1107;
  assign n1110 = ~n1108 & n1109;
  assign n2765 = n1047 | n1049;
  assign n3471 = n1110 & n2765;
  assign n3472 = n1047 & n1110;
  assign n3473 = (n2751 & n3471) | (n2751 & n3472) | (n3471 & n3472);
  assign n3474 = n1110 | n2765;
  assign n3475 = n1047 | n1110;
  assign n3476 = (n2751 & n3474) | (n2751 & n3475) | (n3474 & n3475);
  assign n1113 = ~n3473 & n3476;
  assign n1114 = x21 & x36;
  assign n1115 = n1113 & n1114;
  assign n1116 = n1113 | n1114;
  assign n1117 = ~n1115 & n1116;
  assign n1118 = n2764 & n1117;
  assign n1119 = n2764 | n1117;
  assign n1120 = ~n1118 & n1119;
  assign n1121 = x20 & x37;
  assign n1122 = n1120 & n1121;
  assign n1123 = n1120 | n1121;
  assign n1124 = ~n1122 & n1123;
  assign n1125 = n1087 & n1124;
  assign n1126 = n1087 | n1124;
  assign n1127 = ~n1125 & n1126;
  assign n1128 = x19 & x38;
  assign n1129 = n1127 & n1128;
  assign n1130 = n1127 | n1128;
  assign n1131 = ~n1129 & n1130;
  assign n1132 = n2762 & n1131;
  assign n1133 = n2762 | n1131;
  assign n1134 = ~n1132 & n1133;
  assign n1135 = x18 & x39;
  assign n1136 = n1134 & n1135;
  assign n1137 = n1134 | n1135;
  assign n1138 = ~n1136 & n1137;
  assign n1139 = n2760 & n1138;
  assign n1140 = n2760 | n1138;
  assign n1141 = ~n1139 & n1140;
  assign n1142 = x17 & x40;
  assign n1143 = n1141 & n1142;
  assign n1144 = n1141 | n1142;
  assign n1145 = ~n1143 & n1144;
  assign n1146 = n1082 & n1145;
  assign n1147 = n1082 | n1145;
  assign n1148 = ~n1146 & n1147;
  assign n1149 = x16 & x41;
  assign n1150 = n1148 & n1149;
  assign n1151 = n1148 | n1149;
  assign n1152 = ~n1150 & n1151;
  assign n3901 = n1081 | n1142;
  assign n3902 = (n1080 & n1142) | (n1080 & n3901) | (n1142 & n3901);
  assign n3478 = (n1082 & n1141) | (n1082 & n3902) | (n1141 & n3902);
  assign n2785 = (n1143 & n1145) | (n1143 & n3478) | (n1145 & n3478);
  assign n2786 = n1136 | n2760;
  assign n2787 = (n1136 & n1138) | (n1136 & n2786) | (n1138 & n2786);
  assign n2788 = n1129 | n2762;
  assign n2789 = (n1129 & n1131) | (n1129 & n2788) | (n1131 & n2788);
  assign n2790 = n1122 | n1124;
  assign n2791 = (n1087 & n1122) | (n1087 & n2790) | (n1122 & n2790);
  assign n2766 = (n1047 & n2751) | (n1047 & n2765) | (n2751 & n2765);
  assign n3479 = n1094 | n1096;
  assign n3480 = (n1094 & n3464) | (n1094 & n3479) | (n3464 & n3479);
  assign n3481 = (n1094 & n2770) | (n1094 & n3479) | (n2770 & n3479);
  assign n3482 = (n2739 & n3480) | (n2739 & n3481) | (n3480 & n3481);
  assign n3483 = (n2738 & n3480) | (n2738 & n3481) | (n3480 & n3481);
  assign n3484 = (n2711 & n3482) | (n2711 & n3483) | (n3482 & n3483);
  assign n1161 = x26 & x32;
  assign n1162 = x25 & x33;
  assign n1163 = n1161 & n1162;
  assign n1164 = n1161 | n1162;
  assign n1165 = ~n1163 & n1164;
  assign n1166 = n3484 & n1165;
  assign n1167 = n3484 | n1165;
  assign n1168 = ~n1166 & n1167;
  assign n1169 = x24 & x34;
  assign n1170 = n1168 & n1169;
  assign n1171 = n1168 | n1169;
  assign n1172 = ~n1170 & n1171;
  assign n2799 = n1101 & n1172;
  assign n3485 = (n1172 & n2778) | (n1172 & n2799) | (n2778 & n2799);
  assign n3486 = (n1172 & n2779) | (n1172 & n2799) | (n2779 & n2799);
  assign n3487 = (n2754 & n3485) | (n2754 & n3486) | (n3485 & n3486);
  assign n2801 = n1101 | n1172;
  assign n3488 = n2778 | n2801;
  assign n3489 = n2779 | n2801;
  assign n3490 = (n2754 & n3488) | (n2754 & n3489) | (n3488 & n3489);
  assign n1175 = ~n3487 & n3490;
  assign n1176 = x23 & x35;
  assign n1177 = n1175 & n1176;
  assign n1178 = n1175 | n1176;
  assign n1179 = ~n1177 & n1178;
  assign n2794 = n1108 | n1110;
  assign n2803 = n1179 & n2794;
  assign n2804 = n1108 & n1179;
  assign n2805 = (n2766 & n2803) | (n2766 & n2804) | (n2803 & n2804);
  assign n2806 = n1179 | n2794;
  assign n2807 = n1108 | n1179;
  assign n2808 = (n2766 & n2806) | (n2766 & n2807) | (n2806 & n2807);
  assign n1182 = ~n2805 & n2808;
  assign n1183 = x22 & x36;
  assign n1184 = n1182 & n1183;
  assign n1185 = n1182 | n1183;
  assign n1186 = ~n1184 & n1185;
  assign n2792 = n1115 | n1117;
  assign n3491 = n1186 & n2792;
  assign n3492 = n1115 & n1186;
  assign n3493 = (n2764 & n3491) | (n2764 & n3492) | (n3491 & n3492);
  assign n3494 = n1186 | n2792;
  assign n3495 = n1115 | n1186;
  assign n3496 = (n2764 & n3494) | (n2764 & n3495) | (n3494 & n3495);
  assign n1189 = ~n3493 & n3496;
  assign n1190 = x21 & x37;
  assign n1191 = n1189 & n1190;
  assign n1192 = n1189 | n1190;
  assign n1193 = ~n1191 & n1192;
  assign n1194 = n2791 & n1193;
  assign n1195 = n2791 | n1193;
  assign n1196 = ~n1194 & n1195;
  assign n1197 = x20 & x38;
  assign n1198 = n1196 & n1197;
  assign n1199 = n1196 | n1197;
  assign n1200 = ~n1198 & n1199;
  assign n1201 = n2789 & n1200;
  assign n1202 = n2789 | n1200;
  assign n1203 = ~n1201 & n1202;
  assign n1204 = x19 & x39;
  assign n1205 = n1203 & n1204;
  assign n1206 = n1203 | n1204;
  assign n1207 = ~n1205 & n1206;
  assign n1208 = n2787 & n1207;
  assign n1209 = n2787 | n1207;
  assign n1210 = ~n1208 & n1209;
  assign n1211 = x18 & x40;
  assign n1212 = n1210 & n1211;
  assign n1213 = n1210 | n1211;
  assign n1214 = ~n1212 & n1213;
  assign n1215 = n2785 & n1214;
  assign n1216 = n2785 | n1214;
  assign n1217 = ~n1215 & n1216;
  assign n1218 = x17 & x41;
  assign n1219 = n1217 & n1218;
  assign n1220 = n1217 | n1218;
  assign n1221 = ~n1219 & n1220;
  assign n1222 = n1150 & n1221;
  assign n1223 = n1150 | n1221;
  assign n1224 = ~n1222 & n1223;
  assign n1225 = x16 & x42;
  assign n1226 = n1224 & n1225;
  assign n1227 = n1224 | n1225;
  assign n1228 = ~n1226 & n1227;
  assign n2809 = n1150 | n1219;
  assign n2810 = (n1219 & n1221) | (n1219 & n2809) | (n1221 & n2809);
  assign n1230 = n1212 | n1215;
  assign n1231 = n1205 | n1208;
  assign n2793 = (n1115 & n2764) | (n1115 & n2792) | (n2764 & n2792);
  assign n2816 = n1170 | n1172;
  assign n3497 = n1101 | n1170;
  assign n3498 = (n1170 & n1172) | (n1170 & n3497) | (n1172 & n3497);
  assign n3499 = (n2778 & n2816) | (n2778 & n3498) | (n2816 & n3498);
  assign n3500 = (n2779 & n2816) | (n2779 & n3498) | (n2816 & n3498);
  assign n3501 = (n2754 & n3499) | (n2754 & n3500) | (n3499 & n3500);
  assign n1238 = x27 & x32;
  assign n1239 = x26 & x33;
  assign n1240 = n1238 & n1239;
  assign n1241 = n1238 | n1239;
  assign n1242 = ~n1240 & n1241;
  assign n2818 = n1163 | n1165;
  assign n2820 = n1242 & n2818;
  assign n2821 = n1163 & n1242;
  assign n2822 = (n3484 & n2820) | (n3484 & n2821) | (n2820 & n2821);
  assign n2823 = n1242 | n2818;
  assign n2824 = n1163 | n1242;
  assign n2825 = (n3484 & n2823) | (n3484 & n2824) | (n2823 & n2824);
  assign n1245 = ~n2822 & n2825;
  assign n1246 = x25 & x34;
  assign n1247 = n1245 & n1246;
  assign n1248 = n1245 | n1246;
  assign n1249 = ~n1247 & n1248;
  assign n1250 = n3501 & n1249;
  assign n1251 = n3501 | n1249;
  assign n1252 = ~n1250 & n1251;
  assign n1253 = x24 & x35;
  assign n1254 = n1252 & n1253;
  assign n1255 = n1252 | n1253;
  assign n1256 = ~n1254 & n1255;
  assign n2826 = n1177 & n1256;
  assign n2827 = (n1256 & n2805) | (n1256 & n2826) | (n2805 & n2826);
  assign n2828 = n1177 | n1256;
  assign n2829 = n2805 | n2828;
  assign n1259 = ~n2827 & n2829;
  assign n1260 = x23 & x36;
  assign n1261 = n1259 & n1260;
  assign n1262 = n1259 | n1260;
  assign n1263 = ~n1261 & n1262;
  assign n2813 = n1184 | n1186;
  assign n2830 = n1263 & n2813;
  assign n2831 = n1184 & n1263;
  assign n2832 = (n2793 & n2830) | (n2793 & n2831) | (n2830 & n2831);
  assign n2833 = n1263 | n2813;
  assign n2834 = n1184 | n1263;
  assign n2835 = (n2793 & n2833) | (n2793 & n2834) | (n2833 & n2834);
  assign n1266 = ~n2832 & n2835;
  assign n1267 = x22 & x37;
  assign n1268 = n1266 & n1267;
  assign n1269 = n1266 | n1267;
  assign n1270 = ~n1268 & n1269;
  assign n2811 = n1191 | n1193;
  assign n3502 = n1270 & n2811;
  assign n3503 = n1191 & n1270;
  assign n3504 = (n2791 & n3502) | (n2791 & n3503) | (n3502 & n3503);
  assign n3505 = n1270 | n2811;
  assign n3506 = n1191 | n1270;
  assign n3507 = (n2791 & n3505) | (n2791 & n3506) | (n3505 & n3506);
  assign n1273 = ~n3504 & n3507;
  assign n1274 = x21 & x38;
  assign n1275 = n1273 & n1274;
  assign n1276 = n1273 | n1274;
  assign n1277 = ~n1275 & n1276;
  assign n3508 = n1198 & n1277;
  assign n3509 = (n1201 & n1277) | (n1201 & n3508) | (n1277 & n3508);
  assign n3510 = n1198 | n1277;
  assign n3511 = n1201 | n3510;
  assign n1280 = ~n3509 & n3511;
  assign n1281 = x20 & x39;
  assign n1282 = n1280 & n1281;
  assign n1283 = n1280 | n1281;
  assign n1284 = ~n1282 & n1283;
  assign n1285 = n1231 & n1284;
  assign n1286 = n1231 | n1284;
  assign n1287 = ~n1285 & n1286;
  assign n1288 = x19 & x40;
  assign n1289 = n1287 & n1288;
  assign n1290 = n1287 | n1288;
  assign n1291 = ~n1289 & n1290;
  assign n1292 = n1230 & n1291;
  assign n1293 = n1230 | n1291;
  assign n1294 = ~n1292 & n1293;
  assign n1295 = x18 & x41;
  assign n1296 = n1294 & n1295;
  assign n1297 = n1294 | n1295;
  assign n1298 = ~n1296 & n1297;
  assign n1299 = n2810 & n1298;
  assign n1300 = n2810 | n1298;
  assign n1301 = ~n1299 & n1300;
  assign n1302 = x17 & x42;
  assign n1303 = n1301 & n1302;
  assign n1304 = n1301 | n1302;
  assign n1305 = ~n1303 & n1304;
  assign n1306 = n1226 & n1305;
  assign n1307 = n1226 | n1305;
  assign n1308 = ~n1306 & n1307;
  assign n1309 = x16 & x43;
  assign n1310 = n1308 & n1309;
  assign n1311 = n1308 | n1309;
  assign n1312 = ~n1310 & n1311;
  assign n3903 = n1225 | n1302;
  assign n3904 = (n1224 & n1302) | (n1224 & n3903) | (n1302 & n3903);
  assign n3513 = (n1226 & n1301) | (n1226 & n3904) | (n1301 & n3904);
  assign n2837 = (n1303 & n1305) | (n1303 & n3513) | (n1305 & n3513);
  assign n2838 = n1296 | n2810;
  assign n2839 = (n1296 & n1298) | (n1296 & n2838) | (n1298 & n2838);
  assign n1315 = n1289 | n1292;
  assign n3514 = n1282 | n1284;
  assign n3515 = (n1231 & n1282) | (n1231 & n3514) | (n1282 & n3514);
  assign n1232 = n1198 | n1201;
  assign n2812 = (n1191 & n2791) | (n1191 & n2811) | (n2791 & n2811);
  assign n1323 = x28 & x32;
  assign n1324 = x27 & x33;
  assign n1325 = n1323 & n1324;
  assign n1326 = n1323 | n1324;
  assign n1327 = ~n1325 & n1326;
  assign n3516 = n1240 | n1242;
  assign n3517 = (n1240 & n2818) | (n1240 & n3516) | (n2818 & n3516);
  assign n2849 = n1327 & n3517;
  assign n3518 = n1163 | n1240;
  assign n3519 = (n1240 & n1242) | (n1240 & n3518) | (n1242 & n3518);
  assign n2850 = n1327 & n3519;
  assign n2851 = (n3484 & n2849) | (n3484 & n2850) | (n2849 & n2850);
  assign n2852 = n1327 | n3517;
  assign n2853 = n1327 | n3519;
  assign n2854 = (n3484 & n2852) | (n3484 & n2853) | (n2852 & n2853);
  assign n1330 = ~n2851 & n2854;
  assign n1331 = x26 & x34;
  assign n1332 = n1330 & n1331;
  assign n1333 = n1330 | n1331;
  assign n1334 = ~n1332 & n1333;
  assign n2844 = n1247 | n1249;
  assign n2855 = n1334 & n2844;
  assign n2856 = n1247 & n1334;
  assign n2857 = (n3501 & n2855) | (n3501 & n2856) | (n2855 & n2856);
  assign n2858 = n1334 | n2844;
  assign n2859 = n1247 | n1334;
  assign n2860 = (n3501 & n2858) | (n3501 & n2859) | (n2858 & n2859);
  assign n1337 = ~n2857 & n2860;
  assign n1338 = x25 & x35;
  assign n1339 = n1337 & n1338;
  assign n1340 = n1337 | n1338;
  assign n1341 = ~n1339 & n1340;
  assign n2861 = n1254 & n1341;
  assign n3520 = (n1341 & n2826) | (n1341 & n2861) | (n2826 & n2861);
  assign n3521 = (n1256 & n1341) | (n1256 & n2861) | (n1341 & n2861);
  assign n3522 = (n2805 & n3520) | (n2805 & n3521) | (n3520 & n3521);
  assign n2863 = n1254 | n1341;
  assign n3523 = n2826 | n2863;
  assign n3524 = n1256 | n2863;
  assign n3525 = (n2805 & n3523) | (n2805 & n3524) | (n3523 & n3524);
  assign n1344 = ~n3522 & n3525;
  assign n1345 = x24 & x36;
  assign n1346 = n1344 & n1345;
  assign n1347 = n1344 | n1345;
  assign n1348 = ~n1346 & n1347;
  assign n2865 = n1261 & n1348;
  assign n2866 = (n1348 & n2832) | (n1348 & n2865) | (n2832 & n2865);
  assign n2867 = n1261 | n1348;
  assign n2868 = n2832 | n2867;
  assign n1351 = ~n2866 & n2868;
  assign n1352 = x23 & x37;
  assign n1353 = n1351 & n1352;
  assign n1354 = n1351 | n1352;
  assign n1355 = ~n1353 & n1354;
  assign n2842 = n1268 | n1270;
  assign n2869 = n1355 & n2842;
  assign n2870 = n1268 & n1355;
  assign n2871 = (n2812 & n2869) | (n2812 & n2870) | (n2869 & n2870);
  assign n2872 = n1355 | n2842;
  assign n2873 = n1268 | n1355;
  assign n2874 = (n2812 & n2872) | (n2812 & n2873) | (n2872 & n2873);
  assign n1358 = ~n2871 & n2874;
  assign n1359 = x22 & x38;
  assign n1360 = n1358 & n1359;
  assign n1361 = n1358 | n1359;
  assign n1362 = ~n1360 & n1361;
  assign n2840 = n1275 | n1277;
  assign n3526 = n1362 & n2840;
  assign n3527 = n1275 & n1362;
  assign n3528 = (n1232 & n3526) | (n1232 & n3527) | (n3526 & n3527);
  assign n3529 = n1362 | n2840;
  assign n3530 = n1275 | n1362;
  assign n3531 = (n1232 & n3529) | (n1232 & n3530) | (n3529 & n3530);
  assign n1365 = ~n3528 & n3531;
  assign n1366 = x21 & x39;
  assign n1367 = n1365 & n1366;
  assign n1368 = n1365 | n1366;
  assign n1369 = ~n1367 & n1368;
  assign n1370 = n3515 & n1369;
  assign n1371 = n3515 | n1369;
  assign n1372 = ~n1370 & n1371;
  assign n1373 = x20 & x40;
  assign n1374 = n1372 & n1373;
  assign n1375 = n1372 | n1373;
  assign n1376 = ~n1374 & n1375;
  assign n1377 = n1315 & n1376;
  assign n1378 = n1315 | n1376;
  assign n1379 = ~n1377 & n1378;
  assign n1380 = x19 & x41;
  assign n1381 = n1379 & n1380;
  assign n1382 = n1379 | n1380;
  assign n1383 = ~n1381 & n1382;
  assign n1384 = n2839 & n1383;
  assign n1385 = n2839 | n1383;
  assign n1386 = ~n1384 & n1385;
  assign n1387 = x18 & x42;
  assign n1388 = n1386 & n1387;
  assign n1389 = n1386 | n1387;
  assign n1390 = ~n1388 & n1389;
  assign n1391 = n2837 & n1390;
  assign n1392 = n2837 | n1390;
  assign n1393 = ~n1391 & n1392;
  assign n1394 = x17 & x43;
  assign n1395 = n1393 & n1394;
  assign n1396 = n1393 | n1394;
  assign n1397 = ~n1395 & n1396;
  assign n1398 = n1310 & n1397;
  assign n1399 = n1310 | n1397;
  assign n1400 = ~n1398 & n1399;
  assign n1401 = x16 & x44;
  assign n1402 = n1400 & n1401;
  assign n1403 = n1400 | n1401;
  assign n1404 = ~n1402 & n1403;
  assign n3905 = n1309 | n1394;
  assign n3906 = (n1308 & n1394) | (n1308 & n3905) | (n1394 & n3905);
  assign n3533 = (n1310 & n1393) | (n1310 & n3906) | (n1393 & n3906);
  assign n2876 = (n1395 & n1397) | (n1395 & n3533) | (n1397 & n3533);
  assign n2877 = n1388 | n2837;
  assign n2878 = (n1388 & n1390) | (n1388 & n2877) | (n1390 & n2877);
  assign n2879 = n1381 | n2839;
  assign n2880 = (n1381 & n1383) | (n1381 & n2879) | (n1383 & n2879);
  assign n3534 = n1374 | n1376;
  assign n3535 = (n1315 & n1374) | (n1315 & n3534) | (n1374 & n3534);
  assign n2881 = n1367 | n1369;
  assign n2882 = (n3515 & n1367) | (n3515 & n2881) | (n1367 & n2881);
  assign n2841 = (n1232 & n1275) | (n1232 & n2840) | (n1275 & n2840);
  assign n2886 = n1339 | n1341;
  assign n3536 = n1254 | n1339;
  assign n3537 = (n1339 & n1341) | (n1339 & n3536) | (n1341 & n3536);
  assign n3538 = (n2826 & n2886) | (n2826 & n3537) | (n2886 & n3537);
  assign n3539 = (n1256 & n2886) | (n1256 & n3537) | (n2886 & n3537);
  assign n3540 = (n2805 & n3538) | (n2805 & n3539) | (n3538 & n3539);
  assign n1416 = x29 & x32;
  assign n1417 = x28 & x33;
  assign n1418 = n1416 & n1417;
  assign n1419 = n1416 | n1417;
  assign n1420 = ~n1418 & n1419;
  assign n3545 = n1325 | n1327;
  assign n3907 = n1420 & n3545;
  assign n3908 = n1325 & n1420;
  assign n3909 = (n3517 & n3907) | (n3517 & n3908) | (n3907 & n3908);
  assign n3547 = (n1325 & n3519) | (n1325 & n3545) | (n3519 & n3545);
  assign n3549 = n1420 & n3547;
  assign n3550 = (n3484 & n3909) | (n3484 & n3549) | (n3909 & n3549);
  assign n3910 = n1420 | n3545;
  assign n3911 = n1325 | n1420;
  assign n3912 = (n3517 & n3910) | (n3517 & n3911) | (n3910 & n3911);
  assign n3552 = n1420 | n3547;
  assign n3553 = (n3484 & n3912) | (n3484 & n3552) | (n3912 & n3552);
  assign n1423 = ~n3550 & n3553;
  assign n1424 = x27 & x34;
  assign n1425 = n1423 & n1424;
  assign n1426 = n1423 | n1424;
  assign n1427 = ~n1425 & n1426;
  assign n3541 = n1332 | n1334;
  assign n3542 = (n1332 & n2844) | (n1332 & n3541) | (n2844 & n3541);
  assign n3554 = n1427 & n3542;
  assign n3543 = n1247 | n1332;
  assign n3544 = (n1332 & n1334) | (n1332 & n3543) | (n1334 & n3543);
  assign n3555 = n1427 & n3544;
  assign n3556 = (n3501 & n3554) | (n3501 & n3555) | (n3554 & n3555);
  assign n3557 = n1427 | n3542;
  assign n3558 = n1427 | n3544;
  assign n3559 = (n3501 & n3557) | (n3501 & n3558) | (n3557 & n3558);
  assign n1430 = ~n3556 & n3559;
  assign n1431 = x26 & x35;
  assign n1432 = n1430 & n1431;
  assign n1433 = n1430 | n1431;
  assign n1434 = ~n1432 & n1433;
  assign n1435 = n3540 & n1434;
  assign n1436 = n3540 | n1434;
  assign n1437 = ~n1435 & n1436;
  assign n1438 = x25 & x36;
  assign n1439 = n1437 & n1438;
  assign n1440 = n1437 | n1438;
  assign n1441 = ~n1439 & n1440;
  assign n2894 = n1346 & n1441;
  assign n2895 = (n1441 & n2866) | (n1441 & n2894) | (n2866 & n2894);
  assign n2896 = n1346 | n1441;
  assign n2897 = n2866 | n2896;
  assign n1444 = ~n2895 & n2897;
  assign n1445 = x24 & x37;
  assign n1446 = n1444 & n1445;
  assign n1447 = n1444 | n1445;
  assign n1448 = ~n1446 & n1447;
  assign n2898 = n1353 & n1448;
  assign n2899 = (n1448 & n2871) | (n1448 & n2898) | (n2871 & n2898);
  assign n2900 = n1353 | n1448;
  assign n2901 = n2871 | n2900;
  assign n1451 = ~n2899 & n2901;
  assign n1452 = x23 & x38;
  assign n1453 = n1451 & n1452;
  assign n1454 = n1451 | n1452;
  assign n1455 = ~n1453 & n1454;
  assign n2883 = n1360 | n1362;
  assign n2902 = n1455 & n2883;
  assign n2903 = n1360 & n1455;
  assign n2904 = (n2841 & n2902) | (n2841 & n2903) | (n2902 & n2903);
  assign n2905 = n1455 | n2883;
  assign n2906 = n1360 | n1455;
  assign n2907 = (n2841 & n2905) | (n2841 & n2906) | (n2905 & n2906);
  assign n1458 = ~n2904 & n2907;
  assign n1459 = x22 & x39;
  assign n1460 = n1458 & n1459;
  assign n1461 = n1458 | n1459;
  assign n1462 = ~n1460 & n1461;
  assign n1463 = n2882 & n1462;
  assign n1464 = n2882 | n1462;
  assign n1465 = ~n1463 & n1464;
  assign n1466 = x21 & x40;
  assign n1467 = n1465 & n1466;
  assign n1468 = n1465 | n1466;
  assign n1469 = ~n1467 & n1468;
  assign n1470 = n3535 & n1469;
  assign n1471 = n3535 | n1469;
  assign n1472 = ~n1470 & n1471;
  assign n1473 = x20 & x41;
  assign n1474 = n1472 & n1473;
  assign n1475 = n1472 | n1473;
  assign n1476 = ~n1474 & n1475;
  assign n1477 = n2880 & n1476;
  assign n1478 = n2880 | n1476;
  assign n1479 = ~n1477 & n1478;
  assign n1480 = x19 & x42;
  assign n1481 = n1479 & n1480;
  assign n1482 = n1479 | n1480;
  assign n1483 = ~n1481 & n1482;
  assign n1484 = n2878 & n1483;
  assign n1485 = n2878 | n1483;
  assign n1486 = ~n1484 & n1485;
  assign n1487 = x18 & x43;
  assign n1488 = n1486 & n1487;
  assign n1489 = n1486 | n1487;
  assign n1490 = ~n1488 & n1489;
  assign n1491 = n2876 & n1490;
  assign n1492 = n2876 | n1490;
  assign n1493 = ~n1491 & n1492;
  assign n1494 = x17 & x44;
  assign n1495 = n1493 & n1494;
  assign n1496 = n1493 | n1494;
  assign n1497 = ~n1495 & n1496;
  assign n1498 = n1402 & n1497;
  assign n1499 = n1402 | n1497;
  assign n1500 = ~n1498 & n1499;
  assign n1501 = x16 & x45;
  assign n1502 = n1500 & n1501;
  assign n1503 = n1500 | n1501;
  assign n1504 = ~n1502 & n1503;
  assign n2908 = n1402 | n1495;
  assign n2909 = (n1495 & n1497) | (n1495 & n2908) | (n1497 & n2908);
  assign n2910 = n1488 | n2876;
  assign n2911 = (n1488 & n1490) | (n1488 & n2910) | (n1490 & n2910);
  assign n2912 = n1481 | n2878;
  assign n2913 = (n1481 & n1483) | (n1481 & n2912) | (n1483 & n2912);
  assign n2914 = n1474 | n2880;
  assign n2915 = (n1474 & n1476) | (n1474 & n2914) | (n1476 & n2914);
  assign n2916 = n1467 | n1469;
  assign n2917 = (n3535 & n1467) | (n3535 & n2916) | (n1467 & n2916);
  assign n1517 = x30 & x32;
  assign n1518 = x29 & x33;
  assign n1519 = n1517 & n1518;
  assign n1520 = n1517 | n1518;
  assign n1521 = ~n1519 & n1520;
  assign n2924 = n1418 | n1420;
  assign n2926 = n1521 & n2924;
  assign n2927 = n1418 & n1521;
  assign n3546 = (n1325 & n3517) | (n1325 & n3545) | (n3517 & n3545);
  assign n3560 = (n2926 & n2927) | (n2926 & n3546) | (n2927 & n3546);
  assign n3561 = (n2926 & n2927) | (n2926 & n3547) | (n2927 & n3547);
  assign n3562 = (n3484 & n3560) | (n3484 & n3561) | (n3560 & n3561);
  assign n2929 = n1521 | n2924;
  assign n2930 = n1418 | n1521;
  assign n3563 = (n2929 & n2930) | (n2929 & n3546) | (n2930 & n3546);
  assign n3564 = (n2929 & n2930) | (n2929 & n3547) | (n2930 & n3547);
  assign n3565 = (n3484 & n3563) | (n3484 & n3564) | (n3563 & n3564);
  assign n1524 = ~n3562 & n3565;
  assign n1525 = x28 & x34;
  assign n1526 = n1524 & n1525;
  assign n1527 = n1524 | n1525;
  assign n1528 = ~n1526 & n1527;
  assign n2922 = n1425 | n1427;
  assign n2932 = n1528 & n2922;
  assign n2933 = n1425 & n1528;
  assign n3566 = (n2932 & n2933) | (n2932 & n3542) | (n2933 & n3542);
  assign n3567 = (n2932 & n2933) | (n2932 & n3544) | (n2933 & n3544);
  assign n3568 = (n3501 & n3566) | (n3501 & n3567) | (n3566 & n3567);
  assign n2935 = n1528 | n2922;
  assign n2936 = n1425 | n1528;
  assign n3569 = (n2935 & n2936) | (n2935 & n3542) | (n2936 & n3542);
  assign n3570 = (n2935 & n2936) | (n2935 & n3544) | (n2936 & n3544);
  assign n3571 = (n3501 & n3569) | (n3501 & n3570) | (n3569 & n3570);
  assign n1531 = ~n3568 & n3571;
  assign n1532 = x27 & x35;
  assign n1533 = n1531 & n1532;
  assign n1534 = n1531 | n1532;
  assign n1535 = ~n1533 & n1534;
  assign n2920 = n1432 | n1434;
  assign n2938 = n1535 & n2920;
  assign n2939 = n1432 & n1535;
  assign n2940 = (n3540 & n2938) | (n3540 & n2939) | (n2938 & n2939);
  assign n2941 = n1535 | n2920;
  assign n2942 = n1432 | n1535;
  assign n2943 = (n3540 & n2941) | (n3540 & n2942) | (n2941 & n2942);
  assign n1538 = ~n2940 & n2943;
  assign n1539 = x26 & x36;
  assign n1540 = n1538 & n1539;
  assign n1541 = n1538 | n1539;
  assign n1542 = ~n1540 & n1541;
  assign n2944 = n1439 & n1542;
  assign n3572 = (n1542 & n2894) | (n1542 & n2944) | (n2894 & n2944);
  assign n3573 = (n1441 & n1542) | (n1441 & n2944) | (n1542 & n2944);
  assign n3574 = (n2866 & n3572) | (n2866 & n3573) | (n3572 & n3573);
  assign n2946 = n1439 | n1542;
  assign n3575 = n2894 | n2946;
  assign n3576 = n1441 | n2946;
  assign n3577 = (n2866 & n3575) | (n2866 & n3576) | (n3575 & n3576);
  assign n1545 = ~n3574 & n3577;
  assign n1546 = x25 & x37;
  assign n1547 = n1545 & n1546;
  assign n1548 = n1545 | n1546;
  assign n1549 = ~n1547 & n1548;
  assign n2948 = n1446 & n1549;
  assign n2949 = (n1549 & n2899) | (n1549 & n2948) | (n2899 & n2948);
  assign n2950 = n1446 | n1549;
  assign n2951 = n2899 | n2950;
  assign n1552 = ~n2949 & n2951;
  assign n1553 = x24 & x38;
  assign n1554 = n1552 & n1553;
  assign n1555 = n1552 | n1553;
  assign n1556 = ~n1554 & n1555;
  assign n2952 = n1453 & n1556;
  assign n2953 = (n1556 & n2904) | (n1556 & n2952) | (n2904 & n2952);
  assign n2954 = n1453 | n1556;
  assign n2955 = n2904 | n2954;
  assign n1559 = ~n2953 & n2955;
  assign n1560 = x23 & x39;
  assign n1561 = n1559 & n1560;
  assign n1562 = n1559 | n1560;
  assign n1563 = ~n1561 & n1562;
  assign n2918 = n1460 | n1462;
  assign n2956 = n1563 & n2918;
  assign n2957 = n1460 & n1563;
  assign n2958 = (n2882 & n2956) | (n2882 & n2957) | (n2956 & n2957);
  assign n2959 = n1563 | n2918;
  assign n2960 = n1460 | n1563;
  assign n2961 = (n2882 & n2959) | (n2882 & n2960) | (n2959 & n2960);
  assign n1566 = ~n2958 & n2961;
  assign n1567 = x22 & x40;
  assign n1568 = n1566 & n1567;
  assign n1569 = n1566 | n1567;
  assign n1570 = ~n1568 & n1569;
  assign n1571 = n2917 & n1570;
  assign n1572 = n2917 | n1570;
  assign n1573 = ~n1571 & n1572;
  assign n1574 = x21 & x41;
  assign n1575 = n1573 & n1574;
  assign n1576 = n1573 | n1574;
  assign n1577 = ~n1575 & n1576;
  assign n1578 = n2915 & n1577;
  assign n1579 = n2915 | n1577;
  assign n1580 = ~n1578 & n1579;
  assign n1581 = x20 & x42;
  assign n1582 = n1580 & n1581;
  assign n1583 = n1580 | n1581;
  assign n1584 = ~n1582 & n1583;
  assign n1585 = n2913 & n1584;
  assign n1586 = n2913 | n1584;
  assign n1587 = ~n1585 & n1586;
  assign n1588 = x19 & x43;
  assign n1589 = n1587 & n1588;
  assign n1590 = n1587 | n1588;
  assign n1591 = ~n1589 & n1590;
  assign n1592 = n2911 & n1591;
  assign n1593 = n2911 | n1591;
  assign n1594 = ~n1592 & n1593;
  assign n1595 = x18 & x44;
  assign n1596 = n1594 & n1595;
  assign n1597 = n1594 | n1595;
  assign n1598 = ~n1596 & n1597;
  assign n1599 = n2909 & n1598;
  assign n1600 = n2909 | n1598;
  assign n1601 = ~n1599 & n1600;
  assign n1602 = x17 & x45;
  assign n1603 = n1601 & n1602;
  assign n1604 = n1601 | n1602;
  assign n1605 = ~n1603 & n1604;
  assign n1606 = n1502 & n1605;
  assign n1607 = n1502 | n1605;
  assign n1608 = ~n1606 & n1607;
  assign n1609 = x16 & x46;
  assign n1610 = n1608 & n1609;
  assign n1611 = n1608 | n1609;
  assign n1612 = ~n1610 & n1611;
  assign n3913 = n1501 | n1602;
  assign n3914 = (n1500 & n1602) | (n1500 & n3913) | (n1602 & n3913);
  assign n3579 = (n1502 & n1601) | (n1502 & n3914) | (n1601 & n3914);
  assign n2963 = (n1603 & n1605) | (n1603 & n3579) | (n1605 & n3579);
  assign n3580 = n1596 | n2909;
  assign n3581 = (n1596 & n1598) | (n1596 & n3580) | (n1598 & n3580);
  assign n1615 = n1589 | n1592;
  assign n1616 = n1582 | n1585;
  assign n2967 = n1540 | n1542;
  assign n3582 = n1439 | n1540;
  assign n3583 = (n1540 & n1542) | (n1540 & n3582) | (n1542 & n3582);
  assign n3584 = (n2894 & n2967) | (n2894 & n3583) | (n2967 & n3583);
  assign n3585 = (n1441 & n2967) | (n1441 & n3583) | (n2967 & n3583);
  assign n3586 = (n2866 & n3584) | (n2866 & n3585) | (n3584 & n3585);
  assign n3587 = n1526 | n1528;
  assign n3588 = (n1526 & n2922) | (n1526 & n3587) | (n2922 & n3587);
  assign n3589 = n1425 | n1526;
  assign n3590 = (n1526 & n1528) | (n1526 & n3589) | (n1528 & n3589);
  assign n3591 = (n3542 & n3588) | (n3542 & n3590) | (n3588 & n3590);
  assign n3592 = (n3544 & n3588) | (n3544 & n3590) | (n3588 & n3590);
  assign n3593 = (n3501 & n3591) | (n3501 & n3592) | (n3591 & n3592);
  assign n1626 = x31 & x32;
  assign n1627 = x30 & x33;
  assign n1628 = n1626 & n1627;
  assign n1629 = n1626 | n1627;
  assign n1630 = ~n1628 & n1629;
  assign n3594 = n1519 | n1521;
  assign n3595 = (n1519 & n2924) | (n1519 & n3594) | (n2924 & n3594);
  assign n2975 = n1630 & n3595;
  assign n3596 = n1418 | n1519;
  assign n3597 = (n1519 & n1521) | (n1519 & n3596) | (n1521 & n3596);
  assign n2976 = n1630 & n3597;
  assign n3598 = (n2975 & n2976) | (n2975 & n3546) | (n2976 & n3546);
  assign n3599 = (n2975 & n2976) | (n2975 & n3547) | (n2976 & n3547);
  assign n3600 = (n3484 & n3598) | (n3484 & n3599) | (n3598 & n3599);
  assign n2978 = n1630 | n3595;
  assign n2979 = n1630 | n3597;
  assign n3601 = (n2978 & n2979) | (n2978 & n3546) | (n2979 & n3546);
  assign n3602 = (n2978 & n2979) | (n2978 & n3547) | (n2979 & n3547);
  assign n3603 = (n3484 & n3601) | (n3484 & n3602) | (n3601 & n3602);
  assign n1633 = ~n3600 & n3603;
  assign n1634 = x29 & x34;
  assign n1635 = n1633 & n1634;
  assign n1636 = n1633 | n1634;
  assign n1637 = ~n1635 & n1636;
  assign n1638 = n3593 & n1637;
  assign n1639 = n3593 | n1637;
  assign n1640 = ~n1638 & n1639;
  assign n1641 = x28 & x35;
  assign n1642 = n1640 & n1641;
  assign n1643 = n1640 | n1641;
  assign n1644 = ~n1642 & n1643;
  assign n2981 = n1533 & n1644;
  assign n3604 = (n1644 & n2938) | (n1644 & n2981) | (n2938 & n2981);
  assign n3605 = (n1644 & n2939) | (n1644 & n2981) | (n2939 & n2981);
  assign n3606 = (n3540 & n3604) | (n3540 & n3605) | (n3604 & n3605);
  assign n2983 = n1533 | n1644;
  assign n3607 = n2938 | n2983;
  assign n3608 = n2939 | n2983;
  assign n3609 = (n3540 & n3607) | (n3540 & n3608) | (n3607 & n3608);
  assign n1647 = ~n3606 & n3609;
  assign n1648 = x27 & x36;
  assign n1649 = n1647 & n1648;
  assign n1650 = n1647 | n1648;
  assign n1651 = ~n1649 & n1650;
  assign n1652 = n3586 & n1651;
  assign n1653 = n3586 | n1651;
  assign n1654 = ~n1652 & n1653;
  assign n1655 = x26 & x37;
  assign n1656 = n1654 & n1655;
  assign n1657 = n1654 | n1655;
  assign n1658 = ~n1656 & n1657;
  assign n2985 = n1547 & n1658;
  assign n2986 = (n1658 & n2949) | (n1658 & n2985) | (n2949 & n2985);
  assign n2987 = n1547 | n1658;
  assign n2988 = n2949 | n2987;
  assign n1661 = ~n2986 & n2988;
  assign n1662 = x25 & x38;
  assign n1663 = n1661 & n1662;
  assign n1664 = n1661 | n1662;
  assign n1665 = ~n1663 & n1664;
  assign n2989 = n1554 & n1665;
  assign n2990 = (n1665 & n2953) | (n1665 & n2989) | (n2953 & n2989);
  assign n2991 = n1554 | n1665;
  assign n2992 = n2953 | n2991;
  assign n1668 = ~n2990 & n2992;
  assign n1669 = x24 & x39;
  assign n1670 = n1668 & n1669;
  assign n1671 = n1668 | n1669;
  assign n1672 = ~n1670 & n1671;
  assign n2993 = n1561 & n1672;
  assign n2994 = (n1672 & n2958) | (n1672 & n2993) | (n2958 & n2993);
  assign n2995 = n1561 | n1672;
  assign n2996 = n2958 | n2995;
  assign n1675 = ~n2994 & n2996;
  assign n1676 = x23 & x40;
  assign n1677 = n1675 & n1676;
  assign n1678 = n1675 | n1676;
  assign n1679 = ~n1677 & n1678;
  assign n2964 = n1568 | n1570;
  assign n2997 = n1679 & n2964;
  assign n2998 = n1568 & n1679;
  assign n2999 = (n2917 & n2997) | (n2917 & n2998) | (n2997 & n2998);
  assign n3000 = n1679 | n2964;
  assign n3001 = n1568 | n1679;
  assign n3002 = (n2917 & n3000) | (n2917 & n3001) | (n3000 & n3001);
  assign n1682 = ~n2999 & n3002;
  assign n1683 = x22 & x41;
  assign n1684 = n1682 & n1683;
  assign n1685 = n1682 | n1683;
  assign n1686 = ~n1684 & n1685;
  assign n3003 = n1575 & n1686;
  assign n3004 = (n1578 & n1686) | (n1578 & n3003) | (n1686 & n3003);
  assign n3005 = n1575 | n1686;
  assign n3006 = n1578 | n3005;
  assign n1689 = ~n3004 & n3006;
  assign n1690 = x21 & x42;
  assign n1691 = n1689 & n1690;
  assign n1692 = n1689 | n1690;
  assign n1693 = ~n1691 & n1692;
  assign n1694 = n1616 & n1693;
  assign n1695 = n1616 | n1693;
  assign n1696 = ~n1694 & n1695;
  assign n1697 = x20 & x43;
  assign n1698 = n1696 & n1697;
  assign n1699 = n1696 | n1697;
  assign n1700 = ~n1698 & n1699;
  assign n1701 = n1615 & n1700;
  assign n1702 = n1615 | n1700;
  assign n1703 = ~n1701 & n1702;
  assign n1704 = x19 & x44;
  assign n1705 = n1703 & n1704;
  assign n1706 = n1703 | n1704;
  assign n1707 = ~n1705 & n1706;
  assign n1708 = n3581 & n1707;
  assign n1709 = n3581 | n1707;
  assign n1710 = ~n1708 & n1709;
  assign n1711 = x18 & x45;
  assign n1712 = n1710 & n1711;
  assign n1713 = n1710 | n1711;
  assign n1714 = ~n1712 & n1713;
  assign n1715 = n2963 & n1714;
  assign n1716 = n2963 | n1714;
  assign n1717 = ~n1715 & n1716;
  assign n1718 = x17 & x46;
  assign n1719 = n1717 & n1718;
  assign n1720 = n1717 | n1718;
  assign n1721 = ~n1719 & n1720;
  assign n1722 = n1610 & n1721;
  assign n1723 = n1610 | n1721;
  assign n1724 = ~n1722 & n1723;
  assign n1725 = x16 & x47;
  assign n1726 = n1724 & n1725;
  assign n1727 = n1724 | n1725;
  assign n1728 = ~n1726 & n1727;
  assign n3915 = n1609 | n1718;
  assign n3916 = (n1608 & n1718) | (n1608 & n3915) | (n1718 & n3915);
  assign n3611 = (n1610 & n1717) | (n1610 & n3916) | (n1717 & n3916);
  assign n3008 = (n1719 & n1721) | (n1719 & n3611) | (n1721 & n3611);
  assign n3009 = n1712 | n2963;
  assign n3010 = (n1712 & n1714) | (n1712 & n3009) | (n1714 & n3009);
  assign n3612 = n1705 | n3581;
  assign n3613 = (n1705 & n1707) | (n1705 & n3612) | (n1707 & n3612);
  assign n1732 = n1698 | n1701;
  assign n3011 = n1691 | n1693;
  assign n3012 = (n1616 & n1691) | (n1616 & n3011) | (n1691 & n3011);
  assign n3016 = n1642 | n1644;
  assign n3614 = n1533 | n1642;
  assign n3615 = (n1642 & n1644) | (n1642 & n3614) | (n1644 & n3614);
  assign n3616 = (n2938 & n3016) | (n2938 & n3615) | (n3016 & n3615);
  assign n3617 = (n2939 & n3016) | (n2939 & n3615) | (n3016 & n3615);
  assign n3618 = (n3540 & n3616) | (n3540 & n3617) | (n3616 & n3617);
  assign n1743 = x31 & x33;
  assign n3619 = n1628 | n1630;
  assign n3624 = (n1628 & n3597) | (n1628 & n3619) | (n3597 & n3619);
  assign n3024 = n1743 & n3624;
  assign n3622 = n1628 & n1743;
  assign n3917 = (n1630 & n1743) | (n1630 & n3622) | (n1743 & n3622);
  assign n3623 = (n3595 & n3917) | (n3595 & n3622) | (n3917 & n3622);
  assign n3625 = (n3024 & n3546) | (n3024 & n3623) | (n3546 & n3623);
  assign n3626 = (n3024 & n3547) | (n3024 & n3623) | (n3547 & n3623);
  assign n3627 = (n3484 & n3625) | (n3484 & n3626) | (n3625 & n3626);
  assign n3027 = n1743 | n3624;
  assign n3629 = n1628 | n1743;
  assign n3918 = n1630 | n3629;
  assign n3630 = (n3595 & n3918) | (n3595 & n3629) | (n3918 & n3629);
  assign n3631 = (n3027 & n3546) | (n3027 & n3630) | (n3546 & n3630);
  assign n3632 = (n3027 & n3547) | (n3027 & n3630) | (n3547 & n3630);
  assign n3633 = (n3484 & n3631) | (n3484 & n3632) | (n3631 & n3632);
  assign n1746 = ~n3627 & n3633;
  assign n1747 = x30 & x34;
  assign n1748 = n1746 & n1747;
  assign n1749 = n1746 | n1747;
  assign n1750 = ~n1748 & n1749;
  assign n3018 = n1635 | n1637;
  assign n3029 = n1750 & n3018;
  assign n3030 = n1635 & n1750;
  assign n3031 = (n3593 & n3029) | (n3593 & n3030) | (n3029 & n3030);
  assign n3032 = n1750 | n3018;
  assign n3033 = n1635 | n1750;
  assign n3034 = (n3593 & n3032) | (n3593 & n3033) | (n3032 & n3033);
  assign n1753 = ~n3031 & n3034;
  assign n1754 = x29 & x35;
  assign n1755 = n1753 & n1754;
  assign n1756 = n1753 | n1754;
  assign n1757 = ~n1755 & n1756;
  assign n1758 = n3618 & n1757;
  assign n1759 = n3618 | n1757;
  assign n1760 = ~n1758 & n1759;
  assign n1761 = x28 & x36;
  assign n1762 = n1760 & n1761;
  assign n1763 = n1760 | n1761;
  assign n1764 = ~n1762 & n1763;
  assign n3013 = n1649 | n1651;
  assign n3035 = n1764 & n3013;
  assign n3036 = n1649 & n1764;
  assign n3037 = (n3586 & n3035) | (n3586 & n3036) | (n3035 & n3036);
  assign n3038 = n1764 | n3013;
  assign n3039 = n1649 | n1764;
  assign n3040 = (n3586 & n3038) | (n3586 & n3039) | (n3038 & n3039);
  assign n1767 = ~n3037 & n3040;
  assign n1768 = x27 & x37;
  assign n1769 = n1767 & n1768;
  assign n1770 = n1767 | n1768;
  assign n1771 = ~n1769 & n1770;
  assign n3041 = n1656 & n1771;
  assign n3634 = (n1771 & n2985) | (n1771 & n3041) | (n2985 & n3041);
  assign n3635 = (n1658 & n1771) | (n1658 & n3041) | (n1771 & n3041);
  assign n3636 = (n2949 & n3634) | (n2949 & n3635) | (n3634 & n3635);
  assign n3043 = n1656 | n1771;
  assign n3637 = n2985 | n3043;
  assign n3638 = n1658 | n3043;
  assign n3639 = (n2949 & n3637) | (n2949 & n3638) | (n3637 & n3638);
  assign n1774 = ~n3636 & n3639;
  assign n1775 = x26 & x38;
  assign n1776 = n1774 & n1775;
  assign n1777 = n1774 | n1775;
  assign n1778 = ~n1776 & n1777;
  assign n3045 = n1663 & n1778;
  assign n3046 = (n1778 & n2990) | (n1778 & n3045) | (n2990 & n3045);
  assign n3047 = n1663 | n1778;
  assign n3048 = n2990 | n3047;
  assign n1781 = ~n3046 & n3048;
  assign n1782 = x25 & x39;
  assign n1783 = n1781 & n1782;
  assign n1784 = n1781 | n1782;
  assign n1785 = ~n1783 & n1784;
  assign n3049 = n1670 & n1785;
  assign n3050 = (n1785 & n2994) | (n1785 & n3049) | (n2994 & n3049);
  assign n3051 = n1670 | n1785;
  assign n3052 = n2994 | n3051;
  assign n1788 = ~n3050 & n3052;
  assign n1789 = x24 & x40;
  assign n1790 = n1788 & n1789;
  assign n1791 = n1788 | n1789;
  assign n1792 = ~n1790 & n1791;
  assign n3053 = n1677 & n1792;
  assign n3054 = (n1792 & n2999) | (n1792 & n3053) | (n2999 & n3053);
  assign n3055 = n1677 | n1792;
  assign n3056 = n2999 | n3055;
  assign n1795 = ~n3054 & n3056;
  assign n1796 = x23 & x41;
  assign n1797 = n1795 & n1796;
  assign n1798 = n1795 | n1796;
  assign n1799 = ~n1797 & n1798;
  assign n3057 = n1684 & n1799;
  assign n3058 = (n1799 & n3004) | (n1799 & n3057) | (n3004 & n3057);
  assign n3059 = n1684 | n1799;
  assign n3060 = n3004 | n3059;
  assign n1802 = ~n3058 & n3060;
  assign n1803 = x22 & x42;
  assign n1804 = n1802 & n1803;
  assign n1805 = n1802 | n1803;
  assign n1806 = ~n1804 & n1805;
  assign n1807 = n3012 & n1806;
  assign n1808 = n3012 | n1806;
  assign n1809 = ~n1807 & n1808;
  assign n1810 = x21 & x43;
  assign n1811 = n1809 & n1810;
  assign n1812 = n1809 | n1810;
  assign n1813 = ~n1811 & n1812;
  assign n1814 = n1732 & n1813;
  assign n1815 = n1732 | n1813;
  assign n1816 = ~n1814 & n1815;
  assign n1817 = x20 & x44;
  assign n1818 = n1816 & n1817;
  assign n1819 = n1816 | n1817;
  assign n1820 = ~n1818 & n1819;
  assign n1821 = n3613 & n1820;
  assign n1822 = n3613 | n1820;
  assign n1823 = ~n1821 & n1822;
  assign n1824 = x19 & x45;
  assign n1825 = n1823 & n1824;
  assign n1826 = n1823 | n1824;
  assign n1827 = ~n1825 & n1826;
  assign n1828 = n3010 & n1827;
  assign n1829 = n3010 | n1827;
  assign n1830 = ~n1828 & n1829;
  assign n1831 = x18 & x46;
  assign n1832 = n1830 & n1831;
  assign n1833 = n1830 | n1831;
  assign n1834 = ~n1832 & n1833;
  assign n1835 = n3008 & n1834;
  assign n1836 = n3008 | n1834;
  assign n1837 = ~n1835 & n1836;
  assign n1838 = x17 & x47;
  assign n1839 = n1837 & n1838;
  assign n1840 = n1837 | n1838;
  assign n1841 = ~n1839 & n1840;
  assign n1842 = n1726 & n1841;
  assign n1843 = n1726 | n1841;
  assign n1844 = ~n1842 & n1843;
  assign n3919 = n1725 | n1838;
  assign n3920 = (n1724 & n1838) | (n1724 & n3919) | (n1838 & n3919);
  assign n3641 = (n1726 & n1837) | (n1726 & n3920) | (n1837 & n3920);
  assign n3062 = (n1839 & n1841) | (n1839 & n3641) | (n1841 & n3641);
  assign n3063 = n1832 | n3008;
  assign n3064 = (n1832 & n1834) | (n1832 & n3063) | (n1834 & n3063);
  assign n3065 = n1825 | n3010;
  assign n3066 = (n1825 & n1827) | (n1825 & n3065) | (n1827 & n3065);
  assign n3642 = n1818 | n3613;
  assign n3643 = (n1818 & n1820) | (n1818 & n3642) | (n1820 & n3642);
  assign n3067 = n1811 | n1813;
  assign n3068 = (n1732 & n1811) | (n1732 & n3067) | (n1811 & n3067);
  assign n3069 = n1804 | n1806;
  assign n3070 = (n1804 & n3012) | (n1804 & n3069) | (n3012 & n3069);
  assign n3072 = n1769 | n1771;
  assign n3644 = n1656 | n1769;
  assign n3645 = (n1769 & n1771) | (n1769 & n3644) | (n1771 & n3644);
  assign n3646 = (n2985 & n3072) | (n2985 & n3645) | (n3072 & n3645);
  assign n3647 = (n1658 & n3072) | (n1658 & n3645) | (n3072 & n3645);
  assign n3648 = (n2949 & n3646) | (n2949 & n3647) | (n3646 & n3647);
  assign n1859 = x31 & x34;
  assign n1860 = n3627 & n1859;
  assign n1861 = n3627 | n1859;
  assign n1862 = ~n1860 & n1861;
  assign n3649 = n1748 | n1750;
  assign n3650 = (n1748 & n3018) | (n1748 & n3649) | (n3018 & n3649);
  assign n3079 = n1862 & n3650;
  assign n3651 = n1635 | n1748;
  assign n3652 = (n1748 & n1750) | (n1748 & n3651) | (n1750 & n3651);
  assign n3080 = n1862 & n3652;
  assign n3081 = (n3593 & n3079) | (n3593 & n3080) | (n3079 & n3080);
  assign n3082 = n1862 | n3650;
  assign n3083 = n1862 | n3652;
  assign n3084 = (n3593 & n3082) | (n3593 & n3083) | (n3082 & n3083);
  assign n1865 = ~n3081 & n3084;
  assign n1866 = x30 & x35;
  assign n1867 = n1865 & n1866;
  assign n1868 = n1865 | n1866;
  assign n1869 = ~n1867 & n1868;
  assign n3074 = n1755 | n1757;
  assign n3085 = n1869 & n3074;
  assign n3086 = n1755 & n1869;
  assign n3087 = (n3618 & n3085) | (n3618 & n3086) | (n3085 & n3086);
  assign n3088 = n1869 | n3074;
  assign n3089 = n1755 | n1869;
  assign n3090 = (n3618 & n3088) | (n3618 & n3089) | (n3088 & n3089);
  assign n1872 = ~n3087 & n3090;
  assign n1873 = x29 & x36;
  assign n1874 = n1872 & n1873;
  assign n1875 = n1872 | n1873;
  assign n1876 = ~n1874 & n1875;
  assign n3091 = n1762 & n1876;
  assign n3653 = (n1876 & n3036) | (n1876 & n3091) | (n3036 & n3091);
  assign n3654 = (n1876 & n3035) | (n1876 & n3091) | (n3035 & n3091);
  assign n3655 = (n3586 & n3653) | (n3586 & n3654) | (n3653 & n3654);
  assign n3093 = n1762 | n1876;
  assign n3656 = n3036 | n3093;
  assign n3657 = n3035 | n3093;
  assign n3658 = (n3586 & n3656) | (n3586 & n3657) | (n3656 & n3657);
  assign n1879 = ~n3655 & n3658;
  assign n1880 = x28 & x37;
  assign n1881 = n1879 & n1880;
  assign n1882 = n1879 | n1880;
  assign n1883 = ~n1881 & n1882;
  assign n1884 = n3648 & n1883;
  assign n1885 = n3648 | n1883;
  assign n1886 = ~n1884 & n1885;
  assign n1887 = x27 & x38;
  assign n1888 = n1886 & n1887;
  assign n1889 = n1886 | n1887;
  assign n1890 = ~n1888 & n1889;
  assign n3095 = n1776 & n1890;
  assign n3096 = (n1890 & n3046) | (n1890 & n3095) | (n3046 & n3095);
  assign n3097 = n1776 | n1890;
  assign n3098 = n3046 | n3097;
  assign n1893 = ~n3096 & n3098;
  assign n1894 = x26 & x39;
  assign n1895 = n1893 & n1894;
  assign n1896 = n1893 | n1894;
  assign n1897 = ~n1895 & n1896;
  assign n3099 = n1783 & n1897;
  assign n3100 = (n1897 & n3050) | (n1897 & n3099) | (n3050 & n3099);
  assign n3101 = n1783 | n1897;
  assign n3102 = n3050 | n3101;
  assign n1900 = ~n3100 & n3102;
  assign n1901 = x25 & x40;
  assign n1902 = n1900 & n1901;
  assign n1903 = n1900 | n1901;
  assign n1904 = ~n1902 & n1903;
  assign n3103 = n1790 & n1904;
  assign n3104 = (n1904 & n3054) | (n1904 & n3103) | (n3054 & n3103);
  assign n3105 = n1790 | n1904;
  assign n3106 = n3054 | n3105;
  assign n1907 = ~n3104 & n3106;
  assign n1908 = x24 & x41;
  assign n1909 = n1907 & n1908;
  assign n1910 = n1907 | n1908;
  assign n1911 = ~n1909 & n1910;
  assign n3107 = n1797 & n1911;
  assign n3108 = (n1911 & n3058) | (n1911 & n3107) | (n3058 & n3107);
  assign n3109 = n1797 | n1911;
  assign n3110 = n3058 | n3109;
  assign n1914 = ~n3108 & n3110;
  assign n1915 = x23 & x42;
  assign n1916 = n1914 & n1915;
  assign n1917 = n1914 | n1915;
  assign n1918 = ~n1916 & n1917;
  assign n1919 = n3070 & n1918;
  assign n1920 = n3070 | n1918;
  assign n1921 = ~n1919 & n1920;
  assign n1922 = x22 & x43;
  assign n1923 = n1921 & n1922;
  assign n1924 = n1921 | n1922;
  assign n1925 = ~n1923 & n1924;
  assign n1926 = n3068 & n1925;
  assign n1927 = n3068 | n1925;
  assign n1928 = ~n1926 & n1927;
  assign n1929 = x21 & x44;
  assign n1930 = n1928 & n1929;
  assign n1931 = n1928 | n1929;
  assign n1932 = ~n1930 & n1931;
  assign n1933 = n3643 & n1932;
  assign n1934 = n3643 | n1932;
  assign n1935 = ~n1933 & n1934;
  assign n1936 = x20 & x45;
  assign n1937 = n1935 & n1936;
  assign n1938 = n1935 | n1936;
  assign n1939 = ~n1937 & n1938;
  assign n1940 = n3066 & n1939;
  assign n1941 = n3066 | n1939;
  assign n1942 = ~n1940 & n1941;
  assign n1943 = x19 & x46;
  assign n1944 = n1942 & n1943;
  assign n1945 = n1942 | n1943;
  assign n1946 = ~n1944 & n1945;
  assign n1947 = n3064 & n1946;
  assign n1948 = n3064 | n1946;
  assign n1949 = ~n1947 & n1948;
  assign n1950 = x18 & x47;
  assign n1951 = n1949 & n1950;
  assign n1952 = n1949 | n1950;
  assign n1953 = ~n1951 & n1952;
  assign n1954 = n3062 & n1953;
  assign n1955 = n3062 | n1953;
  assign n1956 = ~n1954 & n1955;
  assign n3111 = n1951 | n3062;
  assign n3112 = (n1951 & n1953) | (n1951 & n3111) | (n1953 & n3111);
  assign n3113 = n1944 | n3064;
  assign n3114 = (n1944 & n1946) | (n1944 & n3113) | (n1946 & n3113);
  assign n3115 = n1937 | n3066;
  assign n3116 = (n1937 & n1939) | (n1937 & n3115) | (n1939 & n3115);
  assign n3117 = n1930 | n1932;
  assign n3118 = (n3643 & n1930) | (n3643 & n3117) | (n1930 & n3117);
  assign n3119 = n1923 | n1925;
  assign n3120 = (n1923 & n3068) | (n1923 & n3119) | (n3068 & n3119);
  assign n3121 = n1916 | n1918;
  assign n3122 = (n1916 & n3070) | (n1916 & n3121) | (n3070 & n3121);
  assign n3126 = n1874 | n1876;
  assign n3659 = n1762 | n1874;
  assign n3660 = (n1874 & n1876) | (n1874 & n3659) | (n1876 & n3659);
  assign n3661 = (n3036 & n3126) | (n3036 & n3660) | (n3126 & n3660);
  assign n3662 = (n3035 & n3126) | (n3035 & n3660) | (n3126 & n3660);
  assign n3663 = (n3586 & n3661) | (n3586 & n3662) | (n3661 & n3662);
  assign n1971 = x31 & x35;
  assign n3668 = n1859 & n1971;
  assign n3669 = n3627 & n3668;
  assign n3921 = (n1862 & n1971) | (n1862 & n3669) | (n1971 & n3669);
  assign n4042 = n1971 & n3668;
  assign n4043 = n3627 & n4042;
  assign n3923 = (n3650 & n3921) | (n3650 & n4043) | (n3921 & n4043);
  assign n3924 = (n3652 & n3921) | (n3652 & n4043) | (n3921 & n4043);
  assign n3672 = (n3593 & n3923) | (n3593 & n3924) | (n3923 & n3924);
  assign n3673 = n1859 | n1971;
  assign n3674 = (n1971 & n3627) | (n1971 & n3673) | (n3627 & n3673);
  assign n3925 = n1862 | n3674;
  assign n3926 = (n3650 & n3674) | (n3650 & n3925) | (n3674 & n3925);
  assign n3927 = (n3652 & n3674) | (n3652 & n3925) | (n3674 & n3925);
  assign n3677 = (n3593 & n3926) | (n3593 & n3927) | (n3926 & n3927);
  assign n1974 = ~n3672 & n3677;
  assign n3664 = n1867 | n1869;
  assign n3665 = (n1867 & n3074) | (n1867 & n3664) | (n3074 & n3664);
  assign n3678 = n1974 & n3665;
  assign n3666 = n1755 | n1867;
  assign n3667 = (n1867 & n1869) | (n1867 & n3666) | (n1869 & n3666);
  assign n3679 = n1974 & n3667;
  assign n3680 = (n3618 & n3678) | (n3618 & n3679) | (n3678 & n3679);
  assign n3681 = n1974 | n3665;
  assign n3682 = n1974 | n3667;
  assign n3683 = (n3618 & n3681) | (n3618 & n3682) | (n3681 & n3682);
  assign n1977 = ~n3680 & n3683;
  assign n1978 = x30 & x36;
  assign n1979 = n1977 & n1978;
  assign n1980 = n1977 | n1978;
  assign n1981 = ~n1979 & n1980;
  assign n1982 = n3663 & n1981;
  assign n1983 = n3663 | n1981;
  assign n1984 = ~n1982 & n1983;
  assign n1985 = x29 & x37;
  assign n1986 = n1984 & n1985;
  assign n1987 = n1984 | n1985;
  assign n1988 = ~n1986 & n1987;
  assign n3123 = n1881 | n1883;
  assign n3135 = n1988 & n3123;
  assign n3136 = n1881 & n1988;
  assign n3137 = (n3648 & n3135) | (n3648 & n3136) | (n3135 & n3136);
  assign n3138 = n1988 | n3123;
  assign n3139 = n1881 | n1988;
  assign n3140 = (n3648 & n3138) | (n3648 & n3139) | (n3138 & n3139);
  assign n1991 = ~n3137 & n3140;
  assign n1992 = x28 & x38;
  assign n1993 = n1991 & n1992;
  assign n1994 = n1991 | n1992;
  assign n1995 = ~n1993 & n1994;
  assign n3141 = n1888 & n1995;
  assign n3684 = (n1995 & n3095) | (n1995 & n3141) | (n3095 & n3141);
  assign n3685 = (n1890 & n1995) | (n1890 & n3141) | (n1995 & n3141);
  assign n3686 = (n3046 & n3684) | (n3046 & n3685) | (n3684 & n3685);
  assign n3143 = n1888 | n1995;
  assign n3687 = n3095 | n3143;
  assign n3688 = n1890 | n3143;
  assign n3689 = (n3046 & n3687) | (n3046 & n3688) | (n3687 & n3688);
  assign n1998 = ~n3686 & n3689;
  assign n1999 = x27 & x39;
  assign n2000 = n1998 & n1999;
  assign n2001 = n1998 | n1999;
  assign n2002 = ~n2000 & n2001;
  assign n3145 = n1895 & n2002;
  assign n3146 = (n2002 & n3100) | (n2002 & n3145) | (n3100 & n3145);
  assign n3147 = n1895 | n2002;
  assign n3148 = n3100 | n3147;
  assign n2005 = ~n3146 & n3148;
  assign n2006 = x26 & x40;
  assign n2007 = n2005 & n2006;
  assign n2008 = n2005 | n2006;
  assign n2009 = ~n2007 & n2008;
  assign n3149 = n1902 & n2009;
  assign n3150 = (n2009 & n3104) | (n2009 & n3149) | (n3104 & n3149);
  assign n3151 = n1902 | n2009;
  assign n3152 = n3104 | n3151;
  assign n2012 = ~n3150 & n3152;
  assign n2013 = x25 & x41;
  assign n2014 = n2012 & n2013;
  assign n2015 = n2012 | n2013;
  assign n2016 = ~n2014 & n2015;
  assign n3153 = n1909 & n2016;
  assign n3154 = (n2016 & n3108) | (n2016 & n3153) | (n3108 & n3153);
  assign n3155 = n1909 | n2016;
  assign n3156 = n3108 | n3155;
  assign n2019 = ~n3154 & n3156;
  assign n2020 = x24 & x42;
  assign n2021 = n2019 & n2020;
  assign n2022 = n2019 | n2020;
  assign n2023 = ~n2021 & n2022;
  assign n2024 = n3122 & n2023;
  assign n2025 = n3122 | n2023;
  assign n2026 = ~n2024 & n2025;
  assign n2027 = x23 & x43;
  assign n2028 = n2026 & n2027;
  assign n2029 = n2026 | n2027;
  assign n2030 = ~n2028 & n2029;
  assign n2031 = n3120 & n2030;
  assign n2032 = n3120 | n2030;
  assign n2033 = ~n2031 & n2032;
  assign n2034 = x22 & x44;
  assign n2035 = n2033 & n2034;
  assign n2036 = n2033 | n2034;
  assign n2037 = ~n2035 & n2036;
  assign n2038 = n3118 & n2037;
  assign n2039 = n3118 | n2037;
  assign n2040 = ~n2038 & n2039;
  assign n2041 = x21 & x45;
  assign n2042 = n2040 & n2041;
  assign n2043 = n2040 | n2041;
  assign n2044 = ~n2042 & n2043;
  assign n2045 = n3116 & n2044;
  assign n2046 = n3116 | n2044;
  assign n2047 = ~n2045 & n2046;
  assign n2048 = x20 & x46;
  assign n2049 = n2047 & n2048;
  assign n2050 = n2047 | n2048;
  assign n2051 = ~n2049 & n2050;
  assign n2052 = n3114 & n2051;
  assign n2053 = n3114 | n2051;
  assign n2054 = ~n2052 & n2053;
  assign n2055 = x19 & x47;
  assign n2056 = n2054 & n2055;
  assign n2057 = n2054 | n2055;
  assign n2058 = ~n2056 & n2057;
  assign n2059 = n3112 & n2058;
  assign n2060 = n3112 | n2058;
  assign n2061 = ~n2059 & n2060;
  assign n2062 = n2056 | n2059;
  assign n2063 = n2049 | n2052;
  assign n2064 = n2042 | n2045;
  assign n3157 = n2035 | n2037;
  assign n3158 = (n2035 & n3118) | (n2035 & n3157) | (n3118 & n3157);
  assign n3159 = n2028 | n2030;
  assign n3160 = (n2028 & n3120) | (n2028 & n3159) | (n3120 & n3159);
  assign n3161 = n2021 | n2023;
  assign n3162 = (n2021 & n3122) | (n2021 & n3161) | (n3122 & n3161);
  assign n3164 = n1993 | n1995;
  assign n3690 = n1888 | n1993;
  assign n3691 = (n1993 & n1995) | (n1993 & n3690) | (n1995 & n3690);
  assign n3692 = (n3095 & n3164) | (n3095 & n3691) | (n3164 & n3691);
  assign n3693 = (n1890 & n3164) | (n1890 & n3691) | (n3164 & n3691);
  assign n3694 = (n3046 & n3692) | (n3046 & n3693) | (n3692 & n3693);
  assign n2075 = x31 & x36;
  assign n4129 = n2075 & n3668;
  assign n4130 = n3627 & n4129;
  assign n4096 = n1971 & n2075;
  assign n4097 = (n1862 & n4130) | (n1862 & n4096) | (n4130 & n4096);
  assign n4131 = n3668 & n4096;
  assign n4099 = n3627 & n4131;
  assign n4046 = (n3650 & n4097) | (n3650 & n4099) | (n4097 & n4099);
  assign n4047 = (n3652 & n4097) | (n3652 & n4099) | (n4097 & n4099);
  assign n3930 = (n3593 & n4046) | (n3593 & n4047) | (n4046 & n4047);
  assign n3696 = (n1974 & n2075) | (n1974 & n3930) | (n2075 & n3930);
  assign n3697 = (n3930 & n3665) | (n3930 & n3696) | (n3665 & n3696);
  assign n3698 = (n3930 & n3667) | (n3930 & n3696) | (n3667 & n3696);
  assign n3699 = (n3618 & n3697) | (n3618 & n3698) | (n3697 & n3698);
  assign n4132 = n2075 | n3668;
  assign n4133 = (n2075 & n3627) | (n2075 & n4132) | (n3627 & n4132);
  assign n4101 = n1971 | n2075;
  assign n4102 = (n1862 & n4133) | (n1862 & n4101) | (n4133 & n4101);
  assign n4134 = (n2075 & n3668) | (n2075 & n4101) | (n3668 & n4101);
  assign n4104 = (n2075 & n3627) | (n2075 & n4134) | (n3627 & n4134);
  assign n4050 = (n3650 & n4102) | (n3650 & n4104) | (n4102 & n4104);
  assign n4051 = (n3652 & n4102) | (n3652 & n4104) | (n4102 & n4104);
  assign n3933 = (n3593 & n4050) | (n3593 & n4051) | (n4050 & n4051);
  assign n3701 = n1974 | n3933;
  assign n3702 = (n3933 & n3665) | (n3933 & n3701) | (n3665 & n3701);
  assign n3703 = (n3933 & n3667) | (n3933 & n3701) | (n3667 & n3701);
  assign n3704 = (n3618 & n3702) | (n3618 & n3703) | (n3702 & n3703);
  assign n2078 = ~n3699 & n3704;
  assign n3177 = n1979 & n2078;
  assign n3705 = (n1981 & n2078) | (n1981 & n3177) | (n2078 & n3177);
  assign n3178 = (n3663 & n3705) | (n3663 & n3177) | (n3705 & n3177);
  assign n3180 = n1979 | n2078;
  assign n3706 = n1981 | n3180;
  assign n3181 = (n3663 & n3706) | (n3663 & n3180) | (n3706 & n3180);
  assign n2081 = ~n3178 & n3181;
  assign n2082 = x30 & x37;
  assign n2083 = n2081 & n2082;
  assign n2084 = n2081 | n2082;
  assign n2085 = ~n2083 & n2084;
  assign n3182 = n1986 & n2085;
  assign n3707 = (n2085 & n3136) | (n2085 & n3182) | (n3136 & n3182);
  assign n3708 = (n2085 & n3135) | (n2085 & n3182) | (n3135 & n3182);
  assign n3709 = (n3648 & n3707) | (n3648 & n3708) | (n3707 & n3708);
  assign n3184 = n1986 | n2085;
  assign n3710 = n3136 | n3184;
  assign n3711 = n3135 | n3184;
  assign n3712 = (n3648 & n3710) | (n3648 & n3711) | (n3710 & n3711);
  assign n2088 = ~n3709 & n3712;
  assign n2089 = x29 & x38;
  assign n2090 = n2088 & n2089;
  assign n2091 = n2088 | n2089;
  assign n2092 = ~n2090 & n2091;
  assign n2093 = n3694 & n2092;
  assign n2094 = n3694 | n2092;
  assign n2095 = ~n2093 & n2094;
  assign n2096 = x28 & x39;
  assign n2097 = n2095 & n2096;
  assign n2098 = n2095 | n2096;
  assign n2099 = ~n2097 & n2098;
  assign n3186 = n2000 & n2099;
  assign n3187 = (n2099 & n3146) | (n2099 & n3186) | (n3146 & n3186);
  assign n3188 = n2000 | n2099;
  assign n3189 = n3146 | n3188;
  assign n2102 = ~n3187 & n3189;
  assign n2103 = x27 & x40;
  assign n2104 = n2102 & n2103;
  assign n2105 = n2102 | n2103;
  assign n2106 = ~n2104 & n2105;
  assign n3190 = n2007 & n2106;
  assign n3191 = (n2106 & n3150) | (n2106 & n3190) | (n3150 & n3190);
  assign n3192 = n2007 | n2106;
  assign n3193 = n3150 | n3192;
  assign n2109 = ~n3191 & n3193;
  assign n2110 = x26 & x41;
  assign n2111 = n2109 & n2110;
  assign n2112 = n2109 | n2110;
  assign n2113 = ~n2111 & n2112;
  assign n3194 = n2014 & n2113;
  assign n3195 = (n2113 & n3154) | (n2113 & n3194) | (n3154 & n3194);
  assign n3196 = n2014 | n2113;
  assign n3197 = n3154 | n3196;
  assign n2116 = ~n3195 & n3197;
  assign n2117 = x25 & x42;
  assign n2118 = n2116 & n2117;
  assign n2119 = n2116 | n2117;
  assign n2120 = ~n2118 & n2119;
  assign n2121 = n3162 & n2120;
  assign n2122 = n3162 | n2120;
  assign n2123 = ~n2121 & n2122;
  assign n2124 = x24 & x43;
  assign n2125 = n2123 & n2124;
  assign n2126 = n2123 | n2124;
  assign n2127 = ~n2125 & n2126;
  assign n2128 = n3160 & n2127;
  assign n2129 = n3160 | n2127;
  assign n2130 = ~n2128 & n2129;
  assign n2131 = x23 & x44;
  assign n2132 = n2130 & n2131;
  assign n2133 = n2130 | n2131;
  assign n2134 = ~n2132 & n2133;
  assign n2135 = n3158 & n2134;
  assign n2136 = n3158 | n2134;
  assign n2137 = ~n2135 & n2136;
  assign n2138 = x22 & x45;
  assign n2139 = n2137 & n2138;
  assign n2140 = n2137 | n2138;
  assign n2141 = ~n2139 & n2140;
  assign n2142 = n2064 & n2141;
  assign n2143 = n2064 | n2141;
  assign n2144 = ~n2142 & n2143;
  assign n2145 = x21 & x46;
  assign n2146 = n2144 & n2145;
  assign n2147 = n2144 | n2145;
  assign n2148 = ~n2146 & n2147;
  assign n2149 = n2063 & n2148;
  assign n2150 = n2063 | n2148;
  assign n2151 = ~n2149 & n2150;
  assign n2152 = x20 & x47;
  assign n2153 = n2151 & n2152;
  assign n2154 = n2151 | n2152;
  assign n2155 = ~n2153 & n2154;
  assign n2156 = n2062 & n2155;
  assign n2157 = n2062 | n2155;
  assign n2158 = ~n2156 & n2157;
  assign n2159 = n2153 | n2156;
  assign n2160 = n2146 | n2149;
  assign n3198 = n2139 | n2141;
  assign n3199 = (n2064 & n2139) | (n2064 & n3198) | (n2139 & n3198);
  assign n3200 = n2132 | n2134;
  assign n3201 = (n2132 & n3158) | (n2132 & n3200) | (n3158 & n3200);
  assign n3202 = n2125 | n2127;
  assign n3203 = (n2125 & n3160) | (n2125 & n3202) | (n3160 & n3202);
  assign n3204 = n2118 | n2120;
  assign n3205 = (n2118 & n3162) | (n2118 & n3204) | (n3162 & n3204);
  assign n3209 = n2083 | n2085;
  assign n3713 = n1986 | n2083;
  assign n3714 = (n2083 & n2085) | (n2083 & n3713) | (n2085 & n3713);
  assign n3715 = (n3136 & n3209) | (n3136 & n3714) | (n3209 & n3714);
  assign n3716 = (n3135 & n3209) | (n3135 & n3714) | (n3209 & n3714);
  assign n3717 = (n3648 & n3715) | (n3648 & n3716) | (n3715 & n3716);
  assign n2171 = x31 & x37;
  assign n3211 = n2171 & n3699;
  assign n3718 = (n2171 & n3211) | (n2171 & n3705) | (n3211 & n3705);
  assign n3934 = (n2078 & n2171) | (n2078 & n3211) | (n2171 & n3211);
  assign n4052 = n2171 & n3699;
  assign n3936 = (n1979 & n3934) | (n1979 & n4052) | (n3934 & n4052);
  assign n3720 = (n3663 & n3718) | (n3663 & n3936) | (n3718 & n3936);
  assign n3213 = n2171 | n3699;
  assign n3721 = n3213 | n3705;
  assign n3937 = n2078 | n3213;
  assign n3938 = (n1979 & n3213) | (n1979 & n3937) | (n3213 & n3937);
  assign n3723 = (n3663 & n3721) | (n3663 & n3938) | (n3721 & n3938);
  assign n2174 = ~n3720 & n3723;
  assign n2175 = n3717 & n2174;
  assign n2176 = n3717 | n2174;
  assign n2177 = ~n2175 & n2176;
  assign n2178 = x30 & x38;
  assign n2179 = n2177 & n2178;
  assign n2180 = n2177 | n2178;
  assign n2181 = ~n2179 & n2180;
  assign n3206 = n2090 | n2092;
  assign n3215 = n2181 & n3206;
  assign n3216 = n2090 & n2181;
  assign n3217 = (n3694 & n3215) | (n3694 & n3216) | (n3215 & n3216);
  assign n3218 = n2181 | n3206;
  assign n3219 = n2090 | n2181;
  assign n3220 = (n3694 & n3218) | (n3694 & n3219) | (n3218 & n3219);
  assign n2184 = ~n3217 & n3220;
  assign n2185 = x29 & x39;
  assign n2186 = n2184 & n2185;
  assign n2187 = n2184 | n2185;
  assign n2188 = ~n2186 & n2187;
  assign n3221 = n2097 & n2188;
  assign n3724 = (n2188 & n3186) | (n2188 & n3221) | (n3186 & n3221);
  assign n3725 = (n2099 & n2188) | (n2099 & n3221) | (n2188 & n3221);
  assign n3726 = (n3146 & n3724) | (n3146 & n3725) | (n3724 & n3725);
  assign n3223 = n2097 | n2188;
  assign n3727 = n3186 | n3223;
  assign n3728 = n2099 | n3223;
  assign n3729 = (n3146 & n3727) | (n3146 & n3728) | (n3727 & n3728);
  assign n2191 = ~n3726 & n3729;
  assign n2192 = x28 & x40;
  assign n2193 = n2191 & n2192;
  assign n2194 = n2191 | n2192;
  assign n2195 = ~n2193 & n2194;
  assign n3225 = n2104 & n2195;
  assign n3226 = (n2195 & n3191) | (n2195 & n3225) | (n3191 & n3225);
  assign n3227 = n2104 | n2195;
  assign n3228 = n3191 | n3227;
  assign n2198 = ~n3226 & n3228;
  assign n2199 = x27 & x41;
  assign n2200 = n2198 & n2199;
  assign n2201 = n2198 | n2199;
  assign n2202 = ~n2200 & n2201;
  assign n3229 = n2111 & n2202;
  assign n3230 = (n2202 & n3195) | (n2202 & n3229) | (n3195 & n3229);
  assign n3231 = n2111 | n2202;
  assign n3232 = n3195 | n3231;
  assign n2205 = ~n3230 & n3232;
  assign n2206 = x26 & x42;
  assign n2207 = n2205 & n2206;
  assign n2208 = n2205 | n2206;
  assign n2209 = ~n2207 & n2208;
  assign n2210 = n3205 & n2209;
  assign n2211 = n3205 | n2209;
  assign n2212 = ~n2210 & n2211;
  assign n2213 = x25 & x43;
  assign n2214 = n2212 & n2213;
  assign n2215 = n2212 | n2213;
  assign n2216 = ~n2214 & n2215;
  assign n2217 = n3203 & n2216;
  assign n2218 = n3203 | n2216;
  assign n2219 = ~n2217 & n2218;
  assign n2220 = x24 & x44;
  assign n2221 = n2219 & n2220;
  assign n2222 = n2219 | n2220;
  assign n2223 = ~n2221 & n2222;
  assign n2224 = n3201 & n2223;
  assign n2225 = n3201 | n2223;
  assign n2226 = ~n2224 & n2225;
  assign n2227 = x23 & x45;
  assign n2228 = n2226 & n2227;
  assign n2229 = n2226 | n2227;
  assign n2230 = ~n2228 & n2229;
  assign n2231 = n3199 & n2230;
  assign n2232 = n3199 | n2230;
  assign n2233 = ~n2231 & n2232;
  assign n2234 = x22 & x46;
  assign n2235 = n2233 & n2234;
  assign n2236 = n2233 | n2234;
  assign n2237 = ~n2235 & n2236;
  assign n2238 = n2160 & n2237;
  assign n2239 = n2160 | n2237;
  assign n2240 = ~n2238 & n2239;
  assign n2241 = x21 & x47;
  assign n2242 = n2240 & n2241;
  assign n2243 = n2240 | n2241;
  assign n2244 = ~n2242 & n2243;
  assign n2245 = n2159 & n2244;
  assign n2246 = n2159 | n2244;
  assign n2247 = ~n2245 & n2246;
  assign n2248 = n2242 | n2245;
  assign n3233 = n2235 | n2237;
  assign n3234 = (n2160 & n2235) | (n2160 & n3233) | (n2235 & n3233);
  assign n3235 = n2228 | n2230;
  assign n3236 = (n2228 & n3199) | (n2228 & n3235) | (n3199 & n3235);
  assign n3237 = n2221 | n2223;
  assign n3238 = (n2221 & n3201) | (n2221 & n3237) | (n3201 & n3237);
  assign n3239 = n2214 | n2216;
  assign n3240 = (n2214 & n3203) | (n2214 & n3239) | (n3203 & n3239);
  assign n3241 = n2207 | n2209;
  assign n3242 = (n2207 & n3205) | (n2207 & n3241) | (n3205 & n3241);
  assign n3244 = n2186 | n2188;
  assign n3730 = n2097 | n2186;
  assign n3731 = (n2186 & n2188) | (n2186 & n3730) | (n2188 & n3730);
  assign n3732 = (n3186 & n3244) | (n3186 & n3731) | (n3244 & n3731);
  assign n3733 = (n2099 & n3244) | (n2099 & n3731) | (n3244 & n3731);
  assign n3734 = (n3146 & n3732) | (n3146 & n3733) | (n3732 & n3733);
  assign n2259 = x31 & x38;
  assign n3942 = n2171 & n2259;
  assign n4053 = n3699 & n3942;
  assign n3943 = (n3705 & n4053) | (n3705 & n3942) | (n4053 & n3942);
  assign n3939 = n2259 & n3936;
  assign n3940 = (n3663 & n3943) | (n3663 & n3939) | (n3943 & n3939);
  assign n3736 = (n2174 & n2259) | (n2174 & n3940) | (n2259 & n3940);
  assign n3738 = n2259 & n3936;
  assign n3739 = (n3663 & n3943) | (n3663 & n3738) | (n3943 & n3738);
  assign n3250 = (n3717 & n3736) | (n3717 & n3739) | (n3736 & n3739);
  assign n3947 = n2171 | n2259;
  assign n4054 = (n2259 & n3699) | (n2259 & n3947) | (n3699 & n3947);
  assign n3948 = (n3705 & n4054) | (n3705 & n3947) | (n4054 & n3947);
  assign n3944 = n2259 | n3936;
  assign n3945 = (n3663 & n3948) | (n3663 & n3944) | (n3948 & n3944);
  assign n3741 = n2174 | n3945;
  assign n3743 = n2259 | n3936;
  assign n3744 = (n3663 & n3948) | (n3663 & n3743) | (n3948 & n3743);
  assign n3253 = (n3717 & n3741) | (n3717 & n3744) | (n3741 & n3744);
  assign n2262 = ~n3250 & n3253;
  assign n3254 = n2179 & n2262;
  assign n3745 = (n2262 & n3216) | (n2262 & n3254) | (n3216 & n3254);
  assign n3746 = (n2262 & n3215) | (n2262 & n3254) | (n3215 & n3254);
  assign n3747 = (n3694 & n3745) | (n3694 & n3746) | (n3745 & n3746);
  assign n3256 = n2179 | n2262;
  assign n3748 = n3216 | n3256;
  assign n3749 = n3215 | n3256;
  assign n3750 = (n3694 & n3748) | (n3694 & n3749) | (n3748 & n3749);
  assign n2265 = ~n3747 & n3750;
  assign n2266 = x30 & x39;
  assign n2267 = n2265 & n2266;
  assign n2268 = n2265 | n2266;
  assign n2269 = ~n2267 & n2268;
  assign n2270 = n3734 & n2269;
  assign n2271 = n3734 | n2269;
  assign n2272 = ~n2270 & n2271;
  assign n2273 = x29 & x40;
  assign n2274 = n2272 & n2273;
  assign n2275 = n2272 | n2273;
  assign n2276 = ~n2274 & n2275;
  assign n3258 = n2193 & n2276;
  assign n3259 = (n2276 & n3226) | (n2276 & n3258) | (n3226 & n3258);
  assign n3260 = n2193 | n2276;
  assign n3261 = n3226 | n3260;
  assign n2279 = ~n3259 & n3261;
  assign n2280 = x28 & x41;
  assign n2281 = n2279 & n2280;
  assign n2282 = n2279 | n2280;
  assign n2283 = ~n2281 & n2282;
  assign n3262 = n2200 & n2283;
  assign n3263 = (n2283 & n3230) | (n2283 & n3262) | (n3230 & n3262);
  assign n3264 = n2200 | n2283;
  assign n3265 = n3230 | n3264;
  assign n2286 = ~n3263 & n3265;
  assign n2287 = x27 & x42;
  assign n2288 = n2286 & n2287;
  assign n2289 = n2286 | n2287;
  assign n2290 = ~n2288 & n2289;
  assign n2291 = n3242 & n2290;
  assign n2292 = n3242 | n2290;
  assign n2293 = ~n2291 & n2292;
  assign n2294 = x26 & x43;
  assign n2295 = n2293 & n2294;
  assign n2296 = n2293 | n2294;
  assign n2297 = ~n2295 & n2296;
  assign n2298 = n3240 & n2297;
  assign n2299 = n3240 | n2297;
  assign n2300 = ~n2298 & n2299;
  assign n2301 = x25 & x44;
  assign n2302 = n2300 & n2301;
  assign n2303 = n2300 | n2301;
  assign n2304 = ~n2302 & n2303;
  assign n2305 = n3238 & n2304;
  assign n2306 = n3238 | n2304;
  assign n2307 = ~n2305 & n2306;
  assign n2308 = x24 & x45;
  assign n2309 = n2307 & n2308;
  assign n2310 = n2307 | n2308;
  assign n2311 = ~n2309 & n2310;
  assign n2312 = n3236 & n2311;
  assign n2313 = n3236 | n2311;
  assign n2314 = ~n2312 & n2313;
  assign n2315 = x23 & x46;
  assign n2316 = n2314 & n2315;
  assign n2317 = n2314 | n2315;
  assign n2318 = ~n2316 & n2317;
  assign n2319 = n3234 & n2318;
  assign n2320 = n3234 | n2318;
  assign n2321 = ~n2319 & n2320;
  assign n2322 = x22 & x47;
  assign n2323 = n2321 & n2322;
  assign n2324 = n2321 | n2322;
  assign n2325 = ~n2323 & n2324;
  assign n2326 = n2248 & n2325;
  assign n2327 = n2248 | n2325;
  assign n2328 = ~n2326 & n2327;
  assign n3266 = n2323 | n2325;
  assign n3267 = (n2248 & n2323) | (n2248 & n3266) | (n2323 & n3266);
  assign n3268 = n2316 | n2318;
  assign n3269 = (n2316 & n3234) | (n2316 & n3268) | (n3234 & n3268);
  assign n3270 = n2309 | n2311;
  assign n3271 = (n2309 & n3236) | (n2309 & n3270) | (n3236 & n3270);
  assign n3272 = n2302 | n2304;
  assign n3273 = (n2302 & n3238) | (n2302 & n3272) | (n3238 & n3272);
  assign n3274 = n2295 | n2297;
  assign n3275 = (n2295 & n3240) | (n2295 & n3274) | (n3240 & n3274);
  assign n3276 = n2288 | n2290;
  assign n3277 = (n2288 & n3242) | (n2288 & n3276) | (n3242 & n3276);
  assign n2339 = x31 & x39;
  assign n3281 = n2262 | n3250;
  assign n3751 = (n2179 & n3250) | (n2179 & n3281) | (n3250 & n3281);
  assign n3283 = n2339 & n3751;
  assign n4108 = n2339 & n3942;
  assign n4135 = n3699 & n4108;
  assign n4109 = (n3705 & n4135) | (n3705 & n4108) | (n4135 & n4108);
  assign n4056 = n2259 & n2339;
  assign n4110 = n3936 & n4056;
  assign n4106 = (n3663 & n4109) | (n3663 & n4110) | (n4109 & n4110);
  assign n4057 = (n2174 & n4106) | (n2174 & n4056) | (n4106 & n4056);
  assign n4060 = (n3663 & n4109) | (n3663 & n4110) | (n4109 & n4110);
  assign n3951 = (n3717 & n4057) | (n3717 & n4060) | (n4057 & n4060);
  assign n3753 = (n2262 & n2339) | (n2262 & n3951) | (n2339 & n3951);
  assign n3754 = (n3216 & n3283) | (n3216 & n3753) | (n3283 & n3753);
  assign n3755 = (n3215 & n3283) | (n3215 & n3753) | (n3283 & n3753);
  assign n3756 = (n3694 & n3754) | (n3694 & n3755) | (n3754 & n3755);
  assign n3286 = n2339 | n3751;
  assign n4114 = n2339 | n3942;
  assign n4136 = (n2339 & n3699) | (n2339 & n4114) | (n3699 & n4114);
  assign n4115 = (n3705 & n4136) | (n3705 & n4114) | (n4136 & n4114);
  assign n4062 = n2259 | n2339;
  assign n4116 = (n2339 & n3936) | (n2339 & n4062) | (n3936 & n4062);
  assign n4112 = (n3663 & n4115) | (n3663 & n4116) | (n4115 & n4116);
  assign n4063 = (n2174 & n4112) | (n2174 & n4062) | (n4112 & n4062);
  assign n4066 = (n3663 & n4115) | (n3663 & n4116) | (n4115 & n4116);
  assign n3954 = (n3717 & n4063) | (n3717 & n4066) | (n4063 & n4066);
  assign n3758 = n2262 | n3954;
  assign n3759 = (n3216 & n3286) | (n3216 & n3758) | (n3286 & n3758);
  assign n3760 = (n3215 & n3286) | (n3215 & n3758) | (n3286 & n3758);
  assign n3761 = (n3694 & n3759) | (n3694 & n3760) | (n3759 & n3760);
  assign n2342 = ~n3756 & n3761;
  assign n3290 = n2267 & n2342;
  assign n3762 = (n2269 & n2342) | (n2269 & n3290) | (n2342 & n3290);
  assign n3291 = (n3734 & n3762) | (n3734 & n3290) | (n3762 & n3290);
  assign n3293 = n2267 | n2342;
  assign n3763 = n2269 | n3293;
  assign n3294 = (n3734 & n3763) | (n3734 & n3293) | (n3763 & n3293);
  assign n2345 = ~n3291 & n3294;
  assign n2346 = x30 & x40;
  assign n2347 = n2345 & n2346;
  assign n2348 = n2345 | n2346;
  assign n2349 = ~n2347 & n2348;
  assign n3295 = n2274 & n2349;
  assign n3764 = (n2349 & n3258) | (n2349 & n3295) | (n3258 & n3295);
  assign n3765 = (n2276 & n2349) | (n2276 & n3295) | (n2349 & n3295);
  assign n3766 = (n3226 & n3764) | (n3226 & n3765) | (n3764 & n3765);
  assign n3297 = n2274 | n2349;
  assign n3767 = n3258 | n3297;
  assign n3768 = n2276 | n3297;
  assign n3769 = (n3226 & n3767) | (n3226 & n3768) | (n3767 & n3768);
  assign n2352 = ~n3766 & n3769;
  assign n2353 = x29 & x41;
  assign n2354 = n2352 & n2353;
  assign n2355 = n2352 | n2353;
  assign n2356 = ~n2354 & n2355;
  assign n3299 = n2281 & n2356;
  assign n3300 = (n2356 & n3263) | (n2356 & n3299) | (n3263 & n3299);
  assign n3301 = n2281 | n2356;
  assign n3302 = n3263 | n3301;
  assign n2359 = ~n3300 & n3302;
  assign n2360 = x28 & x42;
  assign n2361 = n2359 & n2360;
  assign n2362 = n2359 | n2360;
  assign n2363 = ~n2361 & n2362;
  assign n2364 = n3277 & n2363;
  assign n2365 = n3277 | n2363;
  assign n2366 = ~n2364 & n2365;
  assign n2367 = x27 & x43;
  assign n2368 = n2366 & n2367;
  assign n2369 = n2366 | n2367;
  assign n2370 = ~n2368 & n2369;
  assign n2371 = n3275 & n2370;
  assign n2372 = n3275 | n2370;
  assign n2373 = ~n2371 & n2372;
  assign n2374 = x26 & x44;
  assign n2375 = n2373 & n2374;
  assign n2376 = n2373 | n2374;
  assign n2377 = ~n2375 & n2376;
  assign n2378 = n3273 & n2377;
  assign n2379 = n3273 | n2377;
  assign n2380 = ~n2378 & n2379;
  assign n2381 = x25 & x45;
  assign n2382 = n2380 & n2381;
  assign n2383 = n2380 | n2381;
  assign n2384 = ~n2382 & n2383;
  assign n2385 = n3271 & n2384;
  assign n2386 = n3271 | n2384;
  assign n2387 = ~n2385 & n2386;
  assign n2388 = x24 & x46;
  assign n2389 = n2387 & n2388;
  assign n2390 = n2387 | n2388;
  assign n2391 = ~n2389 & n2390;
  assign n2392 = n3269 & n2391;
  assign n2393 = n3269 | n2391;
  assign n2394 = ~n2392 & n2393;
  assign n2395 = x23 & x47;
  assign n2396 = n2394 & n2395;
  assign n2397 = n2394 | n2395;
  assign n2398 = ~n2396 & n2397;
  assign n2399 = n3267 & n2398;
  assign n2400 = n3267 | n2398;
  assign n2401 = ~n2399 & n2400;
  assign n3303 = n2396 | n2398;
  assign n3304 = (n2396 & n3267) | (n2396 & n3303) | (n3267 & n3303);
  assign n3305 = n2389 | n2391;
  assign n3306 = (n2389 & n3269) | (n2389 & n3305) | (n3269 & n3305);
  assign n3307 = n2382 | n2384;
  assign n3308 = (n2382 & n3271) | (n2382 & n3307) | (n3271 & n3307);
  assign n3309 = n2375 | n2377;
  assign n3310 = (n2375 & n3273) | (n2375 & n3309) | (n3273 & n3309);
  assign n3311 = n2368 | n2370;
  assign n3312 = (n2368 & n3275) | (n2368 & n3311) | (n3275 & n3311);
  assign n3313 = n2361 | n2363;
  assign n3314 = (n2361 & n3277) | (n2361 & n3313) | (n3277 & n3313);
  assign n3316 = n2347 | n2349;
  assign n3770 = n2274 | n2347;
  assign n3771 = (n2347 & n2349) | (n2347 & n3770) | (n2349 & n3770);
  assign n3772 = (n3258 & n3316) | (n3258 & n3771) | (n3316 & n3771);
  assign n3773 = (n2276 & n3316) | (n2276 & n3771) | (n3316 & n3771);
  assign n3774 = (n3226 & n3772) | (n3226 & n3773) | (n3772 & n3773);
  assign n2411 = x31 & x40;
  assign n3318 = n2411 & n3756;
  assign n3775 = (n2411 & n3318) | (n2411 & n3762) | (n3318 & n3762);
  assign n3955 = (n2342 & n2411) | (n2342 & n3318) | (n2411 & n3318);
  assign n4067 = n2411 & n3756;
  assign n3957 = (n2267 & n3955) | (n2267 & n4067) | (n3955 & n4067);
  assign n3777 = (n3734 & n3775) | (n3734 & n3957) | (n3775 & n3957);
  assign n3320 = n2411 | n3756;
  assign n3778 = n3320 | n3762;
  assign n3958 = n2342 | n3320;
  assign n3959 = (n2267 & n3320) | (n2267 & n3958) | (n3320 & n3958);
  assign n3780 = (n3734 & n3778) | (n3734 & n3959) | (n3778 & n3959);
  assign n2414 = ~n3777 & n3780;
  assign n2415 = n3774 & n2414;
  assign n2416 = n3774 | n2414;
  assign n2417 = ~n2415 & n2416;
  assign n2418 = x30 & x41;
  assign n2419 = n2417 & n2418;
  assign n2420 = n2417 | n2418;
  assign n2421 = ~n2419 & n2420;
  assign n3322 = n2354 & n2421;
  assign n3323 = (n2421 & n3300) | (n2421 & n3322) | (n3300 & n3322);
  assign n3324 = n2354 | n2421;
  assign n3325 = n3300 | n3324;
  assign n2424 = ~n3323 & n3325;
  assign n2425 = x29 & x42;
  assign n2426 = n2424 & n2425;
  assign n2427 = n2424 | n2425;
  assign n2428 = ~n2426 & n2427;
  assign n2429 = n3314 & n2428;
  assign n2430 = n3314 | n2428;
  assign n2431 = ~n2429 & n2430;
  assign n2432 = x28 & x43;
  assign n2433 = n2431 & n2432;
  assign n2434 = n2431 | n2432;
  assign n2435 = ~n2433 & n2434;
  assign n2436 = n3312 & n2435;
  assign n2437 = n3312 | n2435;
  assign n2438 = ~n2436 & n2437;
  assign n2439 = x27 & x44;
  assign n2440 = n2438 & n2439;
  assign n2441 = n2438 | n2439;
  assign n2442 = ~n2440 & n2441;
  assign n2443 = n3310 & n2442;
  assign n2444 = n3310 | n2442;
  assign n2445 = ~n2443 & n2444;
  assign n2446 = x26 & x45;
  assign n2447 = n2445 & n2446;
  assign n2448 = n2445 | n2446;
  assign n2449 = ~n2447 & n2448;
  assign n2450 = n3308 & n2449;
  assign n2451 = n3308 | n2449;
  assign n2452 = ~n2450 & n2451;
  assign n2453 = x25 & x46;
  assign n2454 = n2452 & n2453;
  assign n2455 = n2452 | n2453;
  assign n2456 = ~n2454 & n2455;
  assign n2457 = n3306 & n2456;
  assign n2458 = n3306 | n2456;
  assign n2459 = ~n2457 & n2458;
  assign n2460 = x24 & x47;
  assign n2461 = n2459 & n2460;
  assign n2462 = n2459 | n2460;
  assign n2463 = ~n2461 & n2462;
  assign n2464 = n3304 & n2463;
  assign n2465 = n3304 | n2463;
  assign n2466 = ~n2464 & n2465;
  assign n3326 = n2461 | n2463;
  assign n3327 = (n2461 & n3304) | (n2461 & n3326) | (n3304 & n3326);
  assign n3328 = n2454 | n2456;
  assign n3329 = (n2454 & n3306) | (n2454 & n3328) | (n3306 & n3328);
  assign n3330 = n2447 | n2449;
  assign n3331 = (n2447 & n3308) | (n2447 & n3330) | (n3308 & n3330);
  assign n3332 = n2440 | n2442;
  assign n3333 = (n2440 & n3310) | (n2440 & n3332) | (n3310 & n3332);
  assign n3334 = n2433 | n2435;
  assign n3335 = (n2433 & n3312) | (n2433 & n3334) | (n3312 & n3334);
  assign n3336 = n2426 | n2428;
  assign n3337 = (n2426 & n3314) | (n2426 & n3336) | (n3314 & n3336);
  assign n2475 = x31 & x41;
  assign n3963 = n2411 & n2475;
  assign n4068 = n3756 & n3963;
  assign n3964 = (n3762 & n4068) | (n3762 & n3963) | (n4068 & n3963);
  assign n3960 = n2475 & n3957;
  assign n3961 = (n3734 & n3964) | (n3734 & n3960) | (n3964 & n3960);
  assign n3782 = (n2414 & n2475) | (n2414 & n3961) | (n2475 & n3961);
  assign n3784 = n2475 & n3957;
  assign n3785 = (n3734 & n3964) | (n3734 & n3784) | (n3964 & n3784);
  assign n3342 = (n3774 & n3782) | (n3774 & n3785) | (n3782 & n3785);
  assign n3968 = n2411 | n2475;
  assign n4069 = (n2475 & n3756) | (n2475 & n3968) | (n3756 & n3968);
  assign n3969 = (n3762 & n4069) | (n3762 & n3968) | (n4069 & n3968);
  assign n3965 = n2475 | n3957;
  assign n3966 = (n3734 & n3969) | (n3734 & n3965) | (n3969 & n3965);
  assign n3787 = n2414 | n3966;
  assign n3789 = n2475 | n3957;
  assign n3790 = (n3734 & n3969) | (n3734 & n3789) | (n3969 & n3789);
  assign n3345 = (n3774 & n3787) | (n3774 & n3790) | (n3787 & n3790);
  assign n2478 = ~n3342 & n3345;
  assign n3346 = n2419 & n2478;
  assign n3791 = (n2478 & n3322) | (n2478 & n3346) | (n3322 & n3346);
  assign n3792 = (n2421 & n2478) | (n2421 & n3346) | (n2478 & n3346);
  assign n3793 = (n3300 & n3791) | (n3300 & n3792) | (n3791 & n3792);
  assign n3348 = n2419 | n2478;
  assign n3794 = n3322 | n3348;
  assign n3795 = n2421 | n3348;
  assign n3796 = (n3300 & n3794) | (n3300 & n3795) | (n3794 & n3795);
  assign n2481 = ~n3793 & n3796;
  assign n2482 = x30 & x42;
  assign n2483 = n2481 & n2482;
  assign n2484 = n2481 | n2482;
  assign n2485 = ~n2483 & n2484;
  assign n2486 = n3337 & n2485;
  assign n2487 = n3337 | n2485;
  assign n2488 = ~n2486 & n2487;
  assign n2489 = x29 & x43;
  assign n2490 = n2488 & n2489;
  assign n2491 = n2488 | n2489;
  assign n2492 = ~n2490 & n2491;
  assign n2493 = n3335 & n2492;
  assign n2494 = n3335 | n2492;
  assign n2495 = ~n2493 & n2494;
  assign n2496 = x28 & x44;
  assign n2497 = n2495 & n2496;
  assign n2498 = n2495 | n2496;
  assign n2499 = ~n2497 & n2498;
  assign n2500 = n3333 & n2499;
  assign n2501 = n3333 | n2499;
  assign n2502 = ~n2500 & n2501;
  assign n2503 = x27 & x45;
  assign n2504 = n2502 & n2503;
  assign n2505 = n2502 | n2503;
  assign n2506 = ~n2504 & n2505;
  assign n2507 = n3331 & n2506;
  assign n2508 = n3331 | n2506;
  assign n2509 = ~n2507 & n2508;
  assign n2510 = x26 & x46;
  assign n2511 = n2509 & n2510;
  assign n2512 = n2509 | n2510;
  assign n2513 = ~n2511 & n2512;
  assign n2514 = n3329 & n2513;
  assign n2515 = n3329 | n2513;
  assign n2516 = ~n2514 & n2515;
  assign n2517 = x25 & x47;
  assign n2518 = n2516 & n2517;
  assign n2519 = n2516 | n2517;
  assign n2520 = ~n2518 & n2519;
  assign n2521 = n3327 & n2520;
  assign n2522 = n3327 | n2520;
  assign n2523 = ~n2521 & n2522;
  assign n3350 = n2518 | n2520;
  assign n3351 = (n2518 & n3327) | (n2518 & n3350) | (n3327 & n3350);
  assign n3352 = n2511 | n2513;
  assign n3353 = (n2511 & n3329) | (n2511 & n3352) | (n3329 & n3352);
  assign n3354 = n2504 | n2506;
  assign n3355 = (n2504 & n3331) | (n2504 & n3354) | (n3331 & n3354);
  assign n3356 = n2497 | n2499;
  assign n3357 = (n2497 & n3333) | (n2497 & n3356) | (n3333 & n3356);
  assign n3358 = n2490 | n2492;
  assign n3359 = (n2490 & n3335) | (n2490 & n3358) | (n3335 & n3358);
  assign n2531 = x31 & x42;
  assign n3363 = n2478 | n3342;
  assign n3797 = (n2419 & n3342) | (n2419 & n3363) | (n3342 & n3363);
  assign n3365 = n2531 & n3797;
  assign n4120 = n2531 & n3963;
  assign n4137 = n3756 & n4120;
  assign n4121 = (n3762 & n4137) | (n3762 & n4120) | (n4137 & n4120);
  assign n4071 = n2475 & n2531;
  assign n4122 = n3957 & n4071;
  assign n4118 = (n3734 & n4121) | (n3734 & n4122) | (n4121 & n4122);
  assign n4072 = (n2414 & n4118) | (n2414 & n4071) | (n4118 & n4071);
  assign n4075 = (n3734 & n4121) | (n3734 & n4122) | (n4121 & n4122);
  assign n3972 = (n3774 & n4072) | (n3774 & n4075) | (n4072 & n4075);
  assign n3799 = (n2478 & n2531) | (n2478 & n3972) | (n2531 & n3972);
  assign n3800 = (n3322 & n3365) | (n3322 & n3799) | (n3365 & n3799);
  assign n3801 = (n2421 & n3365) | (n2421 & n3799) | (n3365 & n3799);
  assign n3802 = (n3300 & n3800) | (n3300 & n3801) | (n3800 & n3801);
  assign n3368 = n2531 | n3797;
  assign n4126 = n2531 | n3963;
  assign n4138 = (n2531 & n3756) | (n2531 & n4126) | (n3756 & n4126);
  assign n4127 = (n3762 & n4138) | (n3762 & n4126) | (n4138 & n4126);
  assign n4077 = n2475 | n2531;
  assign n4128 = (n2531 & n3957) | (n2531 & n4077) | (n3957 & n4077);
  assign n4124 = (n3734 & n4127) | (n3734 & n4128) | (n4127 & n4128);
  assign n4078 = (n2414 & n4124) | (n2414 & n4077) | (n4124 & n4077);
  assign n4081 = (n3734 & n4127) | (n3734 & n4128) | (n4127 & n4128);
  assign n3975 = (n3774 & n4078) | (n3774 & n4081) | (n4078 & n4081);
  assign n3804 = n2478 | n3975;
  assign n3805 = (n3322 & n3368) | (n3322 & n3804) | (n3368 & n3804);
  assign n3806 = (n2421 & n3368) | (n2421 & n3804) | (n3368 & n3804);
  assign n3807 = (n3300 & n3805) | (n3300 & n3806) | (n3805 & n3806);
  assign n2534 = ~n3802 & n3807;
  assign n3809 = n2483 & n2534;
  assign n3976 = (n2485 & n2534) | (n2485 & n3809) | (n2534 & n3809);
  assign n3810 = (n3337 & n3976) | (n3337 & n3809) | (n3976 & n3809);
  assign n3812 = n2483 | n2534;
  assign n3977 = n2485 | n3812;
  assign n3813 = (n3337 & n3977) | (n3337 & n3812) | (n3977 & n3812);
  assign n2537 = ~n3810 & n3813;
  assign n2538 = x30 & x43;
  assign n2539 = n2537 & n2538;
  assign n2540 = n2537 | n2538;
  assign n2541 = ~n2539 & n2540;
  assign n2542 = n3359 & n2541;
  assign n2543 = n3359 | n2541;
  assign n2544 = ~n2542 & n2543;
  assign n2545 = x29 & x44;
  assign n2546 = n2544 & n2545;
  assign n2547 = n2544 | n2545;
  assign n2548 = ~n2546 & n2547;
  assign n2549 = n3357 & n2548;
  assign n2550 = n3357 | n2548;
  assign n2551 = ~n2549 & n2550;
  assign n2552 = x28 & x45;
  assign n2553 = n2551 & n2552;
  assign n2554 = n2551 | n2552;
  assign n2555 = ~n2553 & n2554;
  assign n2556 = n3355 & n2555;
  assign n2557 = n3355 | n2555;
  assign n2558 = ~n2556 & n2557;
  assign n2559 = x27 & x46;
  assign n2560 = n2558 & n2559;
  assign n2561 = n2558 | n2559;
  assign n2562 = ~n2560 & n2561;
  assign n2563 = n3353 & n2562;
  assign n2564 = n3353 | n2562;
  assign n2565 = ~n2563 & n2564;
  assign n2566 = x26 & x47;
  assign n2567 = n2565 & n2566;
  assign n2568 = n2565 | n2566;
  assign n2569 = ~n2567 & n2568;
  assign n2570 = n3351 & n2569;
  assign n2571 = n3351 | n2569;
  assign n2572 = ~n2570 & n2571;
  assign n3371 = n2567 | n2569;
  assign n3372 = (n2567 & n3351) | (n2567 & n3371) | (n3351 & n3371);
  assign n3373 = n2560 | n2562;
  assign n3374 = (n2560 & n3353) | (n2560 & n3373) | (n3353 & n3373);
  assign n3375 = n2553 | n2555;
  assign n3376 = (n2553 & n3355) | (n2553 & n3375) | (n3355 & n3375);
  assign n3377 = n2546 | n2548;
  assign n3378 = (n2546 & n3357) | (n2546 & n3377) | (n3357 & n3377);
  assign n2579 = x31 & x43;
  assign n3384 = n2579 & n3802;
  assign n3814 = n2579 & n3802;
  assign n3815 = (n2534 & n2579) | (n2534 & n3814) | (n2579 & n3814);
  assign n3817 = (n2483 & n3384) | (n2483 & n3815) | (n3384 & n3815);
  assign n3978 = n3384 | n3815;
  assign n3979 = (n2485 & n3817) | (n2485 & n3978) | (n3817 & n3978);
  assign n3818 = (n3337 & n3979) | (n3337 & n3817) | (n3979 & n3817);
  assign n3387 = n2579 | n3802;
  assign n3819 = n2579 | n3802;
  assign n3820 = n2534 | n3819;
  assign n3822 = (n2483 & n3387) | (n2483 & n3820) | (n3387 & n3820);
  assign n3980 = n3387 | n3820;
  assign n3981 = (n2485 & n3822) | (n2485 & n3980) | (n3822 & n3980);
  assign n3823 = (n3337 & n3981) | (n3337 & n3822) | (n3981 & n3822);
  assign n2582 = ~n3818 & n3823;
  assign n3825 = n2539 & n2582;
  assign n3982 = (n2541 & n2582) | (n2541 & n3825) | (n2582 & n3825);
  assign n3826 = (n3359 & n3982) | (n3359 & n3825) | (n3982 & n3825);
  assign n3828 = n2539 | n2582;
  assign n3983 = n2541 | n3828;
  assign n3829 = (n3359 & n3983) | (n3359 & n3828) | (n3983 & n3828);
  assign n2585 = ~n3826 & n3829;
  assign n2586 = x30 & x44;
  assign n2587 = n2585 & n2586;
  assign n2588 = n2585 | n2586;
  assign n2589 = ~n2587 & n2588;
  assign n2590 = n3378 & n2589;
  assign n2591 = n3378 | n2589;
  assign n2592 = ~n2590 & n2591;
  assign n2593 = x29 & x45;
  assign n2594 = n2592 & n2593;
  assign n2595 = n2592 | n2593;
  assign n2596 = ~n2594 & n2595;
  assign n2597 = n3376 & n2596;
  assign n2598 = n3376 | n2596;
  assign n2599 = ~n2597 & n2598;
  assign n2600 = x28 & x46;
  assign n2601 = n2599 & n2600;
  assign n2602 = n2599 | n2600;
  assign n2603 = ~n2601 & n2602;
  assign n2604 = n3374 & n2603;
  assign n2605 = n3374 | n2603;
  assign n2606 = ~n2604 & n2605;
  assign n2607 = x27 & x47;
  assign n2608 = n2606 & n2607;
  assign n2609 = n2606 | n2607;
  assign n2610 = ~n2608 & n2609;
  assign n2611 = n3372 & n2610;
  assign n2612 = n3372 | n2610;
  assign n2613 = ~n2611 & n2612;
  assign n3389 = n2608 | n2610;
  assign n3390 = (n2608 & n3372) | (n2608 & n3389) | (n3372 & n3389);
  assign n3391 = n2601 | n2603;
  assign n3392 = (n2601 & n3374) | (n2601 & n3391) | (n3374 & n3391);
  assign n3393 = n2594 | n2596;
  assign n3394 = (n2594 & n3376) | (n2594 & n3393) | (n3376 & n3393);
  assign n2619 = x31 & x44;
  assign n3984 = n2619 & n3979;
  assign n3985 = n2619 & n3817;
  assign n3986 = (n3337 & n3984) | (n3337 & n3985) | (n3984 & n3985);
  assign n3831 = (n2582 & n2619) | (n2582 & n3986) | (n2619 & n3986);
  assign n3987 = (n2539 & n3831) | (n2539 & n3986) | (n3831 & n3986);
  assign n4082 = n2619 | n3986;
  assign n4083 = (n2582 & n3986) | (n2582 & n4082) | (n3986 & n4082);
  assign n3989 = (n2541 & n3987) | (n2541 & n4083) | (n3987 & n4083);
  assign n3833 = (n2539 & n3986) | (n2539 & n3831) | (n3986 & n3831);
  assign n3834 = (n3359 & n3989) | (n3359 & n3833) | (n3989 & n3833);
  assign n3990 = n2619 | n3979;
  assign n3991 = n2619 | n3817;
  assign n3992 = (n3337 & n3990) | (n3337 & n3991) | (n3990 & n3991);
  assign n3836 = n2582 | n3992;
  assign n3993 = (n2539 & n3836) | (n2539 & n3992) | (n3836 & n3992);
  assign n4084 = n2582 | n3992;
  assign n3995 = (n2541 & n3993) | (n2541 & n4084) | (n3993 & n4084);
  assign n3838 = (n2539 & n3992) | (n2539 & n3836) | (n3992 & n3836);
  assign n3839 = (n3359 & n3995) | (n3359 & n3838) | (n3995 & n3838);
  assign n2622 = ~n3834 & n3839;
  assign n3841 = n2587 & n2622;
  assign n3996 = (n2589 & n2622) | (n2589 & n3841) | (n2622 & n3841);
  assign n3842 = (n3378 & n3996) | (n3378 & n3841) | (n3996 & n3841);
  assign n3844 = n2587 | n2622;
  assign n3997 = n2589 | n3844;
  assign n3845 = (n3378 & n3997) | (n3378 & n3844) | (n3997 & n3844);
  assign n2625 = ~n3842 & n3845;
  assign n2626 = x30 & x45;
  assign n2627 = n2625 & n2626;
  assign n2628 = n2625 | n2626;
  assign n2629 = ~n2627 & n2628;
  assign n2630 = n3394 & n2629;
  assign n2631 = n3394 | n2629;
  assign n2632 = ~n2630 & n2631;
  assign n2633 = x29 & x46;
  assign n2634 = n2632 & n2633;
  assign n2635 = n2632 | n2633;
  assign n2636 = ~n2634 & n2635;
  assign n2637 = n3392 & n2636;
  assign n2638 = n3392 | n2636;
  assign n2639 = ~n2637 & n2638;
  assign n2640 = x28 & x47;
  assign n2641 = n2639 & n2640;
  assign n2642 = n2639 | n2640;
  assign n2643 = ~n2641 & n2642;
  assign n2644 = n3390 & n2643;
  assign n2645 = n3390 | n2643;
  assign n2646 = ~n2644 & n2645;
  assign n3405 = n2641 | n2643;
  assign n3406 = (n2641 & n3390) | (n2641 & n3405) | (n3390 & n3405);
  assign n3407 = n2634 | n2636;
  assign n3408 = (n2634 & n3392) | (n2634 & n3407) | (n3392 & n3407);
  assign n2651 = x31 & x45;
  assign n3998 = n2651 & n3989;
  assign n3999 = n2651 & n3833;
  assign n4000 = (n3359 & n3998) | (n3359 & n3999) | (n3998 & n3999);
  assign n3847 = (n2622 & n2651) | (n2622 & n4000) | (n2651 & n4000);
  assign n4001 = (n2587 & n3847) | (n2587 & n4000) | (n3847 & n4000);
  assign n4085 = n2651 | n4000;
  assign n4086 = (n2622 & n4000) | (n2622 & n4085) | (n4000 & n4085);
  assign n4003 = (n2589 & n4001) | (n2589 & n4086) | (n4001 & n4086);
  assign n3849 = (n2587 & n4000) | (n2587 & n3847) | (n4000 & n3847);
  assign n3850 = (n3378 & n4003) | (n3378 & n3849) | (n4003 & n3849);
  assign n4004 = n2651 | n3989;
  assign n4005 = n2651 | n3833;
  assign n4006 = (n3359 & n4004) | (n3359 & n4005) | (n4004 & n4005);
  assign n3852 = n2622 | n4006;
  assign n4007 = (n2587 & n3852) | (n2587 & n4006) | (n3852 & n4006);
  assign n4087 = n2622 | n4006;
  assign n4009 = (n2589 & n4007) | (n2589 & n4087) | (n4007 & n4087);
  assign n3854 = (n2587 & n4006) | (n2587 & n3852) | (n4006 & n3852);
  assign n3855 = (n3378 & n4009) | (n3378 & n3854) | (n4009 & n3854);
  assign n2654 = ~n3850 & n3855;
  assign n3857 = n2627 & n2654;
  assign n4010 = (n2629 & n2654) | (n2629 & n3857) | (n2654 & n3857);
  assign n3858 = (n3394 & n4010) | (n3394 & n3857) | (n4010 & n3857);
  assign n3860 = n2627 | n2654;
  assign n4011 = n2629 | n3860;
  assign n3861 = (n3394 & n4011) | (n3394 & n3860) | (n4011 & n3860);
  assign n2657 = ~n3858 & n3861;
  assign n2658 = x30 & x46;
  assign n2659 = n2657 & n2658;
  assign n2660 = n2657 | n2658;
  assign n2661 = ~n2659 & n2660;
  assign n2662 = n3408 & n2661;
  assign n2663 = n3408 | n2661;
  assign n2664 = ~n2662 & n2663;
  assign n2665 = x29 & x47;
  assign n2666 = n2664 & n2665;
  assign n2667 = n2664 | n2665;
  assign n2668 = ~n2666 & n2667;
  assign n2669 = n3406 & n2668;
  assign n2670 = n3406 | n2668;
  assign n2671 = ~n2669 & n2670;
  assign n3419 = n2666 | n2668;
  assign n3420 = (n2666 & n3406) | (n2666 & n3419) | (n3406 & n3419);
  assign n2675 = x31 & x46;
  assign n4012 = n2675 & n4003;
  assign n4013 = n2675 & n3849;
  assign n4014 = (n3378 & n4012) | (n3378 & n4013) | (n4012 & n4013);
  assign n3863 = (n2654 & n2675) | (n2654 & n4014) | (n2675 & n4014);
  assign n4015 = (n2627 & n3863) | (n2627 & n4014) | (n3863 & n4014);
  assign n4088 = n2675 | n4014;
  assign n4089 = (n2654 & n4014) | (n2654 & n4088) | (n4014 & n4088);
  assign n4017 = (n2629 & n4015) | (n2629 & n4089) | (n4015 & n4089);
  assign n3865 = (n2627 & n4014) | (n2627 & n3863) | (n4014 & n3863);
  assign n3866 = (n3394 & n4017) | (n3394 & n3865) | (n4017 & n3865);
  assign n4018 = n2675 | n4003;
  assign n4019 = n2675 | n3849;
  assign n4020 = (n3378 & n4018) | (n3378 & n4019) | (n4018 & n4019);
  assign n3868 = n2654 | n4020;
  assign n4021 = (n2627 & n3868) | (n2627 & n4020) | (n3868 & n4020);
  assign n4090 = n2654 | n4020;
  assign n4023 = (n2629 & n4021) | (n2629 & n4090) | (n4021 & n4090);
  assign n3870 = (n2627 & n4020) | (n2627 & n3868) | (n4020 & n3868);
  assign n3871 = (n3394 & n4023) | (n3394 & n3870) | (n4023 & n3870);
  assign n2678 = ~n3866 & n3871;
  assign n3873 = n2659 & n2678;
  assign n4024 = (n2661 & n2678) | (n2661 & n3873) | (n2678 & n3873);
  assign n3874 = (n3408 & n4024) | (n3408 & n3873) | (n4024 & n3873);
  assign n3876 = n2659 | n2678;
  assign n4025 = n2661 | n3876;
  assign n3877 = (n3408 & n4025) | (n3408 & n3876) | (n4025 & n3876);
  assign n2681 = ~n3874 & n3877;
  assign n2682 = x30 & x47;
  assign n2683 = n2681 & n2682;
  assign n2684 = n2681 | n2682;
  assign n2685 = ~n2683 & n2684;
  assign n2686 = n3420 & n2685;
  assign n2687 = n3420 | n2685;
  assign n2688 = ~n2686 & n2687;
  assign n2691 = x31 & x47;
  assign n4026 = n2691 & n4017;
  assign n4027 = n2691 & n3865;
  assign n4028 = (n3394 & n4026) | (n3394 & n4027) | (n4026 & n4027);
  assign n3879 = (n2678 & n2691) | (n2678 & n4028) | (n2691 & n4028);
  assign n4029 = (n2659 & n3879) | (n2659 & n4028) | (n3879 & n4028);
  assign n4091 = n2691 | n4028;
  assign n4092 = (n2678 & n4028) | (n2678 & n4091) | (n4028 & n4091);
  assign n4031 = (n2661 & n4029) | (n2661 & n4092) | (n4029 & n4092);
  assign n3881 = (n2659 & n4028) | (n2659 & n3879) | (n4028 & n3879);
  assign n3882 = (n3408 & n4031) | (n3408 & n3881) | (n4031 & n3881);
  assign n4032 = n2691 | n4017;
  assign n4033 = n2691 | n3865;
  assign n4034 = (n3394 & n4032) | (n3394 & n4033) | (n4032 & n4033);
  assign n3884 = n2678 | n4034;
  assign n4035 = (n2659 & n3884) | (n2659 & n4034) | (n3884 & n4034);
  assign n4093 = n2678 | n4034;
  assign n4037 = (n2661 & n4035) | (n2661 & n4093) | (n4035 & n4093);
  assign n3886 = (n2659 & n4034) | (n2659 & n3884) | (n4034 & n3884);
  assign n3887 = (n3408 & n4037) | (n3408 & n3886) | (n4037 & n3886);
  assign n2694 = ~n3882 & n3887;
  assign n3889 = n2683 & n2694;
  assign n4038 = (n2685 & n2694) | (n2685 & n3889) | (n2694 & n3889);
  assign n3890 = (n3420 & n4038) | (n3420 & n3889) | (n4038 & n3889);
  assign n3892 = n2683 | n2694;
  assign n4039 = n2685 | n3892;
  assign n3893 = (n3420 & n4039) | (n3420 & n3892) | (n4039 & n3892);
  assign n2697 = ~n3890 & n3893;
  assign n3441 = n2694 | n3882;
  assign n3895 = (n2683 & n3441) | (n2683 & n3882) | (n3441 & n3882);
  assign n4094 = n2694 | n3882;
  assign n4041 = (n2685 & n3895) | (n2685 & n4094) | (n3895 & n4094);
  assign n3896 = (n3420 & n4041) | (n3420 & n3895) | (n4041 & n3895);
  assign n4203 = x48 & x80;
  assign n4204 = x49 & x80;
  assign n4205 = x48 & x81;
  assign n4206 = n4204 & n4205;
  assign n4207 = n4204 | n4205;
  assign n4208 = ~n4206 & n4207;
  assign n4209 = x50 & x80;
  assign n4210 = x49 & x81;
  assign n4211 = n4209 & n4210;
  assign n4212 = n4209 | n4210;
  assign n4213 = ~n4211 & n4212;
  assign n4214 = n4206 & n4213;
  assign n4215 = n4206 | n4213;
  assign n4216 = ~n4214 & n4215;
  assign n4217 = x48 & x82;
  assign n4218 = n4216 & n4217;
  assign n4219 = n4216 | n4217;
  assign n4220 = ~n4218 & n4219;
  assign n12043 = n4206 | n4211;
  assign n12044 = (n4211 & n4213) | (n4211 & n12043) | (n4213 & n12043);
  assign n4222 = x51 & x80;
  assign n4223 = x50 & x81;
  assign n4224 = n4222 & n4223;
  assign n4225 = n4222 | n4223;
  assign n4226 = ~n4224 & n4225;
  assign n4227 = n12044 & n4226;
  assign n4228 = n12044 | n4226;
  assign n4229 = ~n4227 & n4228;
  assign n4230 = x49 & x82;
  assign n4231 = n4229 & n4230;
  assign n4232 = n4229 | n4230;
  assign n4233 = ~n4231 & n4232;
  assign n4234 = n4218 & n4233;
  assign n4235 = n4218 | n4233;
  assign n4236 = ~n4234 & n4235;
  assign n4237 = x48 & x83;
  assign n4238 = n4236 & n4237;
  assign n4239 = n4236 | n4237;
  assign n4240 = ~n4238 & n4239;
  assign n12045 = n4218 | n4231;
  assign n12046 = (n4231 & n4233) | (n4231 & n12045) | (n4233 & n12045);
  assign n12047 = n4224 | n4226;
  assign n12048 = (n4224 & n12044) | (n4224 & n12047) | (n12044 & n12047);
  assign n4243 = x52 & x80;
  assign n4244 = x51 & x81;
  assign n4245 = n4243 & n4244;
  assign n4246 = n4243 | n4244;
  assign n4247 = ~n4245 & n4246;
  assign n4248 = n12048 & n4247;
  assign n4249 = n12048 | n4247;
  assign n4250 = ~n4248 & n4249;
  assign n4251 = x50 & x82;
  assign n4252 = n4250 & n4251;
  assign n4253 = n4250 | n4251;
  assign n4254 = ~n4252 & n4253;
  assign n4255 = n12046 & n4254;
  assign n4256 = n12046 | n4254;
  assign n4257 = ~n4255 & n4256;
  assign n4258 = x49 & x83;
  assign n4259 = n4257 & n4258;
  assign n4260 = n4257 | n4258;
  assign n4261 = ~n4259 & n4260;
  assign n4262 = n4238 & n4261;
  assign n4263 = n4238 | n4261;
  assign n4264 = ~n4262 & n4263;
  assign n4265 = x48 & x84;
  assign n4266 = n4264 & n4265;
  assign n4267 = n4264 | n4265;
  assign n4268 = ~n4266 & n4267;
  assign n12049 = n4238 | n4259;
  assign n12050 = (n4259 & n4261) | (n4259 & n12049) | (n4261 & n12049);
  assign n4272 = x53 & x80;
  assign n4273 = x52 & x81;
  assign n4274 = n4272 & n4273;
  assign n4275 = n4272 | n4273;
  assign n4276 = ~n4274 & n4275;
  assign n12051 = n4245 | n4247;
  assign n12053 = n4276 & n12051;
  assign n12054 = n4245 & n4276;
  assign n12055 = (n12048 & n12053) | (n12048 & n12054) | (n12053 & n12054);
  assign n12056 = n4276 | n12051;
  assign n12057 = n4245 | n4276;
  assign n12058 = (n12048 & n12056) | (n12048 & n12057) | (n12056 & n12057);
  assign n4279 = ~n12055 & n12058;
  assign n4280 = x51 & x82;
  assign n4281 = n4279 & n4280;
  assign n4282 = n4279 | n4280;
  assign n4283 = ~n4281 & n4282;
  assign n12059 = n4252 & n4283;
  assign n12060 = (n4255 & n4283) | (n4255 & n12059) | (n4283 & n12059);
  assign n12061 = n4252 | n4283;
  assign n12062 = n4255 | n12061;
  assign n4286 = ~n12060 & n12062;
  assign n4287 = x50 & x83;
  assign n4288 = n4286 & n4287;
  assign n4289 = n4286 | n4287;
  assign n4290 = ~n4288 & n4289;
  assign n4291 = n12050 & n4290;
  assign n4292 = n12050 | n4290;
  assign n4293 = ~n4291 & n4292;
  assign n4294 = x49 & x84;
  assign n4295 = n4293 & n4294;
  assign n4296 = n4293 | n4294;
  assign n4297 = ~n4295 & n4296;
  assign n4298 = n4266 & n4297;
  assign n4299 = n4266 | n4297;
  assign n4300 = ~n4298 & n4299;
  assign n4301 = x48 & x85;
  assign n4302 = n4300 & n4301;
  assign n4303 = n4300 | n4301;
  assign n4304 = ~n4302 & n4303;
  assign n12063 = n4266 | n4295;
  assign n12064 = (n4295 & n4297) | (n4295 & n12063) | (n4297 & n12063);
  assign n4306 = n4288 | n4291;
  assign n4309 = x54 & x80;
  assign n4310 = x53 & x81;
  assign n4311 = n4309 & n4310;
  assign n4312 = n4309 | n4310;
  assign n4313 = ~n4311 & n4312;
  assign n12065 = n4274 & n4313;
  assign n12066 = (n4313 & n12055) | (n4313 & n12065) | (n12055 & n12065);
  assign n12067 = n4274 | n4313;
  assign n12068 = n12055 | n12067;
  assign n4316 = ~n12066 & n12068;
  assign n4317 = x52 & x82;
  assign n4318 = n4316 & n4317;
  assign n4319 = n4316 | n4317;
  assign n4320 = ~n4318 & n4319;
  assign n12069 = n4281 & n4320;
  assign n12070 = (n4320 & n12060) | (n4320 & n12069) | (n12060 & n12069);
  assign n12071 = n4281 | n4320;
  assign n12072 = n12060 | n12071;
  assign n4323 = ~n12070 & n12072;
  assign n4324 = x51 & x83;
  assign n4325 = n4323 & n4324;
  assign n4326 = n4323 | n4324;
  assign n4327 = ~n4325 & n4326;
  assign n4328 = n4306 & n4327;
  assign n4329 = n4306 | n4327;
  assign n4330 = ~n4328 & n4329;
  assign n4331 = x50 & x84;
  assign n4332 = n4330 & n4331;
  assign n4333 = n4330 | n4331;
  assign n4334 = ~n4332 & n4333;
  assign n4335 = n12064 & n4334;
  assign n4336 = n12064 | n4334;
  assign n4337 = ~n4335 & n4336;
  assign n4338 = x49 & x85;
  assign n4339 = n4337 & n4338;
  assign n4340 = n4337 | n4338;
  assign n4341 = ~n4339 & n4340;
  assign n4342 = n4302 & n4341;
  assign n4343 = n4302 | n4341;
  assign n4344 = ~n4342 & n4343;
  assign n4345 = x48 & x86;
  assign n4346 = n4344 & n4345;
  assign n4347 = n4344 | n4345;
  assign n4348 = ~n4346 & n4347;
  assign n17674 = n4301 | n4338;
  assign n17675 = (n4300 & n4338) | (n4300 & n17674) | (n4338 & n17674);
  assign n15621 = (n4302 & n4337) | (n4302 & n17675) | (n4337 & n17675);
  assign n12074 = (n4339 & n4341) | (n4339 & n15621) | (n4341 & n15621);
  assign n12075 = n4332 | n12064;
  assign n12076 = (n4332 & n4334) | (n4332 & n12075) | (n4334 & n12075);
  assign n12077 = n4325 | n4327;
  assign n12078 = (n4306 & n4325) | (n4306 & n12077) | (n4325 & n12077);
  assign n4354 = x55 & x80;
  assign n4355 = x54 & x81;
  assign n4356 = n4354 & n4355;
  assign n4357 = n4354 | n4355;
  assign n4358 = ~n4356 & n4357;
  assign n15622 = n4274 | n4311;
  assign n15623 = (n4311 & n4313) | (n4311 & n15622) | (n4313 & n15622);
  assign n12082 = n4358 & n15623;
  assign n12080 = n4311 | n4313;
  assign n12083 = n4358 & n12080;
  assign n12084 = (n12055 & n12082) | (n12055 & n12083) | (n12082 & n12083);
  assign n12085 = n4358 | n15623;
  assign n12086 = n4358 | n12080;
  assign n12087 = (n12055 & n12085) | (n12055 & n12086) | (n12085 & n12086);
  assign n4361 = ~n12084 & n12087;
  assign n4362 = x53 & x82;
  assign n4363 = n4361 & n4362;
  assign n4364 = n4361 | n4362;
  assign n4365 = ~n4363 & n4364;
  assign n12088 = n4318 & n4365;
  assign n12089 = (n4365 & n12070) | (n4365 & n12088) | (n12070 & n12088);
  assign n12090 = n4318 | n4365;
  assign n12091 = n12070 | n12090;
  assign n4368 = ~n12089 & n12091;
  assign n4369 = x52 & x83;
  assign n4370 = n4368 & n4369;
  assign n4371 = n4368 | n4369;
  assign n4372 = ~n4370 & n4371;
  assign n4373 = n12078 & n4372;
  assign n4374 = n12078 | n4372;
  assign n4375 = ~n4373 & n4374;
  assign n4376 = x51 & x84;
  assign n4377 = n4375 & n4376;
  assign n4378 = n4375 | n4376;
  assign n4379 = ~n4377 & n4378;
  assign n4380 = n12076 & n4379;
  assign n4381 = n12076 | n4379;
  assign n4382 = ~n4380 & n4381;
  assign n4383 = x50 & x85;
  assign n4384 = n4382 & n4383;
  assign n4385 = n4382 | n4383;
  assign n4386 = ~n4384 & n4385;
  assign n4387 = n12074 & n4386;
  assign n4388 = n12074 | n4386;
  assign n4389 = ~n4387 & n4388;
  assign n4390 = x49 & x86;
  assign n4391 = n4389 & n4390;
  assign n4392 = n4389 | n4390;
  assign n4393 = ~n4391 & n4392;
  assign n4394 = n4346 & n4393;
  assign n4395 = n4346 | n4393;
  assign n4396 = ~n4394 & n4395;
  assign n4397 = x48 & x87;
  assign n4398 = n4396 & n4397;
  assign n4399 = n4396 | n4397;
  assign n4400 = ~n4398 & n4399;
  assign n12092 = n4346 | n4391;
  assign n12093 = (n4391 & n4393) | (n4391 & n12092) | (n4393 & n12092);
  assign n4402 = n4384 | n4387;
  assign n4403 = n4377 | n4380;
  assign n12094 = n4370 | n4372;
  assign n12095 = (n4370 & n12078) | (n4370 & n12094) | (n12078 & n12094);
  assign n4407 = x56 & x80;
  assign n4408 = x55 & x81;
  assign n4409 = n4407 & n4408;
  assign n4410 = n4407 | n4408;
  assign n4411 = ~n4409 & n4410;
  assign n12099 = n4356 & n4411;
  assign n15626 = (n4411 & n12083) | (n4411 & n12099) | (n12083 & n12099);
  assign n15627 = (n4411 & n12082) | (n4411 & n12099) | (n12082 & n12099);
  assign n15628 = (n12055 & n15626) | (n12055 & n15627) | (n15626 & n15627);
  assign n12101 = n4356 | n4411;
  assign n15629 = n12083 | n12101;
  assign n15630 = n12082 | n12101;
  assign n15631 = (n12055 & n15629) | (n12055 & n15630) | (n15629 & n15630);
  assign n4414 = ~n15628 & n15631;
  assign n4415 = x54 & x82;
  assign n4416 = n4414 & n4415;
  assign n4417 = n4414 | n4415;
  assign n4418 = ~n4416 & n4417;
  assign n12097 = n4363 | n4365;
  assign n15632 = n4418 & n12097;
  assign n15624 = n4318 | n4363;
  assign n15625 = (n4363 & n4365) | (n4363 & n15624) | (n4365 & n15624);
  assign n15633 = n4418 & n15625;
  assign n15634 = (n12070 & n15632) | (n12070 & n15633) | (n15632 & n15633);
  assign n15635 = n4418 | n12097;
  assign n15636 = n4418 | n15625;
  assign n15637 = (n12070 & n15635) | (n12070 & n15636) | (n15635 & n15636);
  assign n4421 = ~n15634 & n15637;
  assign n4422 = x53 & x83;
  assign n4423 = n4421 & n4422;
  assign n4424 = n4421 | n4422;
  assign n4425 = ~n4423 & n4424;
  assign n4426 = n12095 & n4425;
  assign n4427 = n12095 | n4425;
  assign n4428 = ~n4426 & n4427;
  assign n4429 = x52 & x84;
  assign n4430 = n4428 & n4429;
  assign n4431 = n4428 | n4429;
  assign n4432 = ~n4430 & n4431;
  assign n4433 = n4403 & n4432;
  assign n4434 = n4403 | n4432;
  assign n4435 = ~n4433 & n4434;
  assign n4436 = x51 & x85;
  assign n4437 = n4435 & n4436;
  assign n4438 = n4435 | n4436;
  assign n4439 = ~n4437 & n4438;
  assign n4440 = n4402 & n4439;
  assign n4441 = n4402 | n4439;
  assign n4442 = ~n4440 & n4441;
  assign n4443 = x50 & x86;
  assign n4444 = n4442 & n4443;
  assign n4445 = n4442 | n4443;
  assign n4446 = ~n4444 & n4445;
  assign n4447 = n12093 & n4446;
  assign n4448 = n12093 | n4446;
  assign n4449 = ~n4447 & n4448;
  assign n4450 = x49 & x87;
  assign n4451 = n4449 & n4450;
  assign n4452 = n4449 | n4450;
  assign n4453 = ~n4451 & n4452;
  assign n4454 = n4398 & n4453;
  assign n4455 = n4398 | n4453;
  assign n4456 = ~n4454 & n4455;
  assign n4457 = x48 & x88;
  assign n4458 = n4456 & n4457;
  assign n4459 = n4456 | n4457;
  assign n4460 = ~n4458 & n4459;
  assign n17676 = n4397 | n4450;
  assign n17677 = (n4396 & n4450) | (n4396 & n17676) | (n4450 & n17676);
  assign n15639 = (n4398 & n4449) | (n4398 & n17677) | (n4449 & n17677);
  assign n12104 = (n4451 & n4453) | (n4451 & n15639) | (n4453 & n15639);
  assign n12105 = n4444 | n12093;
  assign n12106 = (n4444 & n4446) | (n4444 & n12105) | (n4446 & n12105);
  assign n4463 = n4437 | n4440;
  assign n12107 = n4430 | n4432;
  assign n12108 = (n4403 & n4430) | (n4403 & n12107) | (n4430 & n12107);
  assign n12098 = (n12070 & n15625) | (n12070 & n12097) | (n15625 & n12097);
  assign n4468 = x57 & x80;
  assign n4469 = x56 & x81;
  assign n4470 = n4468 & n4469;
  assign n4471 = n4468 | n4469;
  assign n4472 = ~n4470 & n4471;
  assign n15640 = n4356 | n4409;
  assign n15641 = (n4409 & n4411) | (n4409 & n15640) | (n4411 & n15640);
  assign n12116 = n4472 & n15641;
  assign n12114 = n4409 | n4411;
  assign n12117 = n4472 & n12114;
  assign n15642 = (n12083 & n12116) | (n12083 & n12117) | (n12116 & n12117);
  assign n15643 = (n12082 & n12116) | (n12082 & n12117) | (n12116 & n12117);
  assign n15644 = (n12055 & n15642) | (n12055 & n15643) | (n15642 & n15643);
  assign n12119 = n4472 | n15641;
  assign n12120 = n4472 | n12114;
  assign n15645 = (n12083 & n12119) | (n12083 & n12120) | (n12119 & n12120);
  assign n15646 = (n12082 & n12119) | (n12082 & n12120) | (n12119 & n12120);
  assign n15647 = (n12055 & n15645) | (n12055 & n15646) | (n15645 & n15646);
  assign n4475 = ~n15644 & n15647;
  assign n4476 = x55 & x82;
  assign n4477 = n4475 & n4476;
  assign n4478 = n4475 | n4476;
  assign n4479 = ~n4477 & n4478;
  assign n12111 = n4416 | n4418;
  assign n12122 = n4479 & n12111;
  assign n12123 = n4416 & n4479;
  assign n12124 = (n12098 & n12122) | (n12098 & n12123) | (n12122 & n12123);
  assign n12125 = n4479 | n12111;
  assign n12126 = n4416 | n4479;
  assign n12127 = (n12098 & n12125) | (n12098 & n12126) | (n12125 & n12126);
  assign n4482 = ~n12124 & n12127;
  assign n4483 = x54 & x83;
  assign n4484 = n4482 & n4483;
  assign n4485 = n4482 | n4483;
  assign n4486 = ~n4484 & n4485;
  assign n12109 = n4423 | n4425;
  assign n15648 = n4486 & n12109;
  assign n15649 = n4423 & n4486;
  assign n15650 = (n12095 & n15648) | (n12095 & n15649) | (n15648 & n15649);
  assign n15651 = n4486 | n12109;
  assign n15652 = n4423 | n4486;
  assign n15653 = (n12095 & n15651) | (n12095 & n15652) | (n15651 & n15652);
  assign n4489 = ~n15650 & n15653;
  assign n4490 = x53 & x84;
  assign n4491 = n4489 & n4490;
  assign n4492 = n4489 | n4490;
  assign n4493 = ~n4491 & n4492;
  assign n4494 = n12108 & n4493;
  assign n4495 = n12108 | n4493;
  assign n4496 = ~n4494 & n4495;
  assign n4497 = x52 & x85;
  assign n4498 = n4496 & n4497;
  assign n4499 = n4496 | n4497;
  assign n4500 = ~n4498 & n4499;
  assign n4501 = n4463 & n4500;
  assign n4502 = n4463 | n4500;
  assign n4503 = ~n4501 & n4502;
  assign n4504 = x51 & x86;
  assign n4505 = n4503 & n4504;
  assign n4506 = n4503 | n4504;
  assign n4507 = ~n4505 & n4506;
  assign n4508 = n12106 & n4507;
  assign n4509 = n12106 | n4507;
  assign n4510 = ~n4508 & n4509;
  assign n4511 = x50 & x87;
  assign n4512 = n4510 & n4511;
  assign n4513 = n4510 | n4511;
  assign n4514 = ~n4512 & n4513;
  assign n4515 = n12104 & n4514;
  assign n4516 = n12104 | n4514;
  assign n4517 = ~n4515 & n4516;
  assign n4518 = x49 & x88;
  assign n4519 = n4517 & n4518;
  assign n4520 = n4517 | n4518;
  assign n4521 = ~n4519 & n4520;
  assign n4522 = n4458 & n4521;
  assign n4523 = n4458 | n4521;
  assign n4524 = ~n4522 & n4523;
  assign n4525 = x48 & x89;
  assign n4526 = n4524 & n4525;
  assign n4527 = n4524 | n4525;
  assign n4528 = ~n4526 & n4527;
  assign n17678 = n4457 | n4518;
  assign n17679 = (n4456 & n4518) | (n4456 & n17678) | (n4518 & n17678);
  assign n15655 = (n4458 & n4517) | (n4458 & n17679) | (n4517 & n17679);
  assign n12129 = (n4519 & n4521) | (n4519 & n15655) | (n4521 & n15655);
  assign n12130 = n4512 | n12104;
  assign n12131 = (n4512 & n4514) | (n4512 & n12130) | (n4514 & n12130);
  assign n12132 = n4505 | n12106;
  assign n12133 = (n4505 & n4507) | (n4505 & n12132) | (n4507 & n12132);
  assign n12134 = n4498 | n4500;
  assign n12135 = (n4463 & n4498) | (n4463 & n12134) | (n4498 & n12134);
  assign n12110 = (n4423 & n12095) | (n4423 & n12109) | (n12095 & n12109);
  assign n15656 = n4470 | n4472;
  assign n15657 = (n4470 & n15641) | (n4470 & n15656) | (n15641 & n15656);
  assign n15658 = (n4470 & n12114) | (n4470 & n15656) | (n12114 & n15656);
  assign n15659 = (n12083 & n15657) | (n12083 & n15658) | (n15657 & n15658);
  assign n15660 = (n12082 & n15657) | (n12082 & n15658) | (n15657 & n15658);
  assign n15661 = (n12055 & n15659) | (n12055 & n15660) | (n15659 & n15660);
  assign n4537 = x58 & x80;
  assign n4538 = x57 & x81;
  assign n4539 = n4537 & n4538;
  assign n4540 = n4537 | n4538;
  assign n4541 = ~n4539 & n4540;
  assign n4542 = n15661 & n4541;
  assign n4543 = n15661 | n4541;
  assign n4544 = ~n4542 & n4543;
  assign n4545 = x56 & x82;
  assign n4546 = n4544 & n4545;
  assign n4547 = n4544 | n4545;
  assign n4548 = ~n4546 & n4547;
  assign n12143 = n4477 & n4548;
  assign n15662 = (n4548 & n12122) | (n4548 & n12143) | (n12122 & n12143);
  assign n15663 = (n4548 & n12123) | (n4548 & n12143) | (n12123 & n12143);
  assign n15664 = (n12098 & n15662) | (n12098 & n15663) | (n15662 & n15663);
  assign n12145 = n4477 | n4548;
  assign n15665 = n12122 | n12145;
  assign n15666 = n12123 | n12145;
  assign n15667 = (n12098 & n15665) | (n12098 & n15666) | (n15665 & n15666);
  assign n4551 = ~n15664 & n15667;
  assign n4552 = x55 & x83;
  assign n4553 = n4551 & n4552;
  assign n4554 = n4551 | n4552;
  assign n4555 = ~n4553 & n4554;
  assign n12138 = n4484 | n4486;
  assign n12147 = n4555 & n12138;
  assign n12148 = n4484 & n4555;
  assign n12149 = (n12110 & n12147) | (n12110 & n12148) | (n12147 & n12148);
  assign n12150 = n4555 | n12138;
  assign n12151 = n4484 | n4555;
  assign n12152 = (n12110 & n12150) | (n12110 & n12151) | (n12150 & n12151);
  assign n4558 = ~n12149 & n12152;
  assign n4559 = x54 & x84;
  assign n4560 = n4558 & n4559;
  assign n4561 = n4558 | n4559;
  assign n4562 = ~n4560 & n4561;
  assign n12136 = n4491 | n4493;
  assign n15668 = n4562 & n12136;
  assign n15669 = n4491 & n4562;
  assign n15670 = (n12108 & n15668) | (n12108 & n15669) | (n15668 & n15669);
  assign n15671 = n4562 | n12136;
  assign n15672 = n4491 | n4562;
  assign n15673 = (n12108 & n15671) | (n12108 & n15672) | (n15671 & n15672);
  assign n4565 = ~n15670 & n15673;
  assign n4566 = x53 & x85;
  assign n4567 = n4565 & n4566;
  assign n4568 = n4565 | n4566;
  assign n4569 = ~n4567 & n4568;
  assign n4570 = n12135 & n4569;
  assign n4571 = n12135 | n4569;
  assign n4572 = ~n4570 & n4571;
  assign n4573 = x52 & x86;
  assign n4574 = n4572 & n4573;
  assign n4575 = n4572 | n4573;
  assign n4576 = ~n4574 & n4575;
  assign n4577 = n12133 & n4576;
  assign n4578 = n12133 | n4576;
  assign n4579 = ~n4577 & n4578;
  assign n4580 = x51 & x87;
  assign n4581 = n4579 & n4580;
  assign n4582 = n4579 | n4580;
  assign n4583 = ~n4581 & n4582;
  assign n4584 = n12131 & n4583;
  assign n4585 = n12131 | n4583;
  assign n4586 = ~n4584 & n4585;
  assign n4587 = x50 & x88;
  assign n4588 = n4586 & n4587;
  assign n4589 = n4586 | n4587;
  assign n4590 = ~n4588 & n4589;
  assign n4591 = n12129 & n4590;
  assign n4592 = n12129 | n4590;
  assign n4593 = ~n4591 & n4592;
  assign n4594 = x49 & x89;
  assign n4595 = n4593 & n4594;
  assign n4596 = n4593 | n4594;
  assign n4597 = ~n4595 & n4596;
  assign n4598 = n4526 & n4597;
  assign n4599 = n4526 | n4597;
  assign n4600 = ~n4598 & n4599;
  assign n4601 = x48 & x90;
  assign n4602 = n4600 & n4601;
  assign n4603 = n4600 | n4601;
  assign n4604 = ~n4602 & n4603;
  assign n12153 = n4526 | n4595;
  assign n12154 = (n4595 & n4597) | (n4595 & n12153) | (n4597 & n12153);
  assign n4606 = n4588 | n4591;
  assign n4607 = n4581 | n4584;
  assign n12137 = (n4491 & n12108) | (n4491 & n12136) | (n12108 & n12136);
  assign n12160 = n4546 | n4548;
  assign n15674 = n4477 | n4546;
  assign n15675 = (n4546 & n4548) | (n4546 & n15674) | (n4548 & n15674);
  assign n15676 = (n12122 & n12160) | (n12122 & n15675) | (n12160 & n15675);
  assign n15677 = (n12123 & n12160) | (n12123 & n15675) | (n12160 & n15675);
  assign n15678 = (n12098 & n15676) | (n12098 & n15677) | (n15676 & n15677);
  assign n4614 = x59 & x80;
  assign n4615 = x58 & x81;
  assign n4616 = n4614 & n4615;
  assign n4617 = n4614 | n4615;
  assign n4618 = ~n4616 & n4617;
  assign n12162 = n4539 | n4541;
  assign n12164 = n4618 & n12162;
  assign n12165 = n4539 & n4618;
  assign n12166 = (n15661 & n12164) | (n15661 & n12165) | (n12164 & n12165);
  assign n12167 = n4618 | n12162;
  assign n12168 = n4539 | n4618;
  assign n12169 = (n15661 & n12167) | (n15661 & n12168) | (n12167 & n12168);
  assign n4621 = ~n12166 & n12169;
  assign n4622 = x57 & x82;
  assign n4623 = n4621 & n4622;
  assign n4624 = n4621 | n4622;
  assign n4625 = ~n4623 & n4624;
  assign n4626 = n15678 & n4625;
  assign n4627 = n15678 | n4625;
  assign n4628 = ~n4626 & n4627;
  assign n4629 = x56 & x83;
  assign n4630 = n4628 & n4629;
  assign n4631 = n4628 | n4629;
  assign n4632 = ~n4630 & n4631;
  assign n12170 = n4553 & n4632;
  assign n12171 = (n4632 & n12149) | (n4632 & n12170) | (n12149 & n12170);
  assign n12172 = n4553 | n4632;
  assign n12173 = n12149 | n12172;
  assign n4635 = ~n12171 & n12173;
  assign n4636 = x55 & x84;
  assign n4637 = n4635 & n4636;
  assign n4638 = n4635 | n4636;
  assign n4639 = ~n4637 & n4638;
  assign n12157 = n4560 | n4562;
  assign n12174 = n4639 & n12157;
  assign n12175 = n4560 & n4639;
  assign n12176 = (n12137 & n12174) | (n12137 & n12175) | (n12174 & n12175);
  assign n12177 = n4639 | n12157;
  assign n12178 = n4560 | n4639;
  assign n12179 = (n12137 & n12177) | (n12137 & n12178) | (n12177 & n12178);
  assign n4642 = ~n12176 & n12179;
  assign n4643 = x54 & x85;
  assign n4644 = n4642 & n4643;
  assign n4645 = n4642 | n4643;
  assign n4646 = ~n4644 & n4645;
  assign n12155 = n4567 | n4569;
  assign n15679 = n4646 & n12155;
  assign n15680 = n4567 & n4646;
  assign n15681 = (n12135 & n15679) | (n12135 & n15680) | (n15679 & n15680);
  assign n15682 = n4646 | n12155;
  assign n15683 = n4567 | n4646;
  assign n15684 = (n12135 & n15682) | (n12135 & n15683) | (n15682 & n15683);
  assign n4649 = ~n15681 & n15684;
  assign n4650 = x53 & x86;
  assign n4651 = n4649 & n4650;
  assign n4652 = n4649 | n4650;
  assign n4653 = ~n4651 & n4652;
  assign n15685 = n4574 & n4653;
  assign n15686 = (n4577 & n4653) | (n4577 & n15685) | (n4653 & n15685);
  assign n15687 = n4574 | n4653;
  assign n15688 = n4577 | n15687;
  assign n4656 = ~n15686 & n15688;
  assign n4657 = x52 & x87;
  assign n4658 = n4656 & n4657;
  assign n4659 = n4656 | n4657;
  assign n4660 = ~n4658 & n4659;
  assign n4661 = n4607 & n4660;
  assign n4662 = n4607 | n4660;
  assign n4663 = ~n4661 & n4662;
  assign n4664 = x51 & x88;
  assign n4665 = n4663 & n4664;
  assign n4666 = n4663 | n4664;
  assign n4667 = ~n4665 & n4666;
  assign n4668 = n4606 & n4667;
  assign n4669 = n4606 | n4667;
  assign n4670 = ~n4668 & n4669;
  assign n4671 = x50 & x89;
  assign n4672 = n4670 & n4671;
  assign n4673 = n4670 | n4671;
  assign n4674 = ~n4672 & n4673;
  assign n4675 = n12154 & n4674;
  assign n4676 = n12154 | n4674;
  assign n4677 = ~n4675 & n4676;
  assign n4678 = x49 & x90;
  assign n4679 = n4677 & n4678;
  assign n4680 = n4677 | n4678;
  assign n4681 = ~n4679 & n4680;
  assign n4682 = n4602 & n4681;
  assign n4683 = n4602 | n4681;
  assign n4684 = ~n4682 & n4683;
  assign n4685 = x48 & x91;
  assign n4686 = n4684 & n4685;
  assign n4687 = n4684 | n4685;
  assign n4688 = ~n4686 & n4687;
  assign n17680 = n4601 | n4678;
  assign n17681 = (n4600 & n4678) | (n4600 & n17680) | (n4678 & n17680);
  assign n15690 = (n4602 & n4677) | (n4602 & n17681) | (n4677 & n17681);
  assign n12181 = (n4679 & n4681) | (n4679 & n15690) | (n4681 & n15690);
  assign n12182 = n4672 | n12154;
  assign n12183 = (n4672 & n4674) | (n4672 & n12182) | (n4674 & n12182);
  assign n4691 = n4665 | n4668;
  assign n15691 = n4658 | n4660;
  assign n15692 = (n4607 & n4658) | (n4607 & n15691) | (n4658 & n15691);
  assign n4608 = n4574 | n4577;
  assign n12156 = (n4567 & n12135) | (n4567 & n12155) | (n12135 & n12155);
  assign n4699 = x60 & x80;
  assign n4700 = x59 & x81;
  assign n4701 = n4699 & n4700;
  assign n4702 = n4699 | n4700;
  assign n4703 = ~n4701 & n4702;
  assign n15693 = n4616 | n4618;
  assign n15694 = (n4616 & n12162) | (n4616 & n15693) | (n12162 & n15693);
  assign n12193 = n4703 & n15694;
  assign n15695 = n4539 | n4616;
  assign n15696 = (n4616 & n4618) | (n4616 & n15695) | (n4618 & n15695);
  assign n12194 = n4703 & n15696;
  assign n12195 = (n15661 & n12193) | (n15661 & n12194) | (n12193 & n12194);
  assign n12196 = n4703 | n15694;
  assign n12197 = n4703 | n15696;
  assign n12198 = (n15661 & n12196) | (n15661 & n12197) | (n12196 & n12197);
  assign n4706 = ~n12195 & n12198;
  assign n4707 = x58 & x82;
  assign n4708 = n4706 & n4707;
  assign n4709 = n4706 | n4707;
  assign n4710 = ~n4708 & n4709;
  assign n12188 = n4623 | n4625;
  assign n12199 = n4710 & n12188;
  assign n12200 = n4623 & n4710;
  assign n12201 = (n15678 & n12199) | (n15678 & n12200) | (n12199 & n12200);
  assign n12202 = n4710 | n12188;
  assign n12203 = n4623 | n4710;
  assign n12204 = (n15678 & n12202) | (n15678 & n12203) | (n12202 & n12203);
  assign n4713 = ~n12201 & n12204;
  assign n4714 = x57 & x83;
  assign n4715 = n4713 & n4714;
  assign n4716 = n4713 | n4714;
  assign n4717 = ~n4715 & n4716;
  assign n12205 = n4630 & n4717;
  assign n15697 = (n4717 & n12170) | (n4717 & n12205) | (n12170 & n12205);
  assign n15698 = (n4632 & n4717) | (n4632 & n12205) | (n4717 & n12205);
  assign n15699 = (n12149 & n15697) | (n12149 & n15698) | (n15697 & n15698);
  assign n12207 = n4630 | n4717;
  assign n15700 = n12170 | n12207;
  assign n15701 = n4632 | n12207;
  assign n15702 = (n12149 & n15700) | (n12149 & n15701) | (n15700 & n15701);
  assign n4720 = ~n15699 & n15702;
  assign n4721 = x56 & x84;
  assign n4722 = n4720 & n4721;
  assign n4723 = n4720 | n4721;
  assign n4724 = ~n4722 & n4723;
  assign n12209 = n4637 & n4724;
  assign n12210 = (n4724 & n12176) | (n4724 & n12209) | (n12176 & n12209);
  assign n12211 = n4637 | n4724;
  assign n12212 = n12176 | n12211;
  assign n4727 = ~n12210 & n12212;
  assign n4728 = x55 & x85;
  assign n4729 = n4727 & n4728;
  assign n4730 = n4727 | n4728;
  assign n4731 = ~n4729 & n4730;
  assign n12186 = n4644 | n4646;
  assign n12213 = n4731 & n12186;
  assign n12214 = n4644 & n4731;
  assign n12215 = (n12156 & n12213) | (n12156 & n12214) | (n12213 & n12214);
  assign n12216 = n4731 | n12186;
  assign n12217 = n4644 | n4731;
  assign n12218 = (n12156 & n12216) | (n12156 & n12217) | (n12216 & n12217);
  assign n4734 = ~n12215 & n12218;
  assign n4735 = x54 & x86;
  assign n4736 = n4734 & n4735;
  assign n4737 = n4734 | n4735;
  assign n4738 = ~n4736 & n4737;
  assign n12184 = n4651 | n4653;
  assign n15703 = n4738 & n12184;
  assign n15704 = n4651 & n4738;
  assign n15705 = (n4608 & n15703) | (n4608 & n15704) | (n15703 & n15704);
  assign n15706 = n4738 | n12184;
  assign n15707 = n4651 | n4738;
  assign n15708 = (n4608 & n15706) | (n4608 & n15707) | (n15706 & n15707);
  assign n4741 = ~n15705 & n15708;
  assign n4742 = x53 & x87;
  assign n4743 = n4741 & n4742;
  assign n4744 = n4741 | n4742;
  assign n4745 = ~n4743 & n4744;
  assign n4746 = n15692 & n4745;
  assign n4747 = n15692 | n4745;
  assign n4748 = ~n4746 & n4747;
  assign n4749 = x52 & x88;
  assign n4750 = n4748 & n4749;
  assign n4751 = n4748 | n4749;
  assign n4752 = ~n4750 & n4751;
  assign n4753 = n4691 & n4752;
  assign n4754 = n4691 | n4752;
  assign n4755 = ~n4753 & n4754;
  assign n4756 = x51 & x89;
  assign n4757 = n4755 & n4756;
  assign n4758 = n4755 | n4756;
  assign n4759 = ~n4757 & n4758;
  assign n4760 = n12183 & n4759;
  assign n4761 = n12183 | n4759;
  assign n4762 = ~n4760 & n4761;
  assign n4763 = x50 & x90;
  assign n4764 = n4762 & n4763;
  assign n4765 = n4762 | n4763;
  assign n4766 = ~n4764 & n4765;
  assign n4767 = n12181 & n4766;
  assign n4768 = n12181 | n4766;
  assign n4769 = ~n4767 & n4768;
  assign n4770 = x49 & x91;
  assign n4771 = n4769 & n4770;
  assign n4772 = n4769 | n4770;
  assign n4773 = ~n4771 & n4772;
  assign n4774 = n4686 & n4773;
  assign n4775 = n4686 | n4773;
  assign n4776 = ~n4774 & n4775;
  assign n4777 = x48 & x92;
  assign n4778 = n4776 & n4777;
  assign n4779 = n4776 | n4777;
  assign n4780 = ~n4778 & n4779;
  assign n17682 = n4685 | n4770;
  assign n17683 = (n4684 & n4770) | (n4684 & n17682) | (n4770 & n17682);
  assign n15710 = (n4686 & n4769) | (n4686 & n17683) | (n4769 & n17683);
  assign n12220 = (n4771 & n4773) | (n4771 & n15710) | (n4773 & n15710);
  assign n12221 = n4764 | n12181;
  assign n12222 = (n4764 & n4766) | (n4764 & n12221) | (n4766 & n12221);
  assign n12223 = n4757 | n12183;
  assign n12224 = (n4757 & n4759) | (n4757 & n12223) | (n4759 & n12223);
  assign n15711 = n4750 | n4752;
  assign n15712 = (n4691 & n4750) | (n4691 & n15711) | (n4750 & n15711);
  assign n12225 = n4743 | n4745;
  assign n12226 = (n15692 & n4743) | (n15692 & n12225) | (n4743 & n12225);
  assign n12185 = (n4608 & n4651) | (n4608 & n12184) | (n4651 & n12184);
  assign n12230 = n4715 | n4717;
  assign n15713 = n4630 | n4715;
  assign n15714 = (n4715 & n4717) | (n4715 & n15713) | (n4717 & n15713);
  assign n15715 = (n12170 & n12230) | (n12170 & n15714) | (n12230 & n15714);
  assign n15716 = (n4632 & n12230) | (n4632 & n15714) | (n12230 & n15714);
  assign n15717 = (n12149 & n15715) | (n12149 & n15716) | (n15715 & n15716);
  assign n4792 = x61 & x80;
  assign n4793 = x60 & x81;
  assign n4794 = n4792 & n4793;
  assign n4795 = n4792 | n4793;
  assign n4796 = ~n4794 & n4795;
  assign n15722 = n4701 | n4703;
  assign n17684 = n4796 & n15722;
  assign n17685 = n4701 & n4796;
  assign n17686 = (n15694 & n17684) | (n15694 & n17685) | (n17684 & n17685);
  assign n15724 = (n4701 & n15696) | (n4701 & n15722) | (n15696 & n15722);
  assign n15726 = n4796 & n15724;
  assign n15727 = (n15661 & n17686) | (n15661 & n15726) | (n17686 & n15726);
  assign n17687 = n4796 | n15722;
  assign n17688 = n4701 | n4796;
  assign n17689 = (n15694 & n17687) | (n15694 & n17688) | (n17687 & n17688);
  assign n15729 = n4796 | n15724;
  assign n15730 = (n15661 & n17689) | (n15661 & n15729) | (n17689 & n15729);
  assign n4799 = ~n15727 & n15730;
  assign n4800 = x59 & x82;
  assign n4801 = n4799 & n4800;
  assign n4802 = n4799 | n4800;
  assign n4803 = ~n4801 & n4802;
  assign n15718 = n4708 | n4710;
  assign n15719 = (n4708 & n12188) | (n4708 & n15718) | (n12188 & n15718);
  assign n15731 = n4803 & n15719;
  assign n15720 = n4623 | n4708;
  assign n15721 = (n4708 & n4710) | (n4708 & n15720) | (n4710 & n15720);
  assign n15732 = n4803 & n15721;
  assign n15733 = (n15678 & n15731) | (n15678 & n15732) | (n15731 & n15732);
  assign n15734 = n4803 | n15719;
  assign n15735 = n4803 | n15721;
  assign n15736 = (n15678 & n15734) | (n15678 & n15735) | (n15734 & n15735);
  assign n4806 = ~n15733 & n15736;
  assign n4807 = x58 & x83;
  assign n4808 = n4806 & n4807;
  assign n4809 = n4806 | n4807;
  assign n4810 = ~n4808 & n4809;
  assign n4811 = n15717 & n4810;
  assign n4812 = n15717 | n4810;
  assign n4813 = ~n4811 & n4812;
  assign n4814 = x57 & x84;
  assign n4815 = n4813 & n4814;
  assign n4816 = n4813 | n4814;
  assign n4817 = ~n4815 & n4816;
  assign n12238 = n4722 & n4817;
  assign n12239 = (n4817 & n12210) | (n4817 & n12238) | (n12210 & n12238);
  assign n12240 = n4722 | n4817;
  assign n12241 = n12210 | n12240;
  assign n4820 = ~n12239 & n12241;
  assign n4821 = x56 & x85;
  assign n4822 = n4820 & n4821;
  assign n4823 = n4820 | n4821;
  assign n4824 = ~n4822 & n4823;
  assign n12242 = n4729 & n4824;
  assign n12243 = (n4824 & n12215) | (n4824 & n12242) | (n12215 & n12242);
  assign n12244 = n4729 | n4824;
  assign n12245 = n12215 | n12244;
  assign n4827 = ~n12243 & n12245;
  assign n4828 = x55 & x86;
  assign n4829 = n4827 & n4828;
  assign n4830 = n4827 | n4828;
  assign n4831 = ~n4829 & n4830;
  assign n12227 = n4736 | n4738;
  assign n12246 = n4831 & n12227;
  assign n12247 = n4736 & n4831;
  assign n12248 = (n12185 & n12246) | (n12185 & n12247) | (n12246 & n12247);
  assign n12249 = n4831 | n12227;
  assign n12250 = n4736 | n4831;
  assign n12251 = (n12185 & n12249) | (n12185 & n12250) | (n12249 & n12250);
  assign n4834 = ~n12248 & n12251;
  assign n4835 = x54 & x87;
  assign n4836 = n4834 & n4835;
  assign n4837 = n4834 | n4835;
  assign n4838 = ~n4836 & n4837;
  assign n4839 = n12226 & n4838;
  assign n4840 = n12226 | n4838;
  assign n4841 = ~n4839 & n4840;
  assign n4842 = x53 & x88;
  assign n4843 = n4841 & n4842;
  assign n4844 = n4841 | n4842;
  assign n4845 = ~n4843 & n4844;
  assign n4846 = n15712 & n4845;
  assign n4847 = n15712 | n4845;
  assign n4848 = ~n4846 & n4847;
  assign n4849 = x52 & x89;
  assign n4850 = n4848 & n4849;
  assign n4851 = n4848 | n4849;
  assign n4852 = ~n4850 & n4851;
  assign n4853 = n12224 & n4852;
  assign n4854 = n12224 | n4852;
  assign n4855 = ~n4853 & n4854;
  assign n4856 = x51 & x90;
  assign n4857 = n4855 & n4856;
  assign n4858 = n4855 | n4856;
  assign n4859 = ~n4857 & n4858;
  assign n4860 = n12222 & n4859;
  assign n4861 = n12222 | n4859;
  assign n4862 = ~n4860 & n4861;
  assign n4863 = x50 & x91;
  assign n4864 = n4862 & n4863;
  assign n4865 = n4862 | n4863;
  assign n4866 = ~n4864 & n4865;
  assign n4867 = n12220 & n4866;
  assign n4868 = n12220 | n4866;
  assign n4869 = ~n4867 & n4868;
  assign n4870 = x49 & x92;
  assign n4871 = n4869 & n4870;
  assign n4872 = n4869 | n4870;
  assign n4873 = ~n4871 & n4872;
  assign n4874 = n4778 & n4873;
  assign n4875 = n4778 | n4873;
  assign n4876 = ~n4874 & n4875;
  assign n4877 = x48 & x93;
  assign n4878 = n4876 & n4877;
  assign n4879 = n4876 | n4877;
  assign n4880 = ~n4878 & n4879;
  assign n12252 = n4778 | n4871;
  assign n12253 = (n4871 & n4873) | (n4871 & n12252) | (n4873 & n12252);
  assign n12254 = n4864 | n12220;
  assign n12255 = (n4864 & n4866) | (n4864 & n12254) | (n4866 & n12254);
  assign n12256 = n4857 | n12222;
  assign n12257 = (n4857 & n4859) | (n4857 & n12256) | (n4859 & n12256);
  assign n12258 = n4850 | n12224;
  assign n12259 = (n4850 & n4852) | (n4850 & n12258) | (n4852 & n12258);
  assign n12260 = n4843 | n4845;
  assign n12261 = (n15712 & n4843) | (n15712 & n12260) | (n4843 & n12260);
  assign n4893 = x62 & x80;
  assign n4894 = x61 & x81;
  assign n4895 = n4893 & n4894;
  assign n4896 = n4893 | n4894;
  assign n4897 = ~n4895 & n4896;
  assign n12268 = n4794 | n4796;
  assign n12270 = n4897 & n12268;
  assign n12271 = n4794 & n4897;
  assign n15723 = (n4701 & n15694) | (n4701 & n15722) | (n15694 & n15722);
  assign n15737 = (n12270 & n12271) | (n12270 & n15723) | (n12271 & n15723);
  assign n15738 = (n12270 & n12271) | (n12270 & n15724) | (n12271 & n15724);
  assign n15739 = (n15661 & n15737) | (n15661 & n15738) | (n15737 & n15738);
  assign n12273 = n4897 | n12268;
  assign n12274 = n4794 | n4897;
  assign n15740 = (n12273 & n12274) | (n12273 & n15723) | (n12274 & n15723);
  assign n15741 = (n12273 & n12274) | (n12273 & n15724) | (n12274 & n15724);
  assign n15742 = (n15661 & n15740) | (n15661 & n15741) | (n15740 & n15741);
  assign n4900 = ~n15739 & n15742;
  assign n4901 = x60 & x82;
  assign n4902 = n4900 & n4901;
  assign n4903 = n4900 | n4901;
  assign n4904 = ~n4902 & n4903;
  assign n12266 = n4801 | n4803;
  assign n12276 = n4904 & n12266;
  assign n12277 = n4801 & n4904;
  assign n15743 = (n12276 & n12277) | (n12276 & n15719) | (n12277 & n15719);
  assign n15744 = (n12276 & n12277) | (n12276 & n15721) | (n12277 & n15721);
  assign n15745 = (n15678 & n15743) | (n15678 & n15744) | (n15743 & n15744);
  assign n12279 = n4904 | n12266;
  assign n12280 = n4801 | n4904;
  assign n15746 = (n12279 & n12280) | (n12279 & n15719) | (n12280 & n15719);
  assign n15747 = (n12279 & n12280) | (n12279 & n15721) | (n12280 & n15721);
  assign n15748 = (n15678 & n15746) | (n15678 & n15747) | (n15746 & n15747);
  assign n4907 = ~n15745 & n15748;
  assign n4908 = x59 & x83;
  assign n4909 = n4907 & n4908;
  assign n4910 = n4907 | n4908;
  assign n4911 = ~n4909 & n4910;
  assign n12264 = n4808 | n4810;
  assign n12282 = n4911 & n12264;
  assign n12283 = n4808 & n4911;
  assign n12284 = (n15717 & n12282) | (n15717 & n12283) | (n12282 & n12283);
  assign n12285 = n4911 | n12264;
  assign n12286 = n4808 | n4911;
  assign n12287 = (n15717 & n12285) | (n15717 & n12286) | (n12285 & n12286);
  assign n4914 = ~n12284 & n12287;
  assign n4915 = x58 & x84;
  assign n4916 = n4914 & n4915;
  assign n4917 = n4914 | n4915;
  assign n4918 = ~n4916 & n4917;
  assign n12288 = n4815 & n4918;
  assign n15749 = (n4918 & n12238) | (n4918 & n12288) | (n12238 & n12288);
  assign n15750 = (n4817 & n4918) | (n4817 & n12288) | (n4918 & n12288);
  assign n15751 = (n12210 & n15749) | (n12210 & n15750) | (n15749 & n15750);
  assign n12290 = n4815 | n4918;
  assign n15752 = n12238 | n12290;
  assign n15753 = n4817 | n12290;
  assign n15754 = (n12210 & n15752) | (n12210 & n15753) | (n15752 & n15753);
  assign n4921 = ~n15751 & n15754;
  assign n4922 = x57 & x85;
  assign n4923 = n4921 & n4922;
  assign n4924 = n4921 | n4922;
  assign n4925 = ~n4923 & n4924;
  assign n12292 = n4822 & n4925;
  assign n12293 = (n4925 & n12243) | (n4925 & n12292) | (n12243 & n12292);
  assign n12294 = n4822 | n4925;
  assign n12295 = n12243 | n12294;
  assign n4928 = ~n12293 & n12295;
  assign n4929 = x56 & x86;
  assign n4930 = n4928 & n4929;
  assign n4931 = n4928 | n4929;
  assign n4932 = ~n4930 & n4931;
  assign n12296 = n4829 & n4932;
  assign n12297 = (n4932 & n12248) | (n4932 & n12296) | (n12248 & n12296);
  assign n12298 = n4829 | n4932;
  assign n12299 = n12248 | n12298;
  assign n4935 = ~n12297 & n12299;
  assign n4936 = x55 & x87;
  assign n4937 = n4935 & n4936;
  assign n4938 = n4935 | n4936;
  assign n4939 = ~n4937 & n4938;
  assign n12262 = n4836 | n4838;
  assign n12300 = n4939 & n12262;
  assign n12301 = n4836 & n4939;
  assign n12302 = (n12226 & n12300) | (n12226 & n12301) | (n12300 & n12301);
  assign n12303 = n4939 | n12262;
  assign n12304 = n4836 | n4939;
  assign n12305 = (n12226 & n12303) | (n12226 & n12304) | (n12303 & n12304);
  assign n4942 = ~n12302 & n12305;
  assign n4943 = x54 & x88;
  assign n4944 = n4942 & n4943;
  assign n4945 = n4942 | n4943;
  assign n4946 = ~n4944 & n4945;
  assign n4947 = n12261 & n4946;
  assign n4948 = n12261 | n4946;
  assign n4949 = ~n4947 & n4948;
  assign n4950 = x53 & x89;
  assign n4951 = n4949 & n4950;
  assign n4952 = n4949 | n4950;
  assign n4953 = ~n4951 & n4952;
  assign n4954 = n12259 & n4953;
  assign n4955 = n12259 | n4953;
  assign n4956 = ~n4954 & n4955;
  assign n4957 = x52 & x90;
  assign n4958 = n4956 & n4957;
  assign n4959 = n4956 | n4957;
  assign n4960 = ~n4958 & n4959;
  assign n4961 = n12257 & n4960;
  assign n4962 = n12257 | n4960;
  assign n4963 = ~n4961 & n4962;
  assign n4964 = x51 & x91;
  assign n4965 = n4963 & n4964;
  assign n4966 = n4963 | n4964;
  assign n4967 = ~n4965 & n4966;
  assign n4968 = n12255 & n4967;
  assign n4969 = n12255 | n4967;
  assign n4970 = ~n4968 & n4969;
  assign n4971 = x50 & x92;
  assign n4972 = n4970 & n4971;
  assign n4973 = n4970 | n4971;
  assign n4974 = ~n4972 & n4973;
  assign n4975 = n12253 & n4974;
  assign n4976 = n12253 | n4974;
  assign n4977 = ~n4975 & n4976;
  assign n4978 = x49 & x93;
  assign n4979 = n4977 & n4978;
  assign n4980 = n4977 | n4978;
  assign n4981 = ~n4979 & n4980;
  assign n4982 = n4878 & n4981;
  assign n4983 = n4878 | n4981;
  assign n4984 = ~n4982 & n4983;
  assign n4985 = x48 & x94;
  assign n4986 = n4984 & n4985;
  assign n4987 = n4984 | n4985;
  assign n4988 = ~n4986 & n4987;
  assign n17690 = n4877 | n4978;
  assign n17691 = (n4876 & n4978) | (n4876 & n17690) | (n4978 & n17690);
  assign n15756 = (n4878 & n4977) | (n4878 & n17691) | (n4977 & n17691);
  assign n12307 = (n4979 & n4981) | (n4979 & n15756) | (n4981 & n15756);
  assign n15757 = n4972 | n12253;
  assign n15758 = (n4972 & n4974) | (n4972 & n15757) | (n4974 & n15757);
  assign n4991 = n4965 | n4968;
  assign n4992 = n4958 | n4961;
  assign n12311 = n4916 | n4918;
  assign n15759 = n4815 | n4916;
  assign n15760 = (n4916 & n4918) | (n4916 & n15759) | (n4918 & n15759);
  assign n15761 = (n12238 & n12311) | (n12238 & n15760) | (n12311 & n15760);
  assign n15762 = (n4817 & n12311) | (n4817 & n15760) | (n12311 & n15760);
  assign n15763 = (n12210 & n15761) | (n12210 & n15762) | (n15761 & n15762);
  assign n15764 = n4902 | n4904;
  assign n15765 = (n4902 & n12266) | (n4902 & n15764) | (n12266 & n15764);
  assign n15766 = n4801 | n4902;
  assign n15767 = (n4902 & n4904) | (n4902 & n15766) | (n4904 & n15766);
  assign n15768 = (n15719 & n15765) | (n15719 & n15767) | (n15765 & n15767);
  assign n15769 = (n15721 & n15765) | (n15721 & n15767) | (n15765 & n15767);
  assign n15770 = (n15678 & n15768) | (n15678 & n15769) | (n15768 & n15769);
  assign n5002 = x63 & x80;
  assign n5003 = x62 & x81;
  assign n5004 = n5002 & n5003;
  assign n5005 = n5002 | n5003;
  assign n5006 = ~n5004 & n5005;
  assign n15771 = n4895 | n4897;
  assign n15772 = (n4895 & n12268) | (n4895 & n15771) | (n12268 & n15771);
  assign n12319 = n5006 & n15772;
  assign n15773 = n4794 | n4895;
  assign n15774 = (n4895 & n4897) | (n4895 & n15773) | (n4897 & n15773);
  assign n12320 = n5006 & n15774;
  assign n15775 = (n12319 & n12320) | (n12319 & n15723) | (n12320 & n15723);
  assign n15776 = (n12319 & n12320) | (n12319 & n15724) | (n12320 & n15724);
  assign n15777 = (n15661 & n15775) | (n15661 & n15776) | (n15775 & n15776);
  assign n12322 = n5006 | n15772;
  assign n12323 = n5006 | n15774;
  assign n15778 = (n12322 & n12323) | (n12322 & n15723) | (n12323 & n15723);
  assign n15779 = (n12322 & n12323) | (n12322 & n15724) | (n12323 & n15724);
  assign n15780 = (n15661 & n15778) | (n15661 & n15779) | (n15778 & n15779);
  assign n5009 = ~n15777 & n15780;
  assign n5010 = x61 & x82;
  assign n5011 = n5009 & n5010;
  assign n5012 = n5009 | n5010;
  assign n5013 = ~n5011 & n5012;
  assign n5014 = n15770 & n5013;
  assign n5015 = n15770 | n5013;
  assign n5016 = ~n5014 & n5015;
  assign n5017 = x60 & x83;
  assign n5018 = n5016 & n5017;
  assign n5019 = n5016 | n5017;
  assign n5020 = ~n5018 & n5019;
  assign n12325 = n4909 & n5020;
  assign n15781 = (n5020 & n12282) | (n5020 & n12325) | (n12282 & n12325);
  assign n15782 = (n5020 & n12283) | (n5020 & n12325) | (n12283 & n12325);
  assign n15783 = (n15717 & n15781) | (n15717 & n15782) | (n15781 & n15782);
  assign n12327 = n4909 | n5020;
  assign n15784 = n12282 | n12327;
  assign n15785 = n12283 | n12327;
  assign n15786 = (n15717 & n15784) | (n15717 & n15785) | (n15784 & n15785);
  assign n5023 = ~n15783 & n15786;
  assign n5024 = x59 & x84;
  assign n5025 = n5023 & n5024;
  assign n5026 = n5023 | n5024;
  assign n5027 = ~n5025 & n5026;
  assign n5028 = n15763 & n5027;
  assign n5029 = n15763 | n5027;
  assign n5030 = ~n5028 & n5029;
  assign n5031 = x58 & x85;
  assign n5032 = n5030 & n5031;
  assign n5033 = n5030 | n5031;
  assign n5034 = ~n5032 & n5033;
  assign n12329 = n4923 & n5034;
  assign n12330 = (n5034 & n12293) | (n5034 & n12329) | (n12293 & n12329);
  assign n12331 = n4923 | n5034;
  assign n12332 = n12293 | n12331;
  assign n5037 = ~n12330 & n12332;
  assign n5038 = x57 & x86;
  assign n5039 = n5037 & n5038;
  assign n5040 = n5037 | n5038;
  assign n5041 = ~n5039 & n5040;
  assign n12333 = n4930 & n5041;
  assign n12334 = (n5041 & n12297) | (n5041 & n12333) | (n12297 & n12333);
  assign n12335 = n4930 | n5041;
  assign n12336 = n12297 | n12335;
  assign n5044 = ~n12334 & n12336;
  assign n5045 = x56 & x87;
  assign n5046 = n5044 & n5045;
  assign n5047 = n5044 | n5045;
  assign n5048 = ~n5046 & n5047;
  assign n12337 = n4937 & n5048;
  assign n12338 = (n5048 & n12302) | (n5048 & n12337) | (n12302 & n12337);
  assign n12339 = n4937 | n5048;
  assign n12340 = n12302 | n12339;
  assign n5051 = ~n12338 & n12340;
  assign n5052 = x55 & x88;
  assign n5053 = n5051 & n5052;
  assign n5054 = n5051 | n5052;
  assign n5055 = ~n5053 & n5054;
  assign n12308 = n4944 | n4946;
  assign n12341 = n5055 & n12308;
  assign n12342 = n4944 & n5055;
  assign n12343 = (n12261 & n12341) | (n12261 & n12342) | (n12341 & n12342);
  assign n12344 = n5055 | n12308;
  assign n12345 = n4944 | n5055;
  assign n12346 = (n12261 & n12344) | (n12261 & n12345) | (n12344 & n12345);
  assign n5058 = ~n12343 & n12346;
  assign n5059 = x54 & x89;
  assign n5060 = n5058 & n5059;
  assign n5061 = n5058 | n5059;
  assign n5062 = ~n5060 & n5061;
  assign n12347 = n4951 & n5062;
  assign n12348 = (n4954 & n5062) | (n4954 & n12347) | (n5062 & n12347);
  assign n12349 = n4951 | n5062;
  assign n12350 = n4954 | n12349;
  assign n5065 = ~n12348 & n12350;
  assign n5066 = x53 & x90;
  assign n5067 = n5065 & n5066;
  assign n5068 = n5065 | n5066;
  assign n5069 = ~n5067 & n5068;
  assign n5070 = n4992 & n5069;
  assign n5071 = n4992 | n5069;
  assign n5072 = ~n5070 & n5071;
  assign n5073 = x52 & x91;
  assign n5074 = n5072 & n5073;
  assign n5075 = n5072 | n5073;
  assign n5076 = ~n5074 & n5075;
  assign n5077 = n4991 & n5076;
  assign n5078 = n4991 | n5076;
  assign n5079 = ~n5077 & n5078;
  assign n5080 = x51 & x92;
  assign n5081 = n5079 & n5080;
  assign n5082 = n5079 | n5080;
  assign n5083 = ~n5081 & n5082;
  assign n5084 = n15758 & n5083;
  assign n5085 = n15758 | n5083;
  assign n5086 = ~n5084 & n5085;
  assign n5087 = x50 & x93;
  assign n5088 = n5086 & n5087;
  assign n5089 = n5086 | n5087;
  assign n5090 = ~n5088 & n5089;
  assign n5091 = n12307 & n5090;
  assign n5092 = n12307 | n5090;
  assign n5093 = ~n5091 & n5092;
  assign n5094 = x49 & x94;
  assign n5095 = n5093 & n5094;
  assign n5096 = n5093 | n5094;
  assign n5097 = ~n5095 & n5096;
  assign n5098 = n4986 & n5097;
  assign n5099 = n4986 | n5097;
  assign n5100 = ~n5098 & n5099;
  assign n5101 = x48 & x95;
  assign n5102 = n5100 & n5101;
  assign n5103 = n5100 | n5101;
  assign n5104 = ~n5102 & n5103;
  assign n17692 = n4985 | n5094;
  assign n17693 = (n4984 & n5094) | (n4984 & n17692) | (n5094 & n17692);
  assign n15788 = (n4986 & n5093) | (n4986 & n17693) | (n5093 & n17693);
  assign n12352 = (n5095 & n5097) | (n5095 & n15788) | (n5097 & n15788);
  assign n12353 = n5088 | n12307;
  assign n12354 = (n5088 & n5090) | (n5088 & n12353) | (n5090 & n12353);
  assign n15789 = n5081 | n15758;
  assign n15790 = (n5081 & n5083) | (n5081 & n15789) | (n5083 & n15789);
  assign n5108 = n5074 | n5077;
  assign n12355 = n5067 | n5069;
  assign n12356 = (n4992 & n5067) | (n4992 & n12355) | (n5067 & n12355);
  assign n12360 = n5018 | n5020;
  assign n15791 = n4909 | n5018;
  assign n15792 = (n5018 & n5020) | (n5018 & n15791) | (n5020 & n15791);
  assign n15793 = (n12282 & n12360) | (n12282 & n15792) | (n12360 & n15792);
  assign n15794 = (n12283 & n12360) | (n12283 & n15792) | (n12360 & n15792);
  assign n15795 = (n15717 & n15793) | (n15717 & n15794) | (n15793 & n15794);
  assign n5119 = x64 & x80;
  assign n5120 = x63 & x81;
  assign n5121 = n5119 & n5120;
  assign n5122 = n5119 | n5120;
  assign n5123 = ~n5121 & n5122;
  assign n15796 = n5004 | n5006;
  assign n15801 = (n5004 & n15774) | (n5004 & n15796) | (n15774 & n15796);
  assign n12368 = n5123 & n15801;
  assign n15798 = n5123 & n15796;
  assign n15799 = n5004 & n5123;
  assign n15800 = (n15772 & n15798) | (n15772 & n15799) | (n15798 & n15799);
  assign n15802 = (n12368 & n15723) | (n12368 & n15800) | (n15723 & n15800);
  assign n15803 = (n12368 & n15724) | (n12368 & n15800) | (n15724 & n15800);
  assign n15804 = (n15661 & n15802) | (n15661 & n15803) | (n15802 & n15803);
  assign n12371 = n5123 | n15801;
  assign n15805 = n5123 | n15796;
  assign n15806 = n5004 | n5123;
  assign n15807 = (n15772 & n15805) | (n15772 & n15806) | (n15805 & n15806);
  assign n15808 = (n12371 & n15723) | (n12371 & n15807) | (n15723 & n15807);
  assign n15809 = (n12371 & n15724) | (n12371 & n15807) | (n15724 & n15807);
  assign n15810 = (n15661 & n15808) | (n15661 & n15809) | (n15808 & n15809);
  assign n5126 = ~n15804 & n15810;
  assign n5127 = x62 & x82;
  assign n5128 = n5126 & n5127;
  assign n5129 = n5126 | n5127;
  assign n5130 = ~n5128 & n5129;
  assign n12362 = n5011 | n5013;
  assign n12373 = n5130 & n12362;
  assign n12374 = n5011 & n5130;
  assign n12375 = (n15770 & n12373) | (n15770 & n12374) | (n12373 & n12374);
  assign n12376 = n5130 | n12362;
  assign n12377 = n5011 | n5130;
  assign n12378 = (n15770 & n12376) | (n15770 & n12377) | (n12376 & n12377);
  assign n5133 = ~n12375 & n12378;
  assign n5134 = x61 & x83;
  assign n5135 = n5133 & n5134;
  assign n5136 = n5133 | n5134;
  assign n5137 = ~n5135 & n5136;
  assign n5138 = n15795 & n5137;
  assign n5139 = n15795 | n5137;
  assign n5140 = ~n5138 & n5139;
  assign n5141 = x60 & x84;
  assign n5142 = n5140 & n5141;
  assign n5143 = n5140 | n5141;
  assign n5144 = ~n5142 & n5143;
  assign n12357 = n5025 | n5027;
  assign n12379 = n5144 & n12357;
  assign n12380 = n5025 & n5144;
  assign n12381 = (n15763 & n12379) | (n15763 & n12380) | (n12379 & n12380);
  assign n12382 = n5144 | n12357;
  assign n12383 = n5025 | n5144;
  assign n12384 = (n15763 & n12382) | (n15763 & n12383) | (n12382 & n12383);
  assign n5147 = ~n12381 & n12384;
  assign n5148 = x59 & x85;
  assign n5149 = n5147 & n5148;
  assign n5150 = n5147 | n5148;
  assign n5151 = ~n5149 & n5150;
  assign n12385 = n5032 & n5151;
  assign n15811 = (n5151 & n12329) | (n5151 & n12385) | (n12329 & n12385);
  assign n15812 = (n5034 & n5151) | (n5034 & n12385) | (n5151 & n12385);
  assign n15813 = (n12293 & n15811) | (n12293 & n15812) | (n15811 & n15812);
  assign n12387 = n5032 | n5151;
  assign n15814 = n12329 | n12387;
  assign n15815 = n5034 | n12387;
  assign n15816 = (n12293 & n15814) | (n12293 & n15815) | (n15814 & n15815);
  assign n5154 = ~n15813 & n15816;
  assign n5155 = x58 & x86;
  assign n5156 = n5154 & n5155;
  assign n5157 = n5154 | n5155;
  assign n5158 = ~n5156 & n5157;
  assign n12389 = n5039 & n5158;
  assign n12390 = (n5158 & n12334) | (n5158 & n12389) | (n12334 & n12389);
  assign n12391 = n5039 | n5158;
  assign n12392 = n12334 | n12391;
  assign n5161 = ~n12390 & n12392;
  assign n5162 = x57 & x87;
  assign n5163 = n5161 & n5162;
  assign n5164 = n5161 | n5162;
  assign n5165 = ~n5163 & n5164;
  assign n12393 = n5046 & n5165;
  assign n12394 = (n5165 & n12338) | (n5165 & n12393) | (n12338 & n12393);
  assign n12395 = n5046 | n5165;
  assign n12396 = n12338 | n12395;
  assign n5168 = ~n12394 & n12396;
  assign n5169 = x56 & x88;
  assign n5170 = n5168 & n5169;
  assign n5171 = n5168 | n5169;
  assign n5172 = ~n5170 & n5171;
  assign n12397 = n5053 & n5172;
  assign n12398 = (n5172 & n12343) | (n5172 & n12397) | (n12343 & n12397);
  assign n12399 = n5053 | n5172;
  assign n12400 = n12343 | n12399;
  assign n5175 = ~n12398 & n12400;
  assign n5176 = x55 & x89;
  assign n5177 = n5175 & n5176;
  assign n5178 = n5175 | n5176;
  assign n5179 = ~n5177 & n5178;
  assign n12401 = n5060 & n5179;
  assign n12402 = (n5179 & n12348) | (n5179 & n12401) | (n12348 & n12401);
  assign n12403 = n5060 | n5179;
  assign n12404 = n12348 | n12403;
  assign n5182 = ~n12402 & n12404;
  assign n5183 = x54 & x90;
  assign n5184 = n5182 & n5183;
  assign n5185 = n5182 | n5183;
  assign n5186 = ~n5184 & n5185;
  assign n5187 = n12356 & n5186;
  assign n5188 = n12356 | n5186;
  assign n5189 = ~n5187 & n5188;
  assign n5190 = x53 & x91;
  assign n5191 = n5189 & n5190;
  assign n5192 = n5189 | n5190;
  assign n5193 = ~n5191 & n5192;
  assign n5194 = n5108 & n5193;
  assign n5195 = n5108 | n5193;
  assign n5196 = ~n5194 & n5195;
  assign n5197 = x52 & x92;
  assign n5198 = n5196 & n5197;
  assign n5199 = n5196 | n5197;
  assign n5200 = ~n5198 & n5199;
  assign n5201 = n15790 & n5200;
  assign n5202 = n15790 | n5200;
  assign n5203 = ~n5201 & n5202;
  assign n5204 = x51 & x93;
  assign n5205 = n5203 & n5204;
  assign n5206 = n5203 | n5204;
  assign n5207 = ~n5205 & n5206;
  assign n5208 = n12354 & n5207;
  assign n5209 = n12354 | n5207;
  assign n5210 = ~n5208 & n5209;
  assign n5211 = x50 & x94;
  assign n5212 = n5210 & n5211;
  assign n5213 = n5210 | n5211;
  assign n5214 = ~n5212 & n5213;
  assign n5215 = n12352 & n5214;
  assign n5216 = n12352 | n5214;
  assign n5217 = ~n5215 & n5216;
  assign n5218 = x49 & x95;
  assign n5219 = n5217 & n5218;
  assign n5220 = n5217 | n5218;
  assign n5221 = ~n5219 & n5220;
  assign n5222 = n5102 & n5221;
  assign n5223 = n5102 | n5221;
  assign n5224 = ~n5222 & n5223;
  assign n5225 = x48 & x96;
  assign n5226 = n5224 & n5225;
  assign n5227 = n5224 | n5225;
  assign n5228 = ~n5226 & n5227;
  assign n17694 = n5101 | n5218;
  assign n17695 = (n5100 & n5218) | (n5100 & n17694) | (n5218 & n17694);
  assign n15818 = (n5102 & n5217) | (n5102 & n17695) | (n5217 & n17695);
  assign n12406 = (n5219 & n5221) | (n5219 & n15818) | (n5221 & n15818);
  assign n12407 = n5212 | n12352;
  assign n12408 = (n5212 & n5214) | (n5212 & n12407) | (n5214 & n12407);
  assign n12409 = n5205 | n12354;
  assign n12410 = (n5205 & n5207) | (n5205 & n12409) | (n5207 & n12409);
  assign n15819 = n5198 | n15790;
  assign n15820 = (n5198 & n5200) | (n5198 & n15819) | (n5200 & n15819);
  assign n12411 = n5191 | n5193;
  assign n12412 = (n5108 & n5191) | (n5108 & n12411) | (n5191 & n12411);
  assign n12413 = n5184 | n5186;
  assign n12414 = (n5184 & n12356) | (n5184 & n12413) | (n12356 & n12413);
  assign n12416 = n5149 | n5151;
  assign n15821 = n5032 | n5149;
  assign n15822 = (n5149 & n5151) | (n5149 & n15821) | (n5151 & n15821);
  assign n15823 = (n12329 & n12416) | (n12329 & n15822) | (n12416 & n15822);
  assign n15824 = (n5034 & n12416) | (n5034 & n15822) | (n12416 & n15822);
  assign n15825 = (n12293 & n15823) | (n12293 & n15824) | (n15823 & n15824);
  assign n5244 = x65 & x80;
  assign n5245 = x64 & x81;
  assign n5246 = n5244 & n5245;
  assign n5247 = n5244 | n5245;
  assign n5248 = ~n5246 & n5247;
  assign n12423 = n5121 & n5248;
  assign n12424 = (n5248 & n15804) | (n5248 & n12423) | (n15804 & n12423);
  assign n12425 = n5121 | n5248;
  assign n12426 = n15804 | n12425;
  assign n5251 = ~n12424 & n12426;
  assign n5252 = x63 & x82;
  assign n5253 = n5251 & n5252;
  assign n5254 = n5251 | n5252;
  assign n5255 = ~n5253 & n5254;
  assign n15826 = n5128 | n5130;
  assign n15827 = (n5128 & n12362) | (n5128 & n15826) | (n12362 & n15826);
  assign n12427 = n5255 & n15827;
  assign n15828 = n5011 | n5128;
  assign n15829 = (n5128 & n5130) | (n5128 & n15828) | (n5130 & n15828);
  assign n12428 = n5255 & n15829;
  assign n12429 = (n15770 & n12427) | (n15770 & n12428) | (n12427 & n12428);
  assign n12430 = n5255 | n15827;
  assign n12431 = n5255 | n15829;
  assign n12432 = (n15770 & n12430) | (n15770 & n12431) | (n12430 & n12431);
  assign n5258 = ~n12429 & n12432;
  assign n5259 = x62 & x83;
  assign n5260 = n5258 & n5259;
  assign n5261 = n5258 | n5259;
  assign n5262 = ~n5260 & n5261;
  assign n12418 = n5135 | n5137;
  assign n12433 = n5262 & n12418;
  assign n12434 = n5135 & n5262;
  assign n12435 = (n15795 & n12433) | (n15795 & n12434) | (n12433 & n12434);
  assign n12436 = n5262 | n12418;
  assign n12437 = n5135 | n5262;
  assign n12438 = (n15795 & n12436) | (n15795 & n12437) | (n12436 & n12437);
  assign n5265 = ~n12435 & n12438;
  assign n5266 = x61 & x84;
  assign n5267 = n5265 & n5266;
  assign n5268 = n5265 | n5266;
  assign n5269 = ~n5267 & n5268;
  assign n12439 = n5142 & n5269;
  assign n15830 = (n5269 & n12380) | (n5269 & n12439) | (n12380 & n12439);
  assign n15831 = (n5269 & n12379) | (n5269 & n12439) | (n12379 & n12439);
  assign n15832 = (n15763 & n15830) | (n15763 & n15831) | (n15830 & n15831);
  assign n12441 = n5142 | n5269;
  assign n15833 = n12380 | n12441;
  assign n15834 = n12379 | n12441;
  assign n15835 = (n15763 & n15833) | (n15763 & n15834) | (n15833 & n15834);
  assign n5272 = ~n15832 & n15835;
  assign n5273 = x60 & x85;
  assign n5274 = n5272 & n5273;
  assign n5275 = n5272 | n5273;
  assign n5276 = ~n5274 & n5275;
  assign n5277 = n15825 & n5276;
  assign n5278 = n15825 | n5276;
  assign n5279 = ~n5277 & n5278;
  assign n5280 = x59 & x86;
  assign n5281 = n5279 & n5280;
  assign n5282 = n5279 | n5280;
  assign n5283 = ~n5281 & n5282;
  assign n12443 = n5156 & n5283;
  assign n12444 = (n5283 & n12390) | (n5283 & n12443) | (n12390 & n12443);
  assign n12445 = n5156 | n5283;
  assign n12446 = n12390 | n12445;
  assign n5286 = ~n12444 & n12446;
  assign n5287 = x58 & x87;
  assign n5288 = n5286 & n5287;
  assign n5289 = n5286 | n5287;
  assign n5290 = ~n5288 & n5289;
  assign n12447 = n5163 & n5290;
  assign n12448 = (n5290 & n12394) | (n5290 & n12447) | (n12394 & n12447);
  assign n12449 = n5163 | n5290;
  assign n12450 = n12394 | n12449;
  assign n5293 = ~n12448 & n12450;
  assign n5294 = x57 & x88;
  assign n5295 = n5293 & n5294;
  assign n5296 = n5293 | n5294;
  assign n5297 = ~n5295 & n5296;
  assign n12451 = n5170 & n5297;
  assign n12452 = (n5297 & n12398) | (n5297 & n12451) | (n12398 & n12451);
  assign n12453 = n5170 | n5297;
  assign n12454 = n12398 | n12453;
  assign n5300 = ~n12452 & n12454;
  assign n5301 = x56 & x89;
  assign n5302 = n5300 & n5301;
  assign n5303 = n5300 | n5301;
  assign n5304 = ~n5302 & n5303;
  assign n12455 = n5177 & n5304;
  assign n12456 = (n5304 & n12402) | (n5304 & n12455) | (n12402 & n12455);
  assign n12457 = n5177 | n5304;
  assign n12458 = n12402 | n12457;
  assign n5307 = ~n12456 & n12458;
  assign n5308 = x55 & x90;
  assign n5309 = n5307 & n5308;
  assign n5310 = n5307 | n5308;
  assign n5311 = ~n5309 & n5310;
  assign n5312 = n12414 & n5311;
  assign n5313 = n12414 | n5311;
  assign n5314 = ~n5312 & n5313;
  assign n5315 = x54 & x91;
  assign n5316 = n5314 & n5315;
  assign n5317 = n5314 | n5315;
  assign n5318 = ~n5316 & n5317;
  assign n5319 = n12412 & n5318;
  assign n5320 = n12412 | n5318;
  assign n5321 = ~n5319 & n5320;
  assign n5322 = x53 & x92;
  assign n5323 = n5321 & n5322;
  assign n5324 = n5321 | n5322;
  assign n5325 = ~n5323 & n5324;
  assign n5326 = n15820 & n5325;
  assign n5327 = n15820 | n5325;
  assign n5328 = ~n5326 & n5327;
  assign n5329 = x52 & x93;
  assign n5330 = n5328 & n5329;
  assign n5331 = n5328 | n5329;
  assign n5332 = ~n5330 & n5331;
  assign n5333 = n12410 & n5332;
  assign n5334 = n12410 | n5332;
  assign n5335 = ~n5333 & n5334;
  assign n5336 = x51 & x94;
  assign n5337 = n5335 & n5336;
  assign n5338 = n5335 | n5336;
  assign n5339 = ~n5337 & n5338;
  assign n5340 = n12408 & n5339;
  assign n5341 = n12408 | n5339;
  assign n5342 = ~n5340 & n5341;
  assign n5343 = x50 & x95;
  assign n5344 = n5342 & n5343;
  assign n5345 = n5342 | n5343;
  assign n5346 = ~n5344 & n5345;
  assign n5347 = n12406 & n5346;
  assign n5348 = n12406 | n5346;
  assign n5349 = ~n5347 & n5348;
  assign n5350 = x49 & x96;
  assign n5351 = n5349 & n5350;
  assign n5352 = n5349 | n5350;
  assign n5353 = ~n5351 & n5352;
  assign n5354 = n5226 & n5353;
  assign n5355 = n5226 | n5353;
  assign n5356 = ~n5354 & n5355;
  assign n5357 = x48 & x97;
  assign n5358 = n5356 & n5357;
  assign n5359 = n5356 | n5357;
  assign n5360 = ~n5358 & n5359;
  assign n12459 = n5226 | n5351;
  assign n12460 = (n5351 & n5353) | (n5351 & n12459) | (n5353 & n12459);
  assign n12461 = n5344 | n12406;
  assign n12462 = (n5344 & n5346) | (n5344 & n12461) | (n5346 & n12461);
  assign n12463 = n5337 | n12408;
  assign n12464 = (n5337 & n5339) | (n5337 & n12463) | (n5339 & n12463);
  assign n12465 = n5330 | n12410;
  assign n12466 = (n5330 & n5332) | (n5330 & n12465) | (n5332 & n12465);
  assign n12467 = n5323 | n5325;
  assign n12468 = (n15820 & n5323) | (n15820 & n12467) | (n5323 & n12467);
  assign n12469 = n5316 | n5318;
  assign n12470 = (n5316 & n12412) | (n5316 & n12469) | (n12412 & n12469);
  assign n12471 = n5309 | n5311;
  assign n12472 = (n5309 & n12414) | (n5309 & n12471) | (n12414 & n12471);
  assign n12476 = n5267 | n5269;
  assign n15836 = n5142 | n5267;
  assign n15837 = (n5267 & n5269) | (n5267 & n15836) | (n5269 & n15836);
  assign n15838 = (n12380 & n12476) | (n12380 & n15837) | (n12476 & n15837);
  assign n15839 = (n12379 & n12476) | (n12379 & n15837) | (n12476 & n15837);
  assign n15840 = (n15763 & n15838) | (n15763 & n15839) | (n15838 & n15839);
  assign n5377 = x66 & x80;
  assign n5378 = x65 & x81;
  assign n5379 = n5377 & n5378;
  assign n5380 = n5377 | n5378;
  assign n5381 = ~n5379 & n5380;
  assign n15845 = n5121 | n5246;
  assign n15846 = (n5246 & n5248) | (n5246 & n15845) | (n5248 & n15845);
  assign n12484 = n5381 & n15846;
  assign n12482 = n5246 | n5248;
  assign n12485 = n5381 & n12482;
  assign n12486 = (n15804 & n12484) | (n15804 & n12485) | (n12484 & n12485);
  assign n12487 = n5381 | n15846;
  assign n12488 = n5381 | n12482;
  assign n12489 = (n15804 & n12487) | (n15804 & n12488) | (n12487 & n12488);
  assign n5384 = ~n12486 & n12489;
  assign n5385 = x64 & x82;
  assign n5386 = n5384 & n5385;
  assign n5387 = n5384 | n5385;
  assign n5388 = ~n5386 & n5387;
  assign n12490 = n5253 & n5388;
  assign n15847 = (n5388 & n12427) | (n5388 & n12490) | (n12427 & n12490);
  assign n15848 = (n5388 & n12428) | (n5388 & n12490) | (n12428 & n12490);
  assign n15849 = (n15770 & n15847) | (n15770 & n15848) | (n15847 & n15848);
  assign n12492 = n5253 | n5388;
  assign n15850 = n12427 | n12492;
  assign n15851 = n12428 | n12492;
  assign n15852 = (n15770 & n15850) | (n15770 & n15851) | (n15850 & n15851);
  assign n5391 = ~n15849 & n15852;
  assign n5392 = x63 & x83;
  assign n5393 = n5391 & n5392;
  assign n5394 = n5391 | n5392;
  assign n5395 = ~n5393 & n5394;
  assign n15841 = n5260 | n5262;
  assign n15842 = (n5260 & n12418) | (n5260 & n15841) | (n12418 & n15841);
  assign n15853 = n5395 & n15842;
  assign n15843 = n5135 | n5260;
  assign n15844 = (n5260 & n5262) | (n5260 & n15843) | (n5262 & n15843);
  assign n15854 = n5395 & n15844;
  assign n15855 = (n15795 & n15853) | (n15795 & n15854) | (n15853 & n15854);
  assign n15856 = n5395 | n15842;
  assign n15857 = n5395 | n15844;
  assign n15858 = (n15795 & n15856) | (n15795 & n15857) | (n15856 & n15857);
  assign n5398 = ~n15855 & n15858;
  assign n5399 = x62 & x84;
  assign n5400 = n5398 & n5399;
  assign n5401 = n5398 | n5399;
  assign n5402 = ~n5400 & n5401;
  assign n5403 = n15840 & n5402;
  assign n5404 = n15840 | n5402;
  assign n5405 = ~n5403 & n5404;
  assign n5406 = x61 & x85;
  assign n5407 = n5405 & n5406;
  assign n5408 = n5405 | n5406;
  assign n5409 = ~n5407 & n5408;
  assign n12473 = n5274 | n5276;
  assign n12494 = n5409 & n12473;
  assign n12495 = n5274 & n5409;
  assign n12496 = (n15825 & n12494) | (n15825 & n12495) | (n12494 & n12495);
  assign n12497 = n5409 | n12473;
  assign n12498 = n5274 | n5409;
  assign n12499 = (n15825 & n12497) | (n15825 & n12498) | (n12497 & n12498);
  assign n5412 = ~n12496 & n12499;
  assign n5413 = x60 & x86;
  assign n5414 = n5412 & n5413;
  assign n5415 = n5412 | n5413;
  assign n5416 = ~n5414 & n5415;
  assign n12500 = n5281 & n5416;
  assign n15859 = (n5416 & n12443) | (n5416 & n12500) | (n12443 & n12500);
  assign n15860 = (n5283 & n5416) | (n5283 & n12500) | (n5416 & n12500);
  assign n15861 = (n12390 & n15859) | (n12390 & n15860) | (n15859 & n15860);
  assign n12502 = n5281 | n5416;
  assign n15862 = n12443 | n12502;
  assign n15863 = n5283 | n12502;
  assign n15864 = (n12390 & n15862) | (n12390 & n15863) | (n15862 & n15863);
  assign n5419 = ~n15861 & n15864;
  assign n5420 = x59 & x87;
  assign n5421 = n5419 & n5420;
  assign n5422 = n5419 | n5420;
  assign n5423 = ~n5421 & n5422;
  assign n12504 = n5288 & n5423;
  assign n12505 = (n5423 & n12448) | (n5423 & n12504) | (n12448 & n12504);
  assign n12506 = n5288 | n5423;
  assign n12507 = n12448 | n12506;
  assign n5426 = ~n12505 & n12507;
  assign n5427 = x58 & x88;
  assign n5428 = n5426 & n5427;
  assign n5429 = n5426 | n5427;
  assign n5430 = ~n5428 & n5429;
  assign n12508 = n5295 & n5430;
  assign n12509 = (n5430 & n12452) | (n5430 & n12508) | (n12452 & n12508);
  assign n12510 = n5295 | n5430;
  assign n12511 = n12452 | n12510;
  assign n5433 = ~n12509 & n12511;
  assign n5434 = x57 & x89;
  assign n5435 = n5433 & n5434;
  assign n5436 = n5433 | n5434;
  assign n5437 = ~n5435 & n5436;
  assign n12512 = n5302 & n5437;
  assign n12513 = (n5437 & n12456) | (n5437 & n12512) | (n12456 & n12512);
  assign n12514 = n5302 | n5437;
  assign n12515 = n12456 | n12514;
  assign n5440 = ~n12513 & n12515;
  assign n5441 = x56 & x90;
  assign n5442 = n5440 & n5441;
  assign n5443 = n5440 | n5441;
  assign n5444 = ~n5442 & n5443;
  assign n5445 = n12472 & n5444;
  assign n5446 = n12472 | n5444;
  assign n5447 = ~n5445 & n5446;
  assign n5448 = x55 & x91;
  assign n5449 = n5447 & n5448;
  assign n5450 = n5447 | n5448;
  assign n5451 = ~n5449 & n5450;
  assign n5452 = n12470 & n5451;
  assign n5453 = n12470 | n5451;
  assign n5454 = ~n5452 & n5453;
  assign n5455 = x54 & x92;
  assign n5456 = n5454 & n5455;
  assign n5457 = n5454 | n5455;
  assign n5458 = ~n5456 & n5457;
  assign n5459 = n12468 & n5458;
  assign n5460 = n12468 | n5458;
  assign n5461 = ~n5459 & n5460;
  assign n5462 = x53 & x93;
  assign n5463 = n5461 & n5462;
  assign n5464 = n5461 | n5462;
  assign n5465 = ~n5463 & n5464;
  assign n5466 = n12466 & n5465;
  assign n5467 = n12466 | n5465;
  assign n5468 = ~n5466 & n5467;
  assign n5469 = x52 & x94;
  assign n5470 = n5468 & n5469;
  assign n5471 = n5468 | n5469;
  assign n5472 = ~n5470 & n5471;
  assign n5473 = n12464 & n5472;
  assign n5474 = n12464 | n5472;
  assign n5475 = ~n5473 & n5474;
  assign n5476 = x51 & x95;
  assign n5477 = n5475 & n5476;
  assign n5478 = n5475 | n5476;
  assign n5479 = ~n5477 & n5478;
  assign n5480 = n12462 & n5479;
  assign n5481 = n12462 | n5479;
  assign n5482 = ~n5480 & n5481;
  assign n5483 = x50 & x96;
  assign n5484 = n5482 & n5483;
  assign n5485 = n5482 | n5483;
  assign n5486 = ~n5484 & n5485;
  assign n5487 = n12460 & n5486;
  assign n5488 = n12460 | n5486;
  assign n5489 = ~n5487 & n5488;
  assign n5490 = x49 & x97;
  assign n5491 = n5489 & n5490;
  assign n5492 = n5489 | n5490;
  assign n5493 = ~n5491 & n5492;
  assign n5494 = n5358 & n5493;
  assign n5495 = n5358 | n5493;
  assign n5496 = ~n5494 & n5495;
  assign n5497 = x48 & x98;
  assign n5498 = n5496 & n5497;
  assign n5499 = n5496 | n5497;
  assign n5500 = ~n5498 & n5499;
  assign n17696 = n5357 | n5490;
  assign n17697 = (n5356 & n5490) | (n5356 & n17696) | (n5490 & n17696);
  assign n15866 = (n5358 & n5489) | (n5358 & n17697) | (n5489 & n17697);
  assign n12517 = (n5491 & n5493) | (n5491 & n15866) | (n5493 & n15866);
  assign n15867 = n5484 | n12460;
  assign n15868 = (n5484 & n5486) | (n5484 & n15867) | (n5486 & n15867);
  assign n5503 = n5477 | n5480;
  assign n5504 = n5470 | n5473;
  assign n5505 = n5463 | n5466;
  assign n12518 = n5456 | n5458;
  assign n12519 = (n5456 & n12468) | (n5456 & n12518) | (n12468 & n12518);
  assign n12520 = n5449 | n5451;
  assign n12521 = (n5449 & n12470) | (n5449 & n12520) | (n12470 & n12520);
  assign n12522 = n5442 | n5444;
  assign n12523 = (n5442 & n12472) | (n5442 & n12522) | (n12472 & n12522);
  assign n12525 = n5414 | n5416;
  assign n15869 = n5281 | n5414;
  assign n15870 = (n5414 & n5416) | (n5414 & n15869) | (n5416 & n15869);
  assign n15871 = (n12443 & n12525) | (n12443 & n15870) | (n12525 & n15870);
  assign n15872 = (n5283 & n12525) | (n5283 & n15870) | (n12525 & n15870);
  assign n15873 = (n12390 & n15871) | (n12390 & n15872) | (n15871 & n15872);
  assign n5518 = x67 & x80;
  assign n5519 = x66 & x81;
  assign n5520 = n5518 & n5519;
  assign n5521 = n5518 | n5519;
  assign n5522 = ~n5520 & n5521;
  assign n15874 = n5379 | n5381;
  assign n15875 = (n5379 & n15846) | (n5379 & n15874) | (n15846 & n15874);
  assign n12537 = n5522 & n15875;
  assign n15876 = (n5379 & n12482) | (n5379 & n15874) | (n12482 & n15874);
  assign n12538 = n5522 & n15876;
  assign n12539 = (n15804 & n12537) | (n15804 & n12538) | (n12537 & n12538);
  assign n12540 = n5522 | n15875;
  assign n12541 = n5522 | n15876;
  assign n12542 = (n15804 & n12540) | (n15804 & n12541) | (n12540 & n12541);
  assign n5525 = ~n12539 & n12542;
  assign n5526 = x65 & x82;
  assign n5527 = n5525 & n5526;
  assign n5528 = n5525 | n5526;
  assign n5529 = ~n5527 & n5528;
  assign n15877 = n5253 | n5386;
  assign n15878 = (n5386 & n5388) | (n5386 & n15877) | (n5388 & n15877);
  assign n12543 = n5529 & n15878;
  assign n12532 = n5386 | n5388;
  assign n12544 = n5529 & n12532;
  assign n15879 = (n12427 & n12543) | (n12427 & n12544) | (n12543 & n12544);
  assign n15880 = (n12428 & n12543) | (n12428 & n12544) | (n12543 & n12544);
  assign n15881 = (n15770 & n15879) | (n15770 & n15880) | (n15879 & n15880);
  assign n12546 = n5529 | n15878;
  assign n12547 = n5529 | n12532;
  assign n15882 = (n12427 & n12546) | (n12427 & n12547) | (n12546 & n12547);
  assign n15883 = (n12428 & n12546) | (n12428 & n12547) | (n12546 & n12547);
  assign n15884 = (n15770 & n15882) | (n15770 & n15883) | (n15882 & n15883);
  assign n5532 = ~n15881 & n15884;
  assign n5533 = x64 & x83;
  assign n5534 = n5532 & n5533;
  assign n5535 = n5532 | n5533;
  assign n5536 = ~n5534 & n5535;
  assign n12529 = n5393 | n5395;
  assign n12549 = n5536 & n12529;
  assign n12550 = n5393 & n5536;
  assign n15885 = (n12549 & n12550) | (n12549 & n15842) | (n12550 & n15842);
  assign n15886 = (n12549 & n12550) | (n12549 & n15844) | (n12550 & n15844);
  assign n15887 = (n15795 & n15885) | (n15795 & n15886) | (n15885 & n15886);
  assign n12552 = n5536 | n12529;
  assign n12553 = n5393 | n5536;
  assign n15888 = (n12552 & n12553) | (n12552 & n15842) | (n12553 & n15842);
  assign n15889 = (n12552 & n12553) | (n12552 & n15844) | (n12553 & n15844);
  assign n15890 = (n15795 & n15888) | (n15795 & n15889) | (n15888 & n15889);
  assign n5539 = ~n15887 & n15890;
  assign n5540 = x63 & x84;
  assign n5541 = n5539 & n5540;
  assign n5542 = n5539 | n5540;
  assign n5543 = ~n5541 & n5542;
  assign n12527 = n5400 | n5402;
  assign n12555 = n5543 & n12527;
  assign n12556 = n5400 & n5543;
  assign n12557 = (n15840 & n12555) | (n15840 & n12556) | (n12555 & n12556);
  assign n12558 = n5543 | n12527;
  assign n12559 = n5400 | n5543;
  assign n12560 = (n15840 & n12558) | (n15840 & n12559) | (n12558 & n12559);
  assign n5546 = ~n12557 & n12560;
  assign n5547 = x62 & x85;
  assign n5548 = n5546 & n5547;
  assign n5549 = n5546 | n5547;
  assign n5550 = ~n5548 & n5549;
  assign n12561 = n5407 & n5550;
  assign n15891 = (n5550 & n12495) | (n5550 & n12561) | (n12495 & n12561);
  assign n15892 = (n5550 & n12494) | (n5550 & n12561) | (n12494 & n12561);
  assign n15893 = (n15825 & n15891) | (n15825 & n15892) | (n15891 & n15892);
  assign n12563 = n5407 | n5550;
  assign n15894 = n12495 | n12563;
  assign n15895 = n12494 | n12563;
  assign n15896 = (n15825 & n15894) | (n15825 & n15895) | (n15894 & n15895);
  assign n5553 = ~n15893 & n15896;
  assign n5554 = x61 & x86;
  assign n5555 = n5553 & n5554;
  assign n5556 = n5553 | n5554;
  assign n5557 = ~n5555 & n5556;
  assign n5558 = n15873 & n5557;
  assign n5559 = n15873 | n5557;
  assign n5560 = ~n5558 & n5559;
  assign n5561 = x60 & x87;
  assign n5562 = n5560 & n5561;
  assign n5563 = n5560 | n5561;
  assign n5564 = ~n5562 & n5563;
  assign n12565 = n5421 & n5564;
  assign n12566 = (n5564 & n12505) | (n5564 & n12565) | (n12505 & n12565);
  assign n12567 = n5421 | n5564;
  assign n12568 = n12505 | n12567;
  assign n5567 = ~n12566 & n12568;
  assign n5568 = x59 & x88;
  assign n5569 = n5567 & n5568;
  assign n5570 = n5567 | n5568;
  assign n5571 = ~n5569 & n5570;
  assign n12569 = n5428 & n5571;
  assign n12570 = (n5571 & n12509) | (n5571 & n12569) | (n12509 & n12569);
  assign n12571 = n5428 | n5571;
  assign n12572 = n12509 | n12571;
  assign n5574 = ~n12570 & n12572;
  assign n5575 = x58 & x89;
  assign n5576 = n5574 & n5575;
  assign n5577 = n5574 | n5575;
  assign n5578 = ~n5576 & n5577;
  assign n12573 = n5435 & n5578;
  assign n12574 = (n5578 & n12513) | (n5578 & n12573) | (n12513 & n12573);
  assign n12575 = n5435 | n5578;
  assign n12576 = n12513 | n12575;
  assign n5581 = ~n12574 & n12576;
  assign n5582 = x57 & x90;
  assign n5583 = n5581 & n5582;
  assign n5584 = n5581 | n5582;
  assign n5585 = ~n5583 & n5584;
  assign n5586 = n12523 & n5585;
  assign n5587 = n12523 | n5585;
  assign n5588 = ~n5586 & n5587;
  assign n5589 = x56 & x91;
  assign n5590 = n5588 & n5589;
  assign n5591 = n5588 | n5589;
  assign n5592 = ~n5590 & n5591;
  assign n5593 = n12521 & n5592;
  assign n5594 = n12521 | n5592;
  assign n5595 = ~n5593 & n5594;
  assign n5596 = x55 & x92;
  assign n5597 = n5595 & n5596;
  assign n5598 = n5595 | n5596;
  assign n5599 = ~n5597 & n5598;
  assign n5600 = n12519 & n5599;
  assign n5601 = n12519 | n5599;
  assign n5602 = ~n5600 & n5601;
  assign n5603 = x54 & x93;
  assign n5604 = n5602 & n5603;
  assign n5605 = n5602 | n5603;
  assign n5606 = ~n5604 & n5605;
  assign n5607 = n5505 & n5606;
  assign n5608 = n5505 | n5606;
  assign n5609 = ~n5607 & n5608;
  assign n5610 = x53 & x94;
  assign n5611 = n5609 & n5610;
  assign n5612 = n5609 | n5610;
  assign n5613 = ~n5611 & n5612;
  assign n5614 = n5504 & n5613;
  assign n5615 = n5504 | n5613;
  assign n5616 = ~n5614 & n5615;
  assign n5617 = x52 & x95;
  assign n5618 = n5616 & n5617;
  assign n5619 = n5616 | n5617;
  assign n5620 = ~n5618 & n5619;
  assign n5621 = n5503 & n5620;
  assign n5622 = n5503 | n5620;
  assign n5623 = ~n5621 & n5622;
  assign n5624 = x51 & x96;
  assign n5625 = n5623 & n5624;
  assign n5626 = n5623 | n5624;
  assign n5627 = ~n5625 & n5626;
  assign n5628 = n15868 & n5627;
  assign n5629 = n15868 | n5627;
  assign n5630 = ~n5628 & n5629;
  assign n5631 = x50 & x97;
  assign n5632 = n5630 & n5631;
  assign n5633 = n5630 | n5631;
  assign n5634 = ~n5632 & n5633;
  assign n5635 = n12517 & n5634;
  assign n5636 = n12517 | n5634;
  assign n5637 = ~n5635 & n5636;
  assign n5638 = x49 & x98;
  assign n5639 = n5637 & n5638;
  assign n5640 = n5637 | n5638;
  assign n5641 = ~n5639 & n5640;
  assign n5642 = n5498 & n5641;
  assign n5643 = n5498 | n5641;
  assign n5644 = ~n5642 & n5643;
  assign n5645 = x48 & x99;
  assign n5646 = n5644 & n5645;
  assign n5647 = n5644 | n5645;
  assign n5648 = ~n5646 & n5647;
  assign n17698 = n5497 | n5638;
  assign n17699 = (n5496 & n5638) | (n5496 & n17698) | (n5638 & n17698);
  assign n15898 = (n5498 & n5637) | (n5498 & n17699) | (n5637 & n17699);
  assign n12578 = (n5639 & n5641) | (n5639 & n15898) | (n5641 & n15898);
  assign n12579 = n5632 | n12517;
  assign n12580 = (n5632 & n5634) | (n5632 & n12579) | (n5634 & n12579);
  assign n15899 = n5625 | n15868;
  assign n15900 = (n5625 & n5627) | (n5625 & n15899) | (n5627 & n15899);
  assign n5652 = n5618 | n5621;
  assign n5653 = n5611 | n5614;
  assign n12581 = n5604 | n5606;
  assign n12582 = (n5505 & n5604) | (n5505 & n12581) | (n5604 & n12581);
  assign n12583 = n5597 | n5599;
  assign n12584 = (n5597 & n12519) | (n5597 & n12583) | (n12519 & n12583);
  assign n12585 = n5590 | n5592;
  assign n12586 = (n5590 & n12521) | (n5590 & n12585) | (n12521 & n12585);
  assign n12587 = n5583 | n5585;
  assign n12588 = (n5583 & n12523) | (n5583 & n12587) | (n12523 & n12587);
  assign n12592 = n5548 | n5550;
  assign n15901 = n5407 | n5548;
  assign n15902 = (n5548 & n5550) | (n5548 & n15901) | (n5550 & n15901);
  assign n15903 = (n12495 & n12592) | (n12495 & n15902) | (n12592 & n15902);
  assign n15904 = (n12494 & n12592) | (n12494 & n15902) | (n12592 & n15902);
  assign n15905 = (n15825 & n15903) | (n15825 & n15904) | (n15903 & n15904);
  assign n15906 = n5534 | n5536;
  assign n15907 = (n5534 & n12529) | (n5534 & n15906) | (n12529 & n15906);
  assign n15908 = n5393 | n5534;
  assign n15909 = (n5534 & n5536) | (n5534 & n15908) | (n5536 & n15908);
  assign n15910 = (n15842 & n15907) | (n15842 & n15909) | (n15907 & n15909);
  assign n15911 = (n15844 & n15907) | (n15844 & n15909) | (n15907 & n15909);
  assign n15912 = (n15795 & n15910) | (n15795 & n15911) | (n15910 & n15911);
  assign n15913 = n5527 | n5529;
  assign n15914 = (n5527 & n15878) | (n5527 & n15913) | (n15878 & n15913);
  assign n15915 = (n5527 & n12532) | (n5527 & n15913) | (n12532 & n15913);
  assign n15916 = (n12427 & n15914) | (n12427 & n15915) | (n15914 & n15915);
  assign n15917 = (n12428 & n15914) | (n12428 & n15915) | (n15914 & n15915);
  assign n15918 = (n15770 & n15916) | (n15770 & n15917) | (n15916 & n15917);
  assign n5667 = x68 & x80;
  assign n5668 = x67 & x81;
  assign n5669 = n5667 & n5668;
  assign n5670 = n5667 | n5668;
  assign n5671 = ~n5669 & n5670;
  assign n15919 = n5520 | n5522;
  assign n15921 = n5671 & n15919;
  assign n15922 = n5520 & n5671;
  assign n15923 = (n15875 & n15921) | (n15875 & n15922) | (n15921 & n15922);
  assign n15925 = (n15876 & n15921) | (n15876 & n15922) | (n15921 & n15922);
  assign n12605 = (n15804 & n15923) | (n15804 & n15925) | (n15923 & n15925);
  assign n15926 = n5671 | n15919;
  assign n15927 = n5520 | n5671;
  assign n15928 = (n15875 & n15926) | (n15875 & n15927) | (n15926 & n15927);
  assign n15929 = (n15876 & n15926) | (n15876 & n15927) | (n15926 & n15927);
  assign n12608 = (n15804 & n15928) | (n15804 & n15929) | (n15928 & n15929);
  assign n5674 = ~n12605 & n12608;
  assign n5675 = x66 & x82;
  assign n5676 = n5674 & n5675;
  assign n5677 = n5674 | n5675;
  assign n5678 = ~n5676 & n5677;
  assign n5679 = n15918 & n5678;
  assign n5680 = n15918 | n5678;
  assign n5681 = ~n5679 & n5680;
  assign n5682 = x65 & x83;
  assign n5683 = n5681 & n5682;
  assign n5684 = n5681 | n5682;
  assign n5685 = ~n5683 & n5684;
  assign n5686 = n15912 & n5685;
  assign n5687 = n15912 | n5685;
  assign n5688 = ~n5686 & n5687;
  assign n5689 = x64 & x84;
  assign n5690 = n5688 & n5689;
  assign n5691 = n5688 | n5689;
  assign n5692 = ~n5690 & n5691;
  assign n12609 = n5541 & n5692;
  assign n15930 = (n5692 & n12555) | (n5692 & n12609) | (n12555 & n12609);
  assign n15931 = (n5692 & n12556) | (n5692 & n12609) | (n12556 & n12609);
  assign n15932 = (n15840 & n15930) | (n15840 & n15931) | (n15930 & n15931);
  assign n12611 = n5541 | n5692;
  assign n15933 = n12555 | n12611;
  assign n15934 = n12556 | n12611;
  assign n15935 = (n15840 & n15933) | (n15840 & n15934) | (n15933 & n15934);
  assign n5695 = ~n15932 & n15935;
  assign n5696 = x63 & x85;
  assign n5697 = n5695 & n5696;
  assign n5698 = n5695 | n5696;
  assign n5699 = ~n5697 & n5698;
  assign n5700 = n15905 & n5699;
  assign n5701 = n15905 | n5699;
  assign n5702 = ~n5700 & n5701;
  assign n5703 = x62 & x86;
  assign n5704 = n5702 & n5703;
  assign n5705 = n5702 | n5703;
  assign n5706 = ~n5704 & n5705;
  assign n12589 = n5555 | n5557;
  assign n12613 = n5706 & n12589;
  assign n12614 = n5555 & n5706;
  assign n12615 = (n15873 & n12613) | (n15873 & n12614) | (n12613 & n12614);
  assign n12616 = n5706 | n12589;
  assign n12617 = n5555 | n5706;
  assign n12618 = (n15873 & n12616) | (n15873 & n12617) | (n12616 & n12617);
  assign n5709 = ~n12615 & n12618;
  assign n5710 = x61 & x87;
  assign n5711 = n5709 & n5710;
  assign n5712 = n5709 | n5710;
  assign n5713 = ~n5711 & n5712;
  assign n12619 = n5562 & n5713;
  assign n15936 = (n5713 & n12565) | (n5713 & n12619) | (n12565 & n12619);
  assign n15937 = (n5564 & n5713) | (n5564 & n12619) | (n5713 & n12619);
  assign n15938 = (n12505 & n15936) | (n12505 & n15937) | (n15936 & n15937);
  assign n12621 = n5562 | n5713;
  assign n15939 = n12565 | n12621;
  assign n15940 = n5564 | n12621;
  assign n15941 = (n12505 & n15939) | (n12505 & n15940) | (n15939 & n15940);
  assign n5716 = ~n15938 & n15941;
  assign n5717 = x60 & x88;
  assign n5718 = n5716 & n5717;
  assign n5719 = n5716 | n5717;
  assign n5720 = ~n5718 & n5719;
  assign n12623 = n5569 & n5720;
  assign n12624 = (n5720 & n12570) | (n5720 & n12623) | (n12570 & n12623);
  assign n12625 = n5569 | n5720;
  assign n12626 = n12570 | n12625;
  assign n5723 = ~n12624 & n12626;
  assign n5724 = x59 & x89;
  assign n5725 = n5723 & n5724;
  assign n5726 = n5723 | n5724;
  assign n5727 = ~n5725 & n5726;
  assign n12627 = n5576 & n5727;
  assign n12628 = (n5727 & n12574) | (n5727 & n12627) | (n12574 & n12627);
  assign n12629 = n5576 | n5727;
  assign n12630 = n12574 | n12629;
  assign n5730 = ~n12628 & n12630;
  assign n5731 = x58 & x90;
  assign n5732 = n5730 & n5731;
  assign n5733 = n5730 | n5731;
  assign n5734 = ~n5732 & n5733;
  assign n5735 = n12588 & n5734;
  assign n5736 = n12588 | n5734;
  assign n5737 = ~n5735 & n5736;
  assign n5738 = x57 & x91;
  assign n5739 = n5737 & n5738;
  assign n5740 = n5737 | n5738;
  assign n5741 = ~n5739 & n5740;
  assign n5742 = n12586 & n5741;
  assign n5743 = n12586 | n5741;
  assign n5744 = ~n5742 & n5743;
  assign n5745 = x56 & x92;
  assign n5746 = n5744 & n5745;
  assign n5747 = n5744 | n5745;
  assign n5748 = ~n5746 & n5747;
  assign n5749 = n12584 & n5748;
  assign n5750 = n12584 | n5748;
  assign n5751 = ~n5749 & n5750;
  assign n5752 = x55 & x93;
  assign n5753 = n5751 & n5752;
  assign n5754 = n5751 | n5752;
  assign n5755 = ~n5753 & n5754;
  assign n5756 = n12582 & n5755;
  assign n5757 = n12582 | n5755;
  assign n5758 = ~n5756 & n5757;
  assign n5759 = x54 & x94;
  assign n5760 = n5758 & n5759;
  assign n5761 = n5758 | n5759;
  assign n5762 = ~n5760 & n5761;
  assign n5763 = n5653 & n5762;
  assign n5764 = n5653 | n5762;
  assign n5765 = ~n5763 & n5764;
  assign n5766 = x53 & x95;
  assign n5767 = n5765 & n5766;
  assign n5768 = n5765 | n5766;
  assign n5769 = ~n5767 & n5768;
  assign n5770 = n5652 & n5769;
  assign n5771 = n5652 | n5769;
  assign n5772 = ~n5770 & n5771;
  assign n5773 = x52 & x96;
  assign n5774 = n5772 & n5773;
  assign n5775 = n5772 | n5773;
  assign n5776 = ~n5774 & n5775;
  assign n5777 = n15900 & n5776;
  assign n5778 = n15900 | n5776;
  assign n5779 = ~n5777 & n5778;
  assign n5780 = x51 & x97;
  assign n5781 = n5779 & n5780;
  assign n5782 = n5779 | n5780;
  assign n5783 = ~n5781 & n5782;
  assign n5784 = n12580 & n5783;
  assign n5785 = n12580 | n5783;
  assign n5786 = ~n5784 & n5785;
  assign n5787 = x50 & x98;
  assign n5788 = n5786 & n5787;
  assign n5789 = n5786 | n5787;
  assign n5790 = ~n5788 & n5789;
  assign n5791 = n12578 & n5790;
  assign n5792 = n12578 | n5790;
  assign n5793 = ~n5791 & n5792;
  assign n5794 = x49 & x99;
  assign n5795 = n5793 & n5794;
  assign n5796 = n5793 | n5794;
  assign n5797 = ~n5795 & n5796;
  assign n5798 = n5646 & n5797;
  assign n5799 = n5646 | n5797;
  assign n5800 = ~n5798 & n5799;
  assign n5801 = x48 & x100;
  assign n5802 = n5800 & n5801;
  assign n5803 = n5800 | n5801;
  assign n5804 = ~n5802 & n5803;
  assign n17700 = n5645 | n5794;
  assign n17701 = (n5644 & n5794) | (n5644 & n17700) | (n5794 & n17700);
  assign n15943 = (n5646 & n5793) | (n5646 & n17701) | (n5793 & n17701);
  assign n12632 = (n5795 & n5797) | (n5795 & n15943) | (n5797 & n15943);
  assign n12633 = n5788 | n12578;
  assign n12634 = (n5788 & n5790) | (n5788 & n12633) | (n5790 & n12633);
  assign n12635 = n5781 | n12580;
  assign n12636 = (n5781 & n5783) | (n5781 & n12635) | (n5783 & n12635);
  assign n15944 = n5774 | n15900;
  assign n15945 = (n5774 & n5776) | (n5774 & n15944) | (n5776 & n15944);
  assign n5809 = n5767 | n5770;
  assign n12637 = n5760 | n5762;
  assign n12638 = (n5653 & n5760) | (n5653 & n12637) | (n5760 & n12637);
  assign n12639 = n5753 | n5755;
  assign n12640 = (n5753 & n12582) | (n5753 & n12639) | (n12582 & n12639);
  assign n12641 = n5746 | n5748;
  assign n12642 = (n5746 & n12584) | (n5746 & n12641) | (n12584 & n12641);
  assign n12643 = n5739 | n5741;
  assign n12644 = (n5739 & n12586) | (n5739 & n12643) | (n12586 & n12643);
  assign n12645 = n5732 | n5734;
  assign n12646 = (n5732 & n12588) | (n5732 & n12645) | (n12588 & n12645);
  assign n12648 = n5711 | n5713;
  assign n15946 = n5562 | n5711;
  assign n15947 = (n5711 & n5713) | (n5711 & n15946) | (n5713 & n15946);
  assign n15948 = (n12565 & n12648) | (n12565 & n15947) | (n12648 & n15947);
  assign n15949 = (n5564 & n12648) | (n5564 & n15947) | (n12648 & n15947);
  assign n15950 = (n12505 & n15948) | (n12505 & n15949) | (n15948 & n15949);
  assign n12653 = n5690 | n5692;
  assign n15951 = n5541 | n5690;
  assign n15952 = (n5690 & n5692) | (n5690 & n15951) | (n5692 & n15951);
  assign n15953 = (n12555 & n12653) | (n12555 & n15952) | (n12653 & n15952);
  assign n15954 = (n12556 & n12653) | (n12556 & n15952) | (n12653 & n15952);
  assign n15955 = (n15840 & n15953) | (n15840 & n15954) | (n15953 & n15954);
  assign n5824 = x69 & x80;
  assign n5825 = x68 & x81;
  assign n5826 = n5824 & n5825;
  assign n5827 = n5824 | n5825;
  assign n5828 = ~n5826 & n5827;
  assign n12659 = n5669 & n5828;
  assign n15956 = (n5828 & n12659) | (n5828 & n15925) | (n12659 & n15925);
  assign n15957 = (n5828 & n12659) | (n5828 & n15923) | (n12659 & n15923);
  assign n15958 = (n15804 & n15956) | (n15804 & n15957) | (n15956 & n15957);
  assign n12661 = n5669 | n5828;
  assign n15959 = n12661 | n15925;
  assign n15960 = n12661 | n15923;
  assign n15961 = (n15804 & n15959) | (n15804 & n15960) | (n15959 & n15960);
  assign n5831 = ~n15958 & n15961;
  assign n5832 = x67 & x82;
  assign n5833 = n5831 & n5832;
  assign n5834 = n5831 | n5832;
  assign n5835 = ~n5833 & n5834;
  assign n12657 = n5676 | n5678;
  assign n12663 = n5835 & n12657;
  assign n12664 = n5676 & n5835;
  assign n12665 = (n15918 & n12663) | (n15918 & n12664) | (n12663 & n12664);
  assign n12666 = n5835 | n12657;
  assign n12667 = n5676 | n5835;
  assign n12668 = (n15918 & n12666) | (n15918 & n12667) | (n12666 & n12667);
  assign n5838 = ~n12665 & n12668;
  assign n5839 = x66 & x83;
  assign n5840 = n5838 & n5839;
  assign n5841 = n5838 | n5839;
  assign n5842 = ~n5840 & n5841;
  assign n12655 = n5683 | n5685;
  assign n12669 = n5842 & n12655;
  assign n12670 = n5683 & n5842;
  assign n12671 = (n15912 & n12669) | (n15912 & n12670) | (n12669 & n12670);
  assign n12672 = n5842 | n12655;
  assign n12673 = n5683 | n5842;
  assign n12674 = (n15912 & n12672) | (n15912 & n12673) | (n12672 & n12673);
  assign n5845 = ~n12671 & n12674;
  assign n5846 = x65 & x84;
  assign n5847 = n5845 & n5846;
  assign n5848 = n5845 | n5846;
  assign n5849 = ~n5847 & n5848;
  assign n5850 = n15955 & n5849;
  assign n5851 = n15955 | n5849;
  assign n5852 = ~n5850 & n5851;
  assign n5853 = x64 & x85;
  assign n5854 = n5852 & n5853;
  assign n5855 = n5852 | n5853;
  assign n5856 = ~n5854 & n5855;
  assign n12650 = n5697 | n5699;
  assign n12675 = n5856 & n12650;
  assign n12676 = n5697 & n5856;
  assign n12677 = (n15905 & n12675) | (n15905 & n12676) | (n12675 & n12676);
  assign n12678 = n5856 | n12650;
  assign n12679 = n5697 | n5856;
  assign n12680 = (n15905 & n12678) | (n15905 & n12679) | (n12678 & n12679);
  assign n5859 = ~n12677 & n12680;
  assign n5860 = x63 & x86;
  assign n5861 = n5859 & n5860;
  assign n5862 = n5859 | n5860;
  assign n5863 = ~n5861 & n5862;
  assign n12681 = n5704 & n5863;
  assign n15962 = (n5863 & n12614) | (n5863 & n12681) | (n12614 & n12681);
  assign n15963 = (n5863 & n12613) | (n5863 & n12681) | (n12613 & n12681);
  assign n15964 = (n15873 & n15962) | (n15873 & n15963) | (n15962 & n15963);
  assign n12683 = n5704 | n5863;
  assign n15965 = n12614 | n12683;
  assign n15966 = n12613 | n12683;
  assign n15967 = (n15873 & n15965) | (n15873 & n15966) | (n15965 & n15966);
  assign n5866 = ~n15964 & n15967;
  assign n5867 = x62 & x87;
  assign n5868 = n5866 & n5867;
  assign n5869 = n5866 | n5867;
  assign n5870 = ~n5868 & n5869;
  assign n5871 = n15950 & n5870;
  assign n5872 = n15950 | n5870;
  assign n5873 = ~n5871 & n5872;
  assign n5874 = x61 & x88;
  assign n5875 = n5873 & n5874;
  assign n5876 = n5873 | n5874;
  assign n5877 = ~n5875 & n5876;
  assign n12685 = n5718 & n5877;
  assign n12686 = (n5877 & n12624) | (n5877 & n12685) | (n12624 & n12685);
  assign n12687 = n5718 | n5877;
  assign n12688 = n12624 | n12687;
  assign n5880 = ~n12686 & n12688;
  assign n5881 = x60 & x89;
  assign n5882 = n5880 & n5881;
  assign n5883 = n5880 | n5881;
  assign n5884 = ~n5882 & n5883;
  assign n12689 = n5725 & n5884;
  assign n12690 = (n5884 & n12628) | (n5884 & n12689) | (n12628 & n12689);
  assign n12691 = n5725 | n5884;
  assign n12692 = n12628 | n12691;
  assign n5887 = ~n12690 & n12692;
  assign n5888 = x59 & x90;
  assign n5889 = n5887 & n5888;
  assign n5890 = n5887 | n5888;
  assign n5891 = ~n5889 & n5890;
  assign n5892 = n12646 & n5891;
  assign n5893 = n12646 | n5891;
  assign n5894 = ~n5892 & n5893;
  assign n5895 = x58 & x91;
  assign n5896 = n5894 & n5895;
  assign n5897 = n5894 | n5895;
  assign n5898 = ~n5896 & n5897;
  assign n5899 = n12644 & n5898;
  assign n5900 = n12644 | n5898;
  assign n5901 = ~n5899 & n5900;
  assign n5902 = x57 & x92;
  assign n5903 = n5901 & n5902;
  assign n5904 = n5901 | n5902;
  assign n5905 = ~n5903 & n5904;
  assign n5906 = n12642 & n5905;
  assign n5907 = n12642 | n5905;
  assign n5908 = ~n5906 & n5907;
  assign n5909 = x56 & x93;
  assign n5910 = n5908 & n5909;
  assign n5911 = n5908 | n5909;
  assign n5912 = ~n5910 & n5911;
  assign n5913 = n12640 & n5912;
  assign n5914 = n12640 | n5912;
  assign n5915 = ~n5913 & n5914;
  assign n5916 = x55 & x94;
  assign n5917 = n5915 & n5916;
  assign n5918 = n5915 | n5916;
  assign n5919 = ~n5917 & n5918;
  assign n5920 = n12638 & n5919;
  assign n5921 = n12638 | n5919;
  assign n5922 = ~n5920 & n5921;
  assign n5923 = x54 & x95;
  assign n5924 = n5922 & n5923;
  assign n5925 = n5922 | n5923;
  assign n5926 = ~n5924 & n5925;
  assign n5927 = n5809 & n5926;
  assign n5928 = n5809 | n5926;
  assign n5929 = ~n5927 & n5928;
  assign n5930 = x53 & x96;
  assign n5931 = n5929 & n5930;
  assign n5932 = n5929 | n5930;
  assign n5933 = ~n5931 & n5932;
  assign n5934 = n15945 & n5933;
  assign n5935 = n15945 | n5933;
  assign n5936 = ~n5934 & n5935;
  assign n5937 = x52 & x97;
  assign n5938 = n5936 & n5937;
  assign n5939 = n5936 | n5937;
  assign n5940 = ~n5938 & n5939;
  assign n5941 = n12636 & n5940;
  assign n5942 = n12636 | n5940;
  assign n5943 = ~n5941 & n5942;
  assign n5944 = x51 & x98;
  assign n5945 = n5943 & n5944;
  assign n5946 = n5943 | n5944;
  assign n5947 = ~n5945 & n5946;
  assign n5948 = n12634 & n5947;
  assign n5949 = n12634 | n5947;
  assign n5950 = ~n5948 & n5949;
  assign n5951 = x50 & x99;
  assign n5952 = n5950 & n5951;
  assign n5953 = n5950 | n5951;
  assign n5954 = ~n5952 & n5953;
  assign n5955 = n12632 & n5954;
  assign n5956 = n12632 | n5954;
  assign n5957 = ~n5955 & n5956;
  assign n5958 = x49 & x100;
  assign n5959 = n5957 & n5958;
  assign n5960 = n5957 | n5958;
  assign n5961 = ~n5959 & n5960;
  assign n5962 = n5802 & n5961;
  assign n5963 = n5802 | n5961;
  assign n5964 = ~n5962 & n5963;
  assign n5965 = x48 & x101;
  assign n5966 = n5964 & n5965;
  assign n5967 = n5964 | n5965;
  assign n5968 = ~n5966 & n5967;
  assign n17702 = n5801 | n5958;
  assign n17703 = (n5800 & n5958) | (n5800 & n17702) | (n5958 & n17702);
  assign n15969 = (n5802 & n5957) | (n5802 & n17703) | (n5957 & n17703);
  assign n12694 = (n5959 & n5961) | (n5959 & n15969) | (n5961 & n15969);
  assign n12695 = n5952 | n12632;
  assign n12696 = (n5952 & n5954) | (n5952 & n12695) | (n5954 & n12695);
  assign n12697 = n5945 | n12634;
  assign n12698 = (n5945 & n5947) | (n5945 & n12697) | (n5947 & n12697);
  assign n12699 = n5938 | n12636;
  assign n12700 = (n5938 & n5940) | (n5938 & n12699) | (n5940 & n12699);
  assign n15970 = n5931 | n15945;
  assign n15971 = (n5931 & n5933) | (n5931 & n15970) | (n5933 & n15970);
  assign n12701 = n5924 | n5926;
  assign n12702 = (n5809 & n5924) | (n5809 & n12701) | (n5924 & n12701);
  assign n12703 = n5917 | n5919;
  assign n12704 = (n5917 & n12638) | (n5917 & n12703) | (n12638 & n12703);
  assign n12705 = n5910 | n5912;
  assign n12706 = (n5910 & n12640) | (n5910 & n12705) | (n12640 & n12705);
  assign n12707 = n5903 | n5905;
  assign n12708 = (n5903 & n12642) | (n5903 & n12707) | (n12642 & n12707);
  assign n12709 = n5896 | n5898;
  assign n12710 = (n5896 & n12644) | (n5896 & n12709) | (n12644 & n12709);
  assign n12711 = n5889 | n5891;
  assign n12712 = (n5889 & n12646) | (n5889 & n12711) | (n12646 & n12711);
  assign n12716 = n5861 | n5863;
  assign n15972 = n5704 | n5861;
  assign n15973 = (n5861 & n5863) | (n5861 & n15972) | (n5863 & n15972);
  assign n15974 = (n12614 & n12716) | (n12614 & n15973) | (n12716 & n15973);
  assign n15975 = (n12613 & n12716) | (n12613 & n15973) | (n12716 & n15973);
  assign n15976 = (n15873 & n15974) | (n15873 & n15975) | (n15974 & n15975);
  assign n5989 = x70 & x80;
  assign n5990 = x69 & x81;
  assign n5991 = n5989 & n5990;
  assign n5992 = n5989 | n5990;
  assign n5993 = ~n5991 & n5992;
  assign n15981 = n5669 | n5826;
  assign n15982 = (n5826 & n5828) | (n5826 & n15981) | (n5828 & n15981);
  assign n12729 = n5993 & n15982;
  assign n12727 = n5826 | n5828;
  assign n12730 = n5993 & n12727;
  assign n15983 = (n12729 & n12730) | (n12729 & n15925) | (n12730 & n15925);
  assign n15984 = (n12729 & n12730) | (n12729 & n15923) | (n12730 & n15923);
  assign n15985 = (n15804 & n15983) | (n15804 & n15984) | (n15983 & n15984);
  assign n12732 = n5993 | n15982;
  assign n12733 = n5993 | n12727;
  assign n15986 = (n12732 & n12733) | (n12732 & n15925) | (n12733 & n15925);
  assign n15987 = (n12732 & n12733) | (n12732 & n15923) | (n12733 & n15923);
  assign n15988 = (n15804 & n15986) | (n15804 & n15987) | (n15986 & n15987);
  assign n5996 = ~n15985 & n15988;
  assign n5997 = x68 & x82;
  assign n5998 = n5996 & n5997;
  assign n5999 = n5996 | n5997;
  assign n6000 = ~n5998 & n5999;
  assign n15989 = n5833 | n5835;
  assign n15990 = (n5833 & n12657) | (n5833 & n15989) | (n12657 & n15989);
  assign n12735 = n6000 & n15990;
  assign n15991 = n5676 | n5833;
  assign n15992 = (n5833 & n5835) | (n5833 & n15991) | (n5835 & n15991);
  assign n12736 = n6000 & n15992;
  assign n12737 = (n15918 & n12735) | (n15918 & n12736) | (n12735 & n12736);
  assign n12738 = n6000 | n15990;
  assign n12739 = n6000 | n15992;
  assign n12740 = (n15918 & n12738) | (n15918 & n12739) | (n12738 & n12739);
  assign n6003 = ~n12737 & n12740;
  assign n6004 = x67 & x83;
  assign n6005 = n6003 & n6004;
  assign n6006 = n6003 | n6004;
  assign n6007 = ~n6005 & n6006;
  assign n15977 = n5840 | n5842;
  assign n15978 = (n5840 & n12655) | (n5840 & n15977) | (n12655 & n15977);
  assign n15993 = n6007 & n15978;
  assign n15979 = n5683 | n5840;
  assign n15980 = (n5840 & n5842) | (n5840 & n15979) | (n5842 & n15979);
  assign n15994 = n6007 & n15980;
  assign n15995 = (n15912 & n15993) | (n15912 & n15994) | (n15993 & n15994);
  assign n15996 = n6007 | n15978;
  assign n15997 = n6007 | n15980;
  assign n15998 = (n15912 & n15996) | (n15912 & n15997) | (n15996 & n15997);
  assign n6010 = ~n15995 & n15998;
  assign n6011 = x66 & x84;
  assign n6012 = n6010 & n6011;
  assign n6013 = n6010 | n6011;
  assign n6014 = ~n6012 & n6013;
  assign n12718 = n5847 | n5849;
  assign n12741 = n6014 & n12718;
  assign n12742 = n5847 & n6014;
  assign n12743 = (n15955 & n12741) | (n15955 & n12742) | (n12741 & n12742);
  assign n12744 = n6014 | n12718;
  assign n12745 = n5847 | n6014;
  assign n12746 = (n15955 & n12744) | (n15955 & n12745) | (n12744 & n12745);
  assign n6017 = ~n12743 & n12746;
  assign n6018 = x65 & x85;
  assign n6019 = n6017 & n6018;
  assign n6020 = n6017 | n6018;
  assign n6021 = ~n6019 & n6020;
  assign n12747 = n5854 & n6021;
  assign n15999 = (n6021 & n12676) | (n6021 & n12747) | (n12676 & n12747);
  assign n16000 = (n6021 & n12675) | (n6021 & n12747) | (n12675 & n12747);
  assign n16001 = (n15905 & n15999) | (n15905 & n16000) | (n15999 & n16000);
  assign n12749 = n5854 | n6021;
  assign n16002 = n12676 | n12749;
  assign n16003 = n12675 | n12749;
  assign n16004 = (n15905 & n16002) | (n15905 & n16003) | (n16002 & n16003);
  assign n6024 = ~n16001 & n16004;
  assign n6025 = x64 & x86;
  assign n6026 = n6024 & n6025;
  assign n6027 = n6024 | n6025;
  assign n6028 = ~n6026 & n6027;
  assign n6029 = n15976 & n6028;
  assign n6030 = n15976 | n6028;
  assign n6031 = ~n6029 & n6030;
  assign n6032 = x63 & x87;
  assign n6033 = n6031 & n6032;
  assign n6034 = n6031 | n6032;
  assign n6035 = ~n6033 & n6034;
  assign n12713 = n5868 | n5870;
  assign n12751 = n6035 & n12713;
  assign n12752 = n5868 & n6035;
  assign n12753 = (n15950 & n12751) | (n15950 & n12752) | (n12751 & n12752);
  assign n12754 = n6035 | n12713;
  assign n12755 = n5868 | n6035;
  assign n12756 = (n15950 & n12754) | (n15950 & n12755) | (n12754 & n12755);
  assign n6038 = ~n12753 & n12756;
  assign n6039 = x62 & x88;
  assign n6040 = n6038 & n6039;
  assign n6041 = n6038 | n6039;
  assign n6042 = ~n6040 & n6041;
  assign n12757 = n5875 & n6042;
  assign n16005 = (n6042 & n12685) | (n6042 & n12757) | (n12685 & n12757);
  assign n16006 = (n5877 & n6042) | (n5877 & n12757) | (n6042 & n12757);
  assign n16007 = (n12624 & n16005) | (n12624 & n16006) | (n16005 & n16006);
  assign n12759 = n5875 | n6042;
  assign n16008 = n12685 | n12759;
  assign n16009 = n5877 | n12759;
  assign n16010 = (n12624 & n16008) | (n12624 & n16009) | (n16008 & n16009);
  assign n6045 = ~n16007 & n16010;
  assign n6046 = x61 & x89;
  assign n6047 = n6045 & n6046;
  assign n6048 = n6045 | n6046;
  assign n6049 = ~n6047 & n6048;
  assign n12761 = n5882 & n6049;
  assign n12762 = (n6049 & n12690) | (n6049 & n12761) | (n12690 & n12761);
  assign n12763 = n5882 | n6049;
  assign n12764 = n12690 | n12763;
  assign n6052 = ~n12762 & n12764;
  assign n6053 = x60 & x90;
  assign n6054 = n6052 & n6053;
  assign n6055 = n6052 | n6053;
  assign n6056 = ~n6054 & n6055;
  assign n6057 = n12712 & n6056;
  assign n6058 = n12712 | n6056;
  assign n6059 = ~n6057 & n6058;
  assign n6060 = x59 & x91;
  assign n6061 = n6059 & n6060;
  assign n6062 = n6059 | n6060;
  assign n6063 = ~n6061 & n6062;
  assign n6064 = n12710 & n6063;
  assign n6065 = n12710 | n6063;
  assign n6066 = ~n6064 & n6065;
  assign n6067 = x58 & x92;
  assign n6068 = n6066 & n6067;
  assign n6069 = n6066 | n6067;
  assign n6070 = ~n6068 & n6069;
  assign n6071 = n12708 & n6070;
  assign n6072 = n12708 | n6070;
  assign n6073 = ~n6071 & n6072;
  assign n6074 = x57 & x93;
  assign n6075 = n6073 & n6074;
  assign n6076 = n6073 | n6074;
  assign n6077 = ~n6075 & n6076;
  assign n6078 = n12706 & n6077;
  assign n6079 = n12706 | n6077;
  assign n6080 = ~n6078 & n6079;
  assign n6081 = x56 & x94;
  assign n6082 = n6080 & n6081;
  assign n6083 = n6080 | n6081;
  assign n6084 = ~n6082 & n6083;
  assign n6085 = n12704 & n6084;
  assign n6086 = n12704 | n6084;
  assign n6087 = ~n6085 & n6086;
  assign n6088 = x55 & x95;
  assign n6089 = n6087 & n6088;
  assign n6090 = n6087 | n6088;
  assign n6091 = ~n6089 & n6090;
  assign n6092 = n12702 & n6091;
  assign n6093 = n12702 | n6091;
  assign n6094 = ~n6092 & n6093;
  assign n6095 = x54 & x96;
  assign n6096 = n6094 & n6095;
  assign n6097 = n6094 | n6095;
  assign n6098 = ~n6096 & n6097;
  assign n6099 = n15971 & n6098;
  assign n6100 = n15971 | n6098;
  assign n6101 = ~n6099 & n6100;
  assign n6102 = x53 & x97;
  assign n6103 = n6101 & n6102;
  assign n6104 = n6101 | n6102;
  assign n6105 = ~n6103 & n6104;
  assign n6106 = n12700 & n6105;
  assign n6107 = n12700 | n6105;
  assign n6108 = ~n6106 & n6107;
  assign n6109 = x52 & x98;
  assign n6110 = n6108 & n6109;
  assign n6111 = n6108 | n6109;
  assign n6112 = ~n6110 & n6111;
  assign n6113 = n12698 & n6112;
  assign n6114 = n12698 | n6112;
  assign n6115 = ~n6113 & n6114;
  assign n6116 = x51 & x99;
  assign n6117 = n6115 & n6116;
  assign n6118 = n6115 | n6116;
  assign n6119 = ~n6117 & n6118;
  assign n6120 = n12696 & n6119;
  assign n6121 = n12696 | n6119;
  assign n6122 = ~n6120 & n6121;
  assign n6123 = x50 & x100;
  assign n6124 = n6122 & n6123;
  assign n6125 = n6122 | n6123;
  assign n6126 = ~n6124 & n6125;
  assign n6127 = n12694 & n6126;
  assign n6128 = n12694 | n6126;
  assign n6129 = ~n6127 & n6128;
  assign n6130 = x49 & x101;
  assign n6131 = n6129 & n6130;
  assign n6132 = n6129 | n6130;
  assign n6133 = ~n6131 & n6132;
  assign n6134 = n5966 & n6133;
  assign n6135 = n5966 | n6133;
  assign n6136 = ~n6134 & n6135;
  assign n6137 = x48 & x102;
  assign n6138 = n6136 & n6137;
  assign n6139 = n6136 | n6137;
  assign n6140 = ~n6138 & n6139;
  assign n12765 = n5966 | n6131;
  assign n12766 = (n6131 & n6133) | (n6131 & n12765) | (n6133 & n12765);
  assign n12767 = n6124 | n12694;
  assign n12768 = (n6124 & n6126) | (n6124 & n12767) | (n6126 & n12767);
  assign n12769 = n6117 | n12696;
  assign n12770 = (n6117 & n6119) | (n6117 & n12769) | (n6119 & n12769);
  assign n12771 = n6110 | n12698;
  assign n12772 = (n6110 & n6112) | (n6110 & n12771) | (n6112 & n12771);
  assign n12773 = n6103 | n12700;
  assign n12774 = (n6103 & n6105) | (n6103 & n12773) | (n6105 & n12773);
  assign n12775 = n6096 | n6098;
  assign n12776 = (n15971 & n6096) | (n15971 & n12775) | (n6096 & n12775);
  assign n12777 = n6089 | n6091;
  assign n12778 = (n6089 & n12702) | (n6089 & n12777) | (n12702 & n12777);
  assign n12779 = n6082 | n6084;
  assign n12780 = (n6082 & n12704) | (n6082 & n12779) | (n12704 & n12779);
  assign n12781 = n6075 | n6077;
  assign n12782 = (n6075 & n12706) | (n6075 & n12781) | (n12706 & n12781);
  assign n12783 = n6068 | n6070;
  assign n12784 = (n6068 & n12708) | (n6068 & n12783) | (n12708 & n12783);
  assign n12785 = n6061 | n6063;
  assign n12786 = (n6061 & n12710) | (n6061 & n12785) | (n12710 & n12785);
  assign n12787 = n6054 | n6056;
  assign n12788 = (n6054 & n12712) | (n6054 & n12787) | (n12712 & n12787);
  assign n12790 = n6040 | n6042;
  assign n16011 = n5875 | n6040;
  assign n16012 = (n6040 & n6042) | (n6040 & n16011) | (n6042 & n16011);
  assign n16013 = (n12685 & n12790) | (n12685 & n16012) | (n12790 & n16012);
  assign n16014 = (n5877 & n12790) | (n5877 & n16012) | (n12790 & n16012);
  assign n16015 = (n12624 & n16013) | (n12624 & n16014) | (n16013 & n16014);
  assign n12795 = n6019 | n6021;
  assign n16016 = n5854 | n6019;
  assign n16017 = (n6019 & n6021) | (n6019 & n16016) | (n6021 & n16016);
  assign n16018 = (n12676 & n12795) | (n12676 & n16017) | (n12795 & n16017);
  assign n16019 = (n12675 & n12795) | (n12675 & n16017) | (n12795 & n16017);
  assign n16020 = (n15905 & n16018) | (n15905 & n16019) | (n16018 & n16019);
  assign n6162 = x71 & x80;
  assign n6163 = x70 & x81;
  assign n6164 = n6162 & n6163;
  assign n6165 = n6162 | n6163;
  assign n6166 = ~n6164 & n6165;
  assign n16028 = n5991 | n5993;
  assign n16029 = (n5991 & n15982) | (n5991 & n16028) | (n15982 & n16028);
  assign n12808 = n6166 & n16029;
  assign n16030 = (n5991 & n12727) | (n5991 & n16028) | (n12727 & n16028);
  assign n12809 = n6166 & n16030;
  assign n16031 = (n12808 & n12809) | (n12808 & n15925) | (n12809 & n15925);
  assign n16032 = (n12808 & n12809) | (n12808 & n15923) | (n12809 & n15923);
  assign n16033 = (n15804 & n16031) | (n15804 & n16032) | (n16031 & n16032);
  assign n12811 = n6166 | n16029;
  assign n12812 = n6166 | n16030;
  assign n16034 = (n12811 & n12812) | (n12811 & n15925) | (n12812 & n15925);
  assign n16035 = (n12811 & n12812) | (n12811 & n15923) | (n12812 & n15923);
  assign n16036 = (n15804 & n16034) | (n15804 & n16035) | (n16034 & n16035);
  assign n6169 = ~n16033 & n16036;
  assign n6170 = x69 & x82;
  assign n6171 = n6169 & n6170;
  assign n6172 = n6169 | n6170;
  assign n6173 = ~n6171 & n6172;
  assign n16025 = n5998 | n6000;
  assign n17704 = n6173 & n16025;
  assign n17705 = n5998 & n6173;
  assign n17706 = (n15990 & n17704) | (n15990 & n17705) | (n17704 & n17705);
  assign n16026 = (n5998 & n15992) | (n5998 & n16025) | (n15992 & n16025);
  assign n16038 = n6173 & n16026;
  assign n16039 = (n15918 & n17706) | (n15918 & n16038) | (n17706 & n16038);
  assign n17707 = n6173 | n16025;
  assign n17708 = n5998 | n6173;
  assign n17709 = (n15990 & n17707) | (n15990 & n17708) | (n17707 & n17708);
  assign n16041 = n6173 | n16026;
  assign n16042 = (n15918 & n17709) | (n15918 & n16041) | (n17709 & n16041);
  assign n6176 = ~n16039 & n16042;
  assign n6177 = x68 & x83;
  assign n6178 = n6176 & n6177;
  assign n6179 = n6176 | n6177;
  assign n6180 = ~n6178 & n6179;
  assign n12800 = n6005 | n6007;
  assign n12814 = n6180 & n12800;
  assign n12815 = n6005 & n6180;
  assign n16043 = (n12814 & n12815) | (n12814 & n15978) | (n12815 & n15978);
  assign n16044 = (n12814 & n12815) | (n12814 & n15980) | (n12815 & n15980);
  assign n16045 = (n15912 & n16043) | (n15912 & n16044) | (n16043 & n16044);
  assign n12817 = n6180 | n12800;
  assign n12818 = n6005 | n6180;
  assign n16046 = (n12817 & n12818) | (n12817 & n15978) | (n12818 & n15978);
  assign n16047 = (n12817 & n12818) | (n12817 & n15980) | (n12818 & n15980);
  assign n16048 = (n15912 & n16046) | (n15912 & n16047) | (n16046 & n16047);
  assign n6183 = ~n16045 & n16048;
  assign n6184 = x67 & x84;
  assign n6185 = n6183 & n6184;
  assign n6186 = n6183 | n6184;
  assign n6187 = ~n6185 & n6186;
  assign n16023 = n6012 | n6014;
  assign n16024 = (n6012 & n12718) | (n6012 & n16023) | (n12718 & n16023);
  assign n16049 = n6187 & n16024;
  assign n16021 = n5847 | n6012;
  assign n16022 = (n6012 & n6014) | (n6012 & n16021) | (n6014 & n16021);
  assign n16050 = n6187 & n16022;
  assign n16051 = (n15955 & n16049) | (n15955 & n16050) | (n16049 & n16050);
  assign n16052 = n6187 | n16024;
  assign n16053 = n6187 | n16022;
  assign n16054 = (n15955 & n16052) | (n15955 & n16053) | (n16052 & n16053);
  assign n6190 = ~n16051 & n16054;
  assign n6191 = x66 & x85;
  assign n6192 = n6190 & n6191;
  assign n6193 = n6190 | n6191;
  assign n6194 = ~n6192 & n6193;
  assign n6195 = n16020 & n6194;
  assign n6196 = n16020 | n6194;
  assign n6197 = ~n6195 & n6196;
  assign n6198 = x65 & x86;
  assign n6199 = n6197 & n6198;
  assign n6200 = n6197 | n6198;
  assign n6201 = ~n6199 & n6200;
  assign n12792 = n6026 | n6028;
  assign n12820 = n6201 & n12792;
  assign n12821 = n6026 & n6201;
  assign n12822 = (n15976 & n12820) | (n15976 & n12821) | (n12820 & n12821);
  assign n12823 = n6201 | n12792;
  assign n12824 = n6026 | n6201;
  assign n12825 = (n15976 & n12823) | (n15976 & n12824) | (n12823 & n12824);
  assign n6204 = ~n12822 & n12825;
  assign n6205 = x64 & x87;
  assign n6206 = n6204 & n6205;
  assign n6207 = n6204 | n6205;
  assign n6208 = ~n6206 & n6207;
  assign n12826 = n6033 & n6208;
  assign n16055 = (n6208 & n12752) | (n6208 & n12826) | (n12752 & n12826);
  assign n16056 = (n6208 & n12751) | (n6208 & n12826) | (n12751 & n12826);
  assign n16057 = (n15950 & n16055) | (n15950 & n16056) | (n16055 & n16056);
  assign n12828 = n6033 | n6208;
  assign n16058 = n12752 | n12828;
  assign n16059 = n12751 | n12828;
  assign n16060 = (n15950 & n16058) | (n15950 & n16059) | (n16058 & n16059);
  assign n6211 = ~n16057 & n16060;
  assign n6212 = x63 & x88;
  assign n6213 = n6211 & n6212;
  assign n6214 = n6211 | n6212;
  assign n6215 = ~n6213 & n6214;
  assign n6216 = n16015 & n6215;
  assign n6217 = n16015 | n6215;
  assign n6218 = ~n6216 & n6217;
  assign n6219 = x62 & x89;
  assign n6220 = n6218 & n6219;
  assign n6221 = n6218 | n6219;
  assign n6222 = ~n6220 & n6221;
  assign n12830 = n6047 & n6222;
  assign n12831 = (n6222 & n12762) | (n6222 & n12830) | (n12762 & n12830);
  assign n12832 = n6047 | n6222;
  assign n12833 = n12762 | n12832;
  assign n6225 = ~n12831 & n12833;
  assign n6226 = x61 & x90;
  assign n6227 = n6225 & n6226;
  assign n6228 = n6225 | n6226;
  assign n6229 = ~n6227 & n6228;
  assign n6230 = n12788 & n6229;
  assign n6231 = n12788 | n6229;
  assign n6232 = ~n6230 & n6231;
  assign n6233 = x60 & x91;
  assign n6234 = n6232 & n6233;
  assign n6235 = n6232 | n6233;
  assign n6236 = ~n6234 & n6235;
  assign n6237 = n12786 & n6236;
  assign n6238 = n12786 | n6236;
  assign n6239 = ~n6237 & n6238;
  assign n6240 = x59 & x92;
  assign n6241 = n6239 & n6240;
  assign n6242 = n6239 | n6240;
  assign n6243 = ~n6241 & n6242;
  assign n6244 = n12784 & n6243;
  assign n6245 = n12784 | n6243;
  assign n6246 = ~n6244 & n6245;
  assign n6247 = x58 & x93;
  assign n6248 = n6246 & n6247;
  assign n6249 = n6246 | n6247;
  assign n6250 = ~n6248 & n6249;
  assign n6251 = n12782 & n6250;
  assign n6252 = n12782 | n6250;
  assign n6253 = ~n6251 & n6252;
  assign n6254 = x57 & x94;
  assign n6255 = n6253 & n6254;
  assign n6256 = n6253 | n6254;
  assign n6257 = ~n6255 & n6256;
  assign n6258 = n12780 & n6257;
  assign n6259 = n12780 | n6257;
  assign n6260 = ~n6258 & n6259;
  assign n6261 = x56 & x95;
  assign n6262 = n6260 & n6261;
  assign n6263 = n6260 | n6261;
  assign n6264 = ~n6262 & n6263;
  assign n6265 = n12778 & n6264;
  assign n6266 = n12778 | n6264;
  assign n6267 = ~n6265 & n6266;
  assign n6268 = x55 & x96;
  assign n6269 = n6267 & n6268;
  assign n6270 = n6267 | n6268;
  assign n6271 = ~n6269 & n6270;
  assign n6272 = n12776 & n6271;
  assign n6273 = n12776 | n6271;
  assign n6274 = ~n6272 & n6273;
  assign n6275 = x54 & x97;
  assign n6276 = n6274 & n6275;
  assign n6277 = n6274 | n6275;
  assign n6278 = ~n6276 & n6277;
  assign n6279 = n12774 & n6278;
  assign n6280 = n12774 | n6278;
  assign n6281 = ~n6279 & n6280;
  assign n6282 = x53 & x98;
  assign n6283 = n6281 & n6282;
  assign n6284 = n6281 | n6282;
  assign n6285 = ~n6283 & n6284;
  assign n6286 = n12772 & n6285;
  assign n6287 = n12772 | n6285;
  assign n6288 = ~n6286 & n6287;
  assign n6289 = x52 & x99;
  assign n6290 = n6288 & n6289;
  assign n6291 = n6288 | n6289;
  assign n6292 = ~n6290 & n6291;
  assign n6293 = n12770 & n6292;
  assign n6294 = n12770 | n6292;
  assign n6295 = ~n6293 & n6294;
  assign n6296 = x51 & x100;
  assign n6297 = n6295 & n6296;
  assign n6298 = n6295 | n6296;
  assign n6299 = ~n6297 & n6298;
  assign n6300 = n12768 & n6299;
  assign n6301 = n12768 | n6299;
  assign n6302 = ~n6300 & n6301;
  assign n6303 = x50 & x101;
  assign n6304 = n6302 & n6303;
  assign n6305 = n6302 | n6303;
  assign n6306 = ~n6304 & n6305;
  assign n6307 = n12766 & n6306;
  assign n6308 = n12766 | n6306;
  assign n6309 = ~n6307 & n6308;
  assign n6310 = x49 & x102;
  assign n6311 = n6309 & n6310;
  assign n6312 = n6309 | n6310;
  assign n6313 = ~n6311 & n6312;
  assign n6314 = n6138 & n6313;
  assign n6315 = n6138 | n6313;
  assign n6316 = ~n6314 & n6315;
  assign n6317 = x48 & x103;
  assign n6318 = n6316 & n6317;
  assign n6319 = n6316 | n6317;
  assign n6320 = ~n6318 & n6319;
  assign n17710 = n6137 | n6310;
  assign n17711 = (n6136 & n6310) | (n6136 & n17710) | (n6310 & n17710);
  assign n16062 = (n6138 & n6309) | (n6138 & n17711) | (n6309 & n17711);
  assign n12835 = (n6311 & n6313) | (n6311 & n16062) | (n6313 & n16062);
  assign n16063 = n6304 | n12766;
  assign n16064 = (n6304 & n6306) | (n6304 & n16063) | (n6306 & n16063);
  assign n6323 = n6297 | n6300;
  assign n6324 = n6290 | n6293;
  assign n6325 = n6283 | n6286;
  assign n6326 = n6276 | n6279;
  assign n12836 = n6269 | n6271;
  assign n12837 = (n6269 & n12776) | (n6269 & n12836) | (n12776 & n12836);
  assign n12838 = n6262 | n6264;
  assign n12839 = (n6262 & n12778) | (n6262 & n12838) | (n12778 & n12838);
  assign n12840 = n6255 | n6257;
  assign n12841 = (n6255 & n12780) | (n6255 & n12840) | (n12780 & n12840);
  assign n12842 = n6248 | n6250;
  assign n12843 = (n6248 & n12782) | (n6248 & n12842) | (n12782 & n12842);
  assign n12844 = n6241 | n6243;
  assign n12845 = (n6241 & n12784) | (n6241 & n12844) | (n12784 & n12844);
  assign n12846 = n6234 | n6236;
  assign n12847 = (n6234 & n12786) | (n6234 & n12846) | (n12786 & n12846);
  assign n12848 = n6227 | n6229;
  assign n12849 = (n6227 & n12788) | (n6227 & n12848) | (n12788 & n12848);
  assign n12853 = n6206 | n6208;
  assign n16065 = n6033 | n6206;
  assign n16066 = (n6206 & n6208) | (n6206 & n16065) | (n6208 & n16065);
  assign n16067 = (n12752 & n12853) | (n12752 & n16066) | (n12853 & n16066);
  assign n16068 = (n12751 & n12853) | (n12751 & n16066) | (n12853 & n16066);
  assign n16069 = (n15950 & n16067) | (n15950 & n16068) | (n16067 & n16068);
  assign n12722 = (n15912 & n15978) | (n15912 & n15980) | (n15978 & n15980);
  assign n6343 = x72 & x80;
  assign n6344 = x71 & x81;
  assign n6345 = n6343 & n6344;
  assign n6346 = n6343 | n6344;
  assign n6347 = ~n6345 & n6346;
  assign n16070 = n6164 | n6166;
  assign n16072 = n6347 & n16070;
  assign n16073 = n6164 & n6347;
  assign n16074 = (n16029 & n16072) | (n16029 & n16073) | (n16072 & n16073);
  assign n16076 = (n16030 & n16072) | (n16030 & n16073) | (n16072 & n16073);
  assign n16077 = (n15925 & n16074) | (n15925 & n16076) | (n16074 & n16076);
  assign n16078 = (n15923 & n16074) | (n15923 & n16076) | (n16074 & n16076);
  assign n16079 = (n15804 & n16077) | (n15804 & n16078) | (n16077 & n16078);
  assign n16080 = n6347 | n16070;
  assign n16081 = n6164 | n6347;
  assign n16082 = (n16029 & n16080) | (n16029 & n16081) | (n16080 & n16081);
  assign n16083 = (n16030 & n16080) | (n16030 & n16081) | (n16080 & n16081);
  assign n16084 = (n15925 & n16082) | (n15925 & n16083) | (n16082 & n16083);
  assign n16085 = (n15923 & n16082) | (n15923 & n16083) | (n16082 & n16083);
  assign n16086 = (n15804 & n16084) | (n15804 & n16085) | (n16084 & n16085);
  assign n6350 = ~n16079 & n16086;
  assign n6351 = x70 & x82;
  assign n6352 = n6350 & n6351;
  assign n6353 = n6350 | n6351;
  assign n6354 = ~n6352 & n6353;
  assign n12862 = n6171 | n6173;
  assign n12873 = n6354 & n12862;
  assign n12874 = n6171 & n6354;
  assign n16027 = (n5998 & n15990) | (n5998 & n16025) | (n15990 & n16025);
  assign n16087 = (n12873 & n12874) | (n12873 & n16027) | (n12874 & n16027);
  assign n16088 = (n12873 & n12874) | (n12873 & n16026) | (n12874 & n16026);
  assign n16089 = (n15918 & n16087) | (n15918 & n16088) | (n16087 & n16088);
  assign n12876 = n6354 | n12862;
  assign n12877 = n6171 | n6354;
  assign n16090 = (n12876 & n12877) | (n12876 & n16027) | (n12877 & n16027);
  assign n16091 = (n12876 & n12877) | (n12876 & n16026) | (n12877 & n16026);
  assign n16092 = (n15918 & n16090) | (n15918 & n16091) | (n16090 & n16091);
  assign n6357 = ~n16089 & n16092;
  assign n6358 = x69 & x83;
  assign n6359 = n6357 & n6358;
  assign n6360 = n6357 | n6358;
  assign n6361 = ~n6359 & n6360;
  assign n16093 = n6178 | n6180;
  assign n16094 = (n6178 & n12800) | (n6178 & n16093) | (n12800 & n16093);
  assign n12879 = n6361 & n16094;
  assign n16095 = n6005 | n6178;
  assign n16096 = (n6178 & n6180) | (n6178 & n16095) | (n6180 & n16095);
  assign n12880 = n6361 & n16096;
  assign n12881 = (n12722 & n12879) | (n12722 & n12880) | (n12879 & n12880);
  assign n12882 = n6361 | n16094;
  assign n12883 = n6361 | n16096;
  assign n12884 = (n12722 & n12882) | (n12722 & n12883) | (n12882 & n12883);
  assign n6364 = ~n12881 & n12884;
  assign n6365 = x68 & x84;
  assign n6366 = n6364 & n6365;
  assign n6367 = n6364 | n6365;
  assign n6368 = ~n6366 & n6367;
  assign n12857 = n6185 | n6187;
  assign n12885 = n6368 & n12857;
  assign n12886 = n6185 & n6368;
  assign n16097 = (n12885 & n12886) | (n12885 & n16024) | (n12886 & n16024);
  assign n16098 = (n12885 & n12886) | (n12885 & n16022) | (n12886 & n16022);
  assign n16099 = (n15955 & n16097) | (n15955 & n16098) | (n16097 & n16098);
  assign n12888 = n6368 | n12857;
  assign n12889 = n6185 | n6368;
  assign n16100 = (n12888 & n12889) | (n12888 & n16024) | (n12889 & n16024);
  assign n16101 = (n12888 & n12889) | (n12888 & n16022) | (n12889 & n16022);
  assign n16102 = (n15955 & n16100) | (n15955 & n16101) | (n16100 & n16101);
  assign n6371 = ~n16099 & n16102;
  assign n6372 = x67 & x85;
  assign n6373 = n6371 & n6372;
  assign n6374 = n6371 | n6372;
  assign n6375 = ~n6373 & n6374;
  assign n12855 = n6192 | n6194;
  assign n12891 = n6375 & n12855;
  assign n12892 = n6192 & n6375;
  assign n12893 = (n16020 & n12891) | (n16020 & n12892) | (n12891 & n12892);
  assign n12894 = n6375 | n12855;
  assign n12895 = n6192 | n6375;
  assign n12896 = (n16020 & n12894) | (n16020 & n12895) | (n12894 & n12895);
  assign n6378 = ~n12893 & n12896;
  assign n6379 = x66 & x86;
  assign n6380 = n6378 & n6379;
  assign n6381 = n6378 | n6379;
  assign n6382 = ~n6380 & n6381;
  assign n12897 = n6199 & n6382;
  assign n16103 = (n6382 & n12821) | (n6382 & n12897) | (n12821 & n12897);
  assign n16104 = (n6382 & n12820) | (n6382 & n12897) | (n12820 & n12897);
  assign n16105 = (n15976 & n16103) | (n15976 & n16104) | (n16103 & n16104);
  assign n12899 = n6199 | n6382;
  assign n16106 = n12821 | n12899;
  assign n16107 = n12820 | n12899;
  assign n16108 = (n15976 & n16106) | (n15976 & n16107) | (n16106 & n16107);
  assign n6385 = ~n16105 & n16108;
  assign n6386 = x65 & x87;
  assign n6387 = n6385 & n6386;
  assign n6388 = n6385 | n6386;
  assign n6389 = ~n6387 & n6388;
  assign n6390 = n16069 & n6389;
  assign n6391 = n16069 | n6389;
  assign n6392 = ~n6390 & n6391;
  assign n6393 = x64 & x88;
  assign n6394 = n6392 & n6393;
  assign n6395 = n6392 | n6393;
  assign n6396 = ~n6394 & n6395;
  assign n12850 = n6213 | n6215;
  assign n12901 = n6396 & n12850;
  assign n12902 = n6213 & n6396;
  assign n12903 = (n16015 & n12901) | (n16015 & n12902) | (n12901 & n12902);
  assign n12904 = n6396 | n12850;
  assign n12905 = n6213 | n6396;
  assign n12906 = (n16015 & n12904) | (n16015 & n12905) | (n12904 & n12905);
  assign n6399 = ~n12903 & n12906;
  assign n6400 = x63 & x89;
  assign n6401 = n6399 & n6400;
  assign n6402 = n6399 | n6400;
  assign n6403 = ~n6401 & n6402;
  assign n12907 = n6220 & n6403;
  assign n16109 = (n6403 & n12830) | (n6403 & n12907) | (n12830 & n12907);
  assign n16110 = (n6222 & n6403) | (n6222 & n12907) | (n6403 & n12907);
  assign n16111 = (n12762 & n16109) | (n12762 & n16110) | (n16109 & n16110);
  assign n12909 = n6220 | n6403;
  assign n16112 = n12830 | n12909;
  assign n16113 = n6222 | n12909;
  assign n16114 = (n12762 & n16112) | (n12762 & n16113) | (n16112 & n16113);
  assign n6406 = ~n16111 & n16114;
  assign n6407 = x62 & x90;
  assign n6408 = n6406 & n6407;
  assign n6409 = n6406 | n6407;
  assign n6410 = ~n6408 & n6409;
  assign n6411 = n12849 & n6410;
  assign n6412 = n12849 | n6410;
  assign n6413 = ~n6411 & n6412;
  assign n6414 = x61 & x91;
  assign n6415 = n6413 & n6414;
  assign n6416 = n6413 | n6414;
  assign n6417 = ~n6415 & n6416;
  assign n6418 = n12847 & n6417;
  assign n6419 = n12847 | n6417;
  assign n6420 = ~n6418 & n6419;
  assign n6421 = x60 & x92;
  assign n6422 = n6420 & n6421;
  assign n6423 = n6420 | n6421;
  assign n6424 = ~n6422 & n6423;
  assign n6425 = n12845 & n6424;
  assign n6426 = n12845 | n6424;
  assign n6427 = ~n6425 & n6426;
  assign n6428 = x59 & x93;
  assign n6429 = n6427 & n6428;
  assign n6430 = n6427 | n6428;
  assign n6431 = ~n6429 & n6430;
  assign n6432 = n12843 & n6431;
  assign n6433 = n12843 | n6431;
  assign n6434 = ~n6432 & n6433;
  assign n6435 = x58 & x94;
  assign n6436 = n6434 & n6435;
  assign n6437 = n6434 | n6435;
  assign n6438 = ~n6436 & n6437;
  assign n6439 = n12841 & n6438;
  assign n6440 = n12841 | n6438;
  assign n6441 = ~n6439 & n6440;
  assign n6442 = x57 & x95;
  assign n6443 = n6441 & n6442;
  assign n6444 = n6441 | n6442;
  assign n6445 = ~n6443 & n6444;
  assign n6446 = n12839 & n6445;
  assign n6447 = n12839 | n6445;
  assign n6448 = ~n6446 & n6447;
  assign n6449 = x56 & x96;
  assign n6450 = n6448 & n6449;
  assign n6451 = n6448 | n6449;
  assign n6452 = ~n6450 & n6451;
  assign n6453 = n12837 & n6452;
  assign n6454 = n12837 | n6452;
  assign n6455 = ~n6453 & n6454;
  assign n6456 = x55 & x97;
  assign n6457 = n6455 & n6456;
  assign n6458 = n6455 | n6456;
  assign n6459 = ~n6457 & n6458;
  assign n6460 = n6326 & n6459;
  assign n6461 = n6326 | n6459;
  assign n6462 = ~n6460 & n6461;
  assign n6463 = x54 & x98;
  assign n6464 = n6462 & n6463;
  assign n6465 = n6462 | n6463;
  assign n6466 = ~n6464 & n6465;
  assign n6467 = n6325 & n6466;
  assign n6468 = n6325 | n6466;
  assign n6469 = ~n6467 & n6468;
  assign n6470 = x53 & x99;
  assign n6471 = n6469 & n6470;
  assign n6472 = n6469 | n6470;
  assign n6473 = ~n6471 & n6472;
  assign n6474 = n6324 & n6473;
  assign n6475 = n6324 | n6473;
  assign n6476 = ~n6474 & n6475;
  assign n6477 = x52 & x100;
  assign n6478 = n6476 & n6477;
  assign n6479 = n6476 | n6477;
  assign n6480 = ~n6478 & n6479;
  assign n6481 = n6323 & n6480;
  assign n6482 = n6323 | n6480;
  assign n6483 = ~n6481 & n6482;
  assign n6484 = x51 & x101;
  assign n6485 = n6483 & n6484;
  assign n6486 = n6483 | n6484;
  assign n6487 = ~n6485 & n6486;
  assign n6488 = n16064 & n6487;
  assign n6489 = n16064 | n6487;
  assign n6490 = ~n6488 & n6489;
  assign n6491 = x50 & x102;
  assign n6492 = n6490 & n6491;
  assign n6493 = n6490 | n6491;
  assign n6494 = ~n6492 & n6493;
  assign n6495 = n12835 & n6494;
  assign n6496 = n12835 | n6494;
  assign n6497 = ~n6495 & n6496;
  assign n6498 = x49 & x103;
  assign n6499 = n6497 & n6498;
  assign n6500 = n6497 | n6498;
  assign n6501 = ~n6499 & n6500;
  assign n6502 = n6318 & n6501;
  assign n6503 = n6318 | n6501;
  assign n6504 = ~n6502 & n6503;
  assign n6505 = x48 & x104;
  assign n6506 = n6504 & n6505;
  assign n6507 = n6504 | n6505;
  assign n6508 = ~n6506 & n6507;
  assign n17712 = n6317 | n6498;
  assign n17713 = (n6316 & n6498) | (n6316 & n17712) | (n6498 & n17712);
  assign n16116 = (n6318 & n6497) | (n6318 & n17713) | (n6497 & n17713);
  assign n12912 = (n6499 & n6501) | (n6499 & n16116) | (n6501 & n16116);
  assign n12913 = n6492 | n12835;
  assign n12914 = (n6492 & n6494) | (n6492 & n12913) | (n6494 & n12913);
  assign n16117 = n6485 | n16064;
  assign n16118 = (n6485 & n6487) | (n6485 & n16117) | (n6487 & n16117);
  assign n6512 = n6478 | n6481;
  assign n6513 = n6471 | n6474;
  assign n6514 = n6464 | n6467;
  assign n12915 = n6457 | n6459;
  assign n12916 = (n6326 & n6457) | (n6326 & n12915) | (n6457 & n12915);
  assign n12917 = n6450 | n6452;
  assign n12918 = (n6450 & n12837) | (n6450 & n12917) | (n12837 & n12917);
  assign n12919 = n6443 | n6445;
  assign n12920 = (n6443 & n12839) | (n6443 & n12919) | (n12839 & n12919);
  assign n12921 = n6436 | n6438;
  assign n12922 = (n6436 & n12841) | (n6436 & n12921) | (n12841 & n12921);
  assign n12923 = n6429 | n6431;
  assign n12924 = (n6429 & n12843) | (n6429 & n12923) | (n12843 & n12923);
  assign n12925 = n6422 | n6424;
  assign n12926 = (n6422 & n12845) | (n6422 & n12925) | (n12845 & n12925);
  assign n12927 = n6415 | n6417;
  assign n12928 = (n6415 & n12847) | (n6415 & n12927) | (n12847 & n12927);
  assign n12932 = n6401 | n6403;
  assign n16119 = n6220 | n6401;
  assign n16120 = (n6401 & n6403) | (n6401 & n16119) | (n6403 & n16119);
  assign n16121 = (n12830 & n12932) | (n12830 & n16120) | (n12932 & n16120);
  assign n16122 = (n6222 & n12932) | (n6222 & n16120) | (n12932 & n16120);
  assign n16123 = (n12762 & n16121) | (n12762 & n16122) | (n16121 & n16122);
  assign n12937 = n6380 | n6382;
  assign n16124 = n6199 | n6380;
  assign n16125 = (n6380 & n6382) | (n6380 & n16124) | (n6382 & n16124);
  assign n16126 = (n12821 & n12937) | (n12821 & n16125) | (n12937 & n16125);
  assign n16127 = (n12820 & n12937) | (n12820 & n16125) | (n12937 & n16125);
  assign n16128 = (n15976 & n16126) | (n15976 & n16127) | (n16126 & n16127);
  assign n12799 = (n15955 & n16022) | (n15955 & n16024) | (n16022 & n16024);
  assign n12945 = n6345 | n16074;
  assign n12946 = n6345 | n16076;
  assign n16131 = (n12945 & n12946) | (n12945 & n15925) | (n12946 & n15925);
  assign n16132 = (n12945 & n12946) | (n12945 & n15923) | (n12946 & n15923);
  assign n16133 = (n15804 & n16131) | (n15804 & n16132) | (n16131 & n16132);
  assign n6532 = x73 & x80;
  assign n6533 = x72 & x81;
  assign n6534 = n6532 & n6533;
  assign n6535 = n6532 | n6533;
  assign n6536 = ~n6534 & n6535;
  assign n6537 = n16133 & n6536;
  assign n6538 = n16133 | n6536;
  assign n6539 = ~n6537 & n6538;
  assign n6540 = x71 & x82;
  assign n6541 = n6539 & n6540;
  assign n6542 = n6539 | n6540;
  assign n6543 = ~n6541 & n6542;
  assign n16134 = n6352 | n6354;
  assign n16135 = (n6352 & n12862) | (n6352 & n16134) | (n12862 & n16134);
  assign n12948 = n6543 & n16135;
  assign n16136 = n6171 | n6352;
  assign n16137 = (n6352 & n6354) | (n6352 & n16136) | (n6354 & n16136);
  assign n12949 = n6543 & n16137;
  assign n16138 = (n12948 & n12949) | (n12948 & n16027) | (n12949 & n16027);
  assign n16139 = (n12948 & n12949) | (n12948 & n16026) | (n12949 & n16026);
  assign n16140 = (n15918 & n16138) | (n15918 & n16139) | (n16138 & n16139);
  assign n12951 = n6543 | n16135;
  assign n12952 = n6543 | n16137;
  assign n16141 = (n12951 & n12952) | (n12951 & n16027) | (n12952 & n16027);
  assign n16142 = (n12951 & n12952) | (n12951 & n16026) | (n12952 & n16026);
  assign n16143 = (n15918 & n16141) | (n15918 & n16142) | (n16141 & n16142);
  assign n6546 = ~n16140 & n16143;
  assign n6547 = x70 & x83;
  assign n6548 = n6546 & n6547;
  assign n6549 = n6546 | n6547;
  assign n6550 = ~n6548 & n6549;
  assign n12954 = n6359 & n6550;
  assign n17714 = (n6361 & n6550) | (n6361 & n12954) | (n6550 & n12954);
  assign n17715 = n6550 & n12954;
  assign n17716 = (n16094 & n17714) | (n16094 & n17715) | (n17714 & n17715);
  assign n16145 = (n6550 & n12880) | (n6550 & n12954) | (n12880 & n12954);
  assign n16146 = (n12722 & n17716) | (n12722 & n16145) | (n17716 & n16145);
  assign n12956 = n6359 | n6550;
  assign n17717 = n6361 | n12956;
  assign n17718 = (n12956 & n16094) | (n12956 & n17717) | (n16094 & n17717);
  assign n16148 = n12880 | n12956;
  assign n16149 = (n12722 & n17718) | (n12722 & n16148) | (n17718 & n16148);
  assign n6553 = ~n16146 & n16149;
  assign n6554 = x69 & x84;
  assign n6555 = n6553 & n6554;
  assign n6556 = n6553 | n6554;
  assign n6557 = ~n6555 & n6556;
  assign n17719 = n6366 & n6557;
  assign n17720 = (n6557 & n12885) | (n6557 & n17719) | (n12885 & n17719);
  assign n16129 = n6185 | n6366;
  assign n16130 = (n6366 & n6368) | (n6366 & n16129) | (n6368 & n16129);
  assign n16151 = n6557 & n16130;
  assign n16152 = (n12799 & n17720) | (n12799 & n16151) | (n17720 & n16151);
  assign n17721 = n6366 | n6557;
  assign n17722 = n12885 | n17721;
  assign n16154 = n6557 | n16130;
  assign n16155 = (n12799 & n17722) | (n12799 & n16154) | (n17722 & n16154);
  assign n6560 = ~n16152 & n16155;
  assign n6561 = x68 & x85;
  assign n6562 = n6560 & n6561;
  assign n6563 = n6560 | n6561;
  assign n6564 = ~n6562 & n6563;
  assign n12958 = n6373 & n6564;
  assign n16156 = (n6564 & n12891) | (n6564 & n12958) | (n12891 & n12958);
  assign n16157 = (n6564 & n12892) | (n6564 & n12958) | (n12892 & n12958);
  assign n16158 = (n16020 & n16156) | (n16020 & n16157) | (n16156 & n16157);
  assign n12960 = n6373 | n6564;
  assign n16159 = n12891 | n12960;
  assign n16160 = n12892 | n12960;
  assign n16161 = (n16020 & n16159) | (n16020 & n16160) | (n16159 & n16160);
  assign n6567 = ~n16158 & n16161;
  assign n6568 = x67 & x86;
  assign n6569 = n6567 & n6568;
  assign n6570 = n6567 | n6568;
  assign n6571 = ~n6569 & n6570;
  assign n6572 = n16128 & n6571;
  assign n6573 = n16128 | n6571;
  assign n6574 = ~n6572 & n6573;
  assign n6575 = x66 & x87;
  assign n6576 = n6574 & n6575;
  assign n6577 = n6574 | n6575;
  assign n6578 = ~n6576 & n6577;
  assign n12934 = n6387 | n6389;
  assign n12962 = n6578 & n12934;
  assign n12963 = n6387 & n6578;
  assign n12964 = (n16069 & n12962) | (n16069 & n12963) | (n12962 & n12963);
  assign n12965 = n6578 | n12934;
  assign n12966 = n6387 | n6578;
  assign n12967 = (n16069 & n12965) | (n16069 & n12966) | (n12965 & n12966);
  assign n6581 = ~n12964 & n12967;
  assign n6582 = x65 & x88;
  assign n6583 = n6581 & n6582;
  assign n6584 = n6581 | n6582;
  assign n6585 = ~n6583 & n6584;
  assign n12968 = n6394 & n6585;
  assign n16162 = (n6585 & n12902) | (n6585 & n12968) | (n12902 & n12968);
  assign n16163 = (n6585 & n12901) | (n6585 & n12968) | (n12901 & n12968);
  assign n16164 = (n16015 & n16162) | (n16015 & n16163) | (n16162 & n16163);
  assign n12970 = n6394 | n6585;
  assign n16165 = n12902 | n12970;
  assign n16166 = n12901 | n12970;
  assign n16167 = (n16015 & n16165) | (n16015 & n16166) | (n16165 & n16166);
  assign n6588 = ~n16164 & n16167;
  assign n6589 = x64 & x89;
  assign n6590 = n6588 & n6589;
  assign n6591 = n6588 | n6589;
  assign n6592 = ~n6590 & n6591;
  assign n6593 = n16123 & n6592;
  assign n6594 = n16123 | n6592;
  assign n6595 = ~n6593 & n6594;
  assign n6596 = x63 & x90;
  assign n6597 = n6595 & n6596;
  assign n6598 = n6595 | n6596;
  assign n6599 = ~n6597 & n6598;
  assign n12929 = n6408 | n6410;
  assign n16168 = n6599 & n12929;
  assign n16169 = n6408 & n6599;
  assign n16170 = (n12849 & n16168) | (n12849 & n16169) | (n16168 & n16169);
  assign n16171 = n6599 | n12929;
  assign n16172 = n6408 | n6599;
  assign n16173 = (n12849 & n16171) | (n12849 & n16172) | (n16171 & n16172);
  assign n6602 = ~n16170 & n16173;
  assign n6603 = x62 & x91;
  assign n6604 = n6602 & n6603;
  assign n6605 = n6602 | n6603;
  assign n6606 = ~n6604 & n6605;
  assign n6607 = n12928 & n6606;
  assign n6608 = n12928 | n6606;
  assign n6609 = ~n6607 & n6608;
  assign n6610 = x61 & x92;
  assign n6611 = n6609 & n6610;
  assign n6612 = n6609 | n6610;
  assign n6613 = ~n6611 & n6612;
  assign n6614 = n12926 & n6613;
  assign n6615 = n12926 | n6613;
  assign n6616 = ~n6614 & n6615;
  assign n6617 = x60 & x93;
  assign n6618 = n6616 & n6617;
  assign n6619 = n6616 | n6617;
  assign n6620 = ~n6618 & n6619;
  assign n6621 = n12924 & n6620;
  assign n6622 = n12924 | n6620;
  assign n6623 = ~n6621 & n6622;
  assign n6624 = x59 & x94;
  assign n6625 = n6623 & n6624;
  assign n6626 = n6623 | n6624;
  assign n6627 = ~n6625 & n6626;
  assign n6628 = n12922 & n6627;
  assign n6629 = n12922 | n6627;
  assign n6630 = ~n6628 & n6629;
  assign n6631 = x58 & x95;
  assign n6632 = n6630 & n6631;
  assign n6633 = n6630 | n6631;
  assign n6634 = ~n6632 & n6633;
  assign n6635 = n12920 & n6634;
  assign n6636 = n12920 | n6634;
  assign n6637 = ~n6635 & n6636;
  assign n6638 = x57 & x96;
  assign n6639 = n6637 & n6638;
  assign n6640 = n6637 | n6638;
  assign n6641 = ~n6639 & n6640;
  assign n6642 = n12918 & n6641;
  assign n6643 = n12918 | n6641;
  assign n6644 = ~n6642 & n6643;
  assign n6645 = x56 & x97;
  assign n6646 = n6644 & n6645;
  assign n6647 = n6644 | n6645;
  assign n6648 = ~n6646 & n6647;
  assign n6649 = n12916 & n6648;
  assign n6650 = n12916 | n6648;
  assign n6651 = ~n6649 & n6650;
  assign n6652 = x55 & x98;
  assign n6653 = n6651 & n6652;
  assign n6654 = n6651 | n6652;
  assign n6655 = ~n6653 & n6654;
  assign n6656 = n6514 & n6655;
  assign n6657 = n6514 | n6655;
  assign n6658 = ~n6656 & n6657;
  assign n6659 = x54 & x99;
  assign n6660 = n6658 & n6659;
  assign n6661 = n6658 | n6659;
  assign n6662 = ~n6660 & n6661;
  assign n6663 = n6513 & n6662;
  assign n6664 = n6513 | n6662;
  assign n6665 = ~n6663 & n6664;
  assign n6666 = x53 & x100;
  assign n6667 = n6665 & n6666;
  assign n6668 = n6665 | n6666;
  assign n6669 = ~n6667 & n6668;
  assign n6670 = n6512 & n6669;
  assign n6671 = n6512 | n6669;
  assign n6672 = ~n6670 & n6671;
  assign n6673 = x52 & x101;
  assign n6674 = n6672 & n6673;
  assign n6675 = n6672 | n6673;
  assign n6676 = ~n6674 & n6675;
  assign n6677 = n16118 & n6676;
  assign n6678 = n16118 | n6676;
  assign n6679 = ~n6677 & n6678;
  assign n6680 = x51 & x102;
  assign n6681 = n6679 & n6680;
  assign n6682 = n6679 | n6680;
  assign n6683 = ~n6681 & n6682;
  assign n6684 = n12914 & n6683;
  assign n6685 = n12914 | n6683;
  assign n6686 = ~n6684 & n6685;
  assign n6687 = x50 & x103;
  assign n6688 = n6686 & n6687;
  assign n6689 = n6686 | n6687;
  assign n6690 = ~n6688 & n6689;
  assign n6691 = n12912 & n6690;
  assign n6692 = n12912 | n6690;
  assign n6693 = ~n6691 & n6692;
  assign n6694 = x49 & x104;
  assign n6695 = n6693 & n6694;
  assign n6696 = n6693 | n6694;
  assign n6697 = ~n6695 & n6696;
  assign n6698 = n6506 & n6697;
  assign n6699 = n6506 | n6697;
  assign n6700 = ~n6698 & n6699;
  assign n6701 = x48 & x105;
  assign n6702 = n6700 & n6701;
  assign n6703 = n6700 | n6701;
  assign n6704 = ~n6702 & n6703;
  assign n17723 = n6505 | n6694;
  assign n17724 = (n6504 & n6694) | (n6504 & n17723) | (n6694 & n17723);
  assign n16175 = (n6506 & n6693) | (n6506 & n17724) | (n6693 & n17724);
  assign n12973 = (n6695 & n6697) | (n6695 & n16175) | (n6697 & n16175);
  assign n12974 = n6688 | n12912;
  assign n12975 = (n6688 & n6690) | (n6688 & n12974) | (n6690 & n12974);
  assign n12976 = n6681 | n12914;
  assign n12977 = (n6681 & n6683) | (n6681 & n12976) | (n6683 & n12976);
  assign n16176 = n6674 | n16118;
  assign n16177 = (n6674 & n6676) | (n6674 & n16176) | (n6676 & n16176);
  assign n6709 = n6667 | n6670;
  assign n6710 = n6660 | n6663;
  assign n12978 = n6653 | n6655;
  assign n12979 = (n6514 & n6653) | (n6514 & n12978) | (n6653 & n12978);
  assign n12980 = n6646 | n6648;
  assign n12981 = (n6646 & n12916) | (n6646 & n12980) | (n12916 & n12980);
  assign n12982 = n6639 | n6641;
  assign n12983 = (n6639 & n12918) | (n6639 & n12982) | (n12918 & n12982);
  assign n12984 = n6632 | n6634;
  assign n12985 = (n6632 & n12920) | (n6632 & n12984) | (n12920 & n12984);
  assign n12986 = n6625 | n6627;
  assign n12987 = (n6625 & n12922) | (n6625 & n12986) | (n12922 & n12986);
  assign n12988 = n6618 | n6620;
  assign n12989 = (n6618 & n12924) | (n6618 & n12988) | (n12924 & n12988);
  assign n12990 = n6611 | n6613;
  assign n12991 = (n6611 & n12926) | (n6611 & n12990) | (n12926 & n12990);
  assign n12930 = (n6408 & n12849) | (n6408 & n12929) | (n12849 & n12929);
  assign n12999 = n6583 | n6585;
  assign n16178 = n6394 | n6583;
  assign n16179 = (n6583 & n6585) | (n6583 & n16178) | (n6585 & n16178);
  assign n16180 = (n12902 & n12999) | (n12902 & n16179) | (n12999 & n16179);
  assign n16181 = (n12901 & n12999) | (n12901 & n16179) | (n12999 & n16179);
  assign n16182 = (n16015 & n16180) | (n16015 & n16181) | (n16180 & n16181);
  assign n13004 = n6562 | n6564;
  assign n16183 = n6373 | n6562;
  assign n16184 = (n6562 & n6564) | (n6562 & n16183) | (n6564 & n16183);
  assign n16185 = (n12891 & n13004) | (n12891 & n16184) | (n13004 & n16184);
  assign n16186 = (n12892 & n13004) | (n12892 & n16184) | (n13004 & n16184);
  assign n16187 = (n16020 & n16185) | (n16020 & n16186) | (n16185 & n16186);
  assign n12939 = n6366 | n12885;
  assign n13012 = n6541 | n12949;
  assign n16188 = n6541 | n6543;
  assign n16189 = (n6541 & n16135) | (n6541 & n16188) | (n16135 & n16188);
  assign n16190 = (n13012 & n16027) | (n13012 & n16189) | (n16027 & n16189);
  assign n16191 = (n13012 & n16026) | (n13012 & n16189) | (n16026 & n16189);
  assign n16192 = (n15918 & n16190) | (n15918 & n16191) | (n16190 & n16191);
  assign n6729 = x74 & x80;
  assign n6730 = x73 & x81;
  assign n6731 = n6729 & n6730;
  assign n6732 = n6729 | n6730;
  assign n6733 = ~n6731 & n6732;
  assign n13014 = n6534 | n6536;
  assign n13016 = n6733 & n13014;
  assign n13017 = n6534 & n6733;
  assign n13018 = (n16133 & n13016) | (n16133 & n13017) | (n13016 & n13017);
  assign n13019 = n6733 | n13014;
  assign n13020 = n6534 | n6733;
  assign n13021 = (n16133 & n13019) | (n16133 & n13020) | (n13019 & n13020);
  assign n6736 = ~n13018 & n13021;
  assign n6737 = x72 & x82;
  assign n6738 = n6736 & n6737;
  assign n6739 = n6736 | n6737;
  assign n6740 = ~n6738 & n6739;
  assign n6741 = n16192 & n6740;
  assign n6742 = n16192 | n6740;
  assign n6743 = ~n6741 & n6742;
  assign n6744 = x71 & x83;
  assign n6745 = n6743 & n6744;
  assign n6746 = n6743 | n6744;
  assign n6747 = ~n6745 & n6746;
  assign n16193 = n6359 | n6548;
  assign n16194 = (n6548 & n6550) | (n6548 & n16193) | (n6550 & n16193);
  assign n13022 = n6747 & n16194;
  assign n13009 = n6548 | n6550;
  assign n13023 = n6747 & n13009;
  assign n16195 = (n12879 & n13022) | (n12879 & n13023) | (n13022 & n13023);
  assign n16196 = (n12880 & n13022) | (n12880 & n13023) | (n13022 & n13023);
  assign n16197 = (n12722 & n16195) | (n12722 & n16196) | (n16195 & n16196);
  assign n13025 = n6747 | n16194;
  assign n13026 = n6747 | n13009;
  assign n16198 = (n12879 & n13025) | (n12879 & n13026) | (n13025 & n13026);
  assign n16199 = (n12880 & n13025) | (n12880 & n13026) | (n13025 & n13026);
  assign n16200 = (n12722 & n16198) | (n12722 & n16199) | (n16198 & n16199);
  assign n6750 = ~n16197 & n16200;
  assign n6751 = x70 & x84;
  assign n6752 = n6750 & n6751;
  assign n6753 = n6750 | n6751;
  assign n6754 = ~n6752 & n6753;
  assign n13006 = n6555 | n6557;
  assign n13028 = n6754 & n13006;
  assign n13029 = n6555 & n6754;
  assign n16201 = (n12939 & n13028) | (n12939 & n13029) | (n13028 & n13029);
  assign n16202 = (n13028 & n13029) | (n13028 & n16130) | (n13029 & n16130);
  assign n16203 = (n12799 & n16201) | (n12799 & n16202) | (n16201 & n16202);
  assign n13031 = n6754 | n13006;
  assign n13032 = n6555 | n6754;
  assign n16204 = (n12939 & n13031) | (n12939 & n13032) | (n13031 & n13032);
  assign n16205 = (n13031 & n13032) | (n13031 & n16130) | (n13032 & n16130);
  assign n16206 = (n12799 & n16204) | (n12799 & n16205) | (n16204 & n16205);
  assign n6757 = ~n16203 & n16206;
  assign n6758 = x69 & x85;
  assign n6759 = n6757 & n6758;
  assign n6760 = n6757 | n6758;
  assign n6761 = ~n6759 & n6760;
  assign n6762 = n16187 & n6761;
  assign n6763 = n16187 | n6761;
  assign n6764 = ~n6762 & n6763;
  assign n6765 = x68 & x86;
  assign n6766 = n6764 & n6765;
  assign n6767 = n6764 | n6765;
  assign n6768 = ~n6766 & n6767;
  assign n13001 = n6569 | n6571;
  assign n13034 = n6768 & n13001;
  assign n13035 = n6569 & n6768;
  assign n13036 = (n16128 & n13034) | (n16128 & n13035) | (n13034 & n13035);
  assign n13037 = n6768 | n13001;
  assign n13038 = n6569 | n6768;
  assign n13039 = (n16128 & n13037) | (n16128 & n13038) | (n13037 & n13038);
  assign n6771 = ~n13036 & n13039;
  assign n6772 = x67 & x87;
  assign n6773 = n6771 & n6772;
  assign n6774 = n6771 | n6772;
  assign n6775 = ~n6773 & n6774;
  assign n13040 = n6576 & n6775;
  assign n16207 = (n6775 & n12963) | (n6775 & n13040) | (n12963 & n13040);
  assign n16208 = (n6775 & n12962) | (n6775 & n13040) | (n12962 & n13040);
  assign n16209 = (n16069 & n16207) | (n16069 & n16208) | (n16207 & n16208);
  assign n13042 = n6576 | n6775;
  assign n16210 = n12963 | n13042;
  assign n16211 = n12962 | n13042;
  assign n16212 = (n16069 & n16210) | (n16069 & n16211) | (n16210 & n16211);
  assign n6778 = ~n16209 & n16212;
  assign n6779 = x66 & x88;
  assign n6780 = n6778 & n6779;
  assign n6781 = n6778 | n6779;
  assign n6782 = ~n6780 & n6781;
  assign n6783 = n16182 & n6782;
  assign n6784 = n16182 | n6782;
  assign n6785 = ~n6783 & n6784;
  assign n6786 = x65 & x89;
  assign n6787 = n6785 & n6786;
  assign n6788 = n6785 | n6786;
  assign n6789 = ~n6787 & n6788;
  assign n12996 = n6590 | n6592;
  assign n13044 = n6789 & n12996;
  assign n13045 = n6590 & n6789;
  assign n13046 = (n16123 & n13044) | (n16123 & n13045) | (n13044 & n13045);
  assign n13047 = n6789 | n12996;
  assign n13048 = n6590 | n6789;
  assign n13049 = (n16123 & n13047) | (n16123 & n13048) | (n13047 & n13048);
  assign n6792 = ~n13046 & n13049;
  assign n6793 = x64 & x90;
  assign n6794 = n6792 & n6793;
  assign n6795 = n6792 | n6793;
  assign n6796 = ~n6794 & n6795;
  assign n12994 = n6597 | n6599;
  assign n16213 = n6796 & n12994;
  assign n16214 = n6597 & n6796;
  assign n16215 = (n12930 & n16213) | (n12930 & n16214) | (n16213 & n16214);
  assign n16216 = n6796 | n12994;
  assign n16217 = n6597 | n6796;
  assign n16218 = (n12930 & n16216) | (n12930 & n16217) | (n16216 & n16217);
  assign n6799 = ~n16215 & n16218;
  assign n6800 = x63 & x91;
  assign n6801 = n6799 & n6800;
  assign n6802 = n6799 | n6800;
  assign n6803 = ~n6801 & n6802;
  assign n12992 = n6604 | n6606;
  assign n16219 = n6803 & n12992;
  assign n16220 = n6604 & n6803;
  assign n16221 = (n12928 & n16219) | (n12928 & n16220) | (n16219 & n16220);
  assign n16222 = n6803 | n12992;
  assign n16223 = n6604 | n6803;
  assign n16224 = (n12928 & n16222) | (n12928 & n16223) | (n16222 & n16223);
  assign n6806 = ~n16221 & n16224;
  assign n6807 = x62 & x92;
  assign n6808 = n6806 & n6807;
  assign n6809 = n6806 | n6807;
  assign n6810 = ~n6808 & n6809;
  assign n6811 = n12991 & n6810;
  assign n6812 = n12991 | n6810;
  assign n6813 = ~n6811 & n6812;
  assign n6814 = x61 & x93;
  assign n6815 = n6813 & n6814;
  assign n6816 = n6813 | n6814;
  assign n6817 = ~n6815 & n6816;
  assign n6818 = n12989 & n6817;
  assign n6819 = n12989 | n6817;
  assign n6820 = ~n6818 & n6819;
  assign n6821 = x60 & x94;
  assign n6822 = n6820 & n6821;
  assign n6823 = n6820 | n6821;
  assign n6824 = ~n6822 & n6823;
  assign n6825 = n12987 & n6824;
  assign n6826 = n12987 | n6824;
  assign n6827 = ~n6825 & n6826;
  assign n6828 = x59 & x95;
  assign n6829 = n6827 & n6828;
  assign n6830 = n6827 | n6828;
  assign n6831 = ~n6829 & n6830;
  assign n6832 = n12985 & n6831;
  assign n6833 = n12985 | n6831;
  assign n6834 = ~n6832 & n6833;
  assign n6835 = x58 & x96;
  assign n6836 = n6834 & n6835;
  assign n6837 = n6834 | n6835;
  assign n6838 = ~n6836 & n6837;
  assign n6839 = n12983 & n6838;
  assign n6840 = n12983 | n6838;
  assign n6841 = ~n6839 & n6840;
  assign n6842 = x57 & x97;
  assign n6843 = n6841 & n6842;
  assign n6844 = n6841 | n6842;
  assign n6845 = ~n6843 & n6844;
  assign n6846 = n12981 & n6845;
  assign n6847 = n12981 | n6845;
  assign n6848 = ~n6846 & n6847;
  assign n6849 = x56 & x98;
  assign n6850 = n6848 & n6849;
  assign n6851 = n6848 | n6849;
  assign n6852 = ~n6850 & n6851;
  assign n6853 = n12979 & n6852;
  assign n6854 = n12979 | n6852;
  assign n6855 = ~n6853 & n6854;
  assign n6856 = x55 & x99;
  assign n6857 = n6855 & n6856;
  assign n6858 = n6855 | n6856;
  assign n6859 = ~n6857 & n6858;
  assign n6860 = n6710 & n6859;
  assign n6861 = n6710 | n6859;
  assign n6862 = ~n6860 & n6861;
  assign n6863 = x54 & x100;
  assign n6864 = n6862 & n6863;
  assign n6865 = n6862 | n6863;
  assign n6866 = ~n6864 & n6865;
  assign n6867 = n6709 & n6866;
  assign n6868 = n6709 | n6866;
  assign n6869 = ~n6867 & n6868;
  assign n6870 = x53 & x101;
  assign n6871 = n6869 & n6870;
  assign n6872 = n6869 | n6870;
  assign n6873 = ~n6871 & n6872;
  assign n6874 = n16177 & n6873;
  assign n6875 = n16177 | n6873;
  assign n6876 = ~n6874 & n6875;
  assign n6877 = x52 & x102;
  assign n6878 = n6876 & n6877;
  assign n6879 = n6876 | n6877;
  assign n6880 = ~n6878 & n6879;
  assign n6881 = n12977 & n6880;
  assign n6882 = n12977 | n6880;
  assign n6883 = ~n6881 & n6882;
  assign n6884 = x51 & x103;
  assign n6885 = n6883 & n6884;
  assign n6886 = n6883 | n6884;
  assign n6887 = ~n6885 & n6886;
  assign n6888 = n12975 & n6887;
  assign n6889 = n12975 | n6887;
  assign n6890 = ~n6888 & n6889;
  assign n6891 = x50 & x104;
  assign n6892 = n6890 & n6891;
  assign n6893 = n6890 | n6891;
  assign n6894 = ~n6892 & n6893;
  assign n6895 = n12973 & n6894;
  assign n6896 = n12973 | n6894;
  assign n6897 = ~n6895 & n6896;
  assign n6898 = x49 & x105;
  assign n6899 = n6897 & n6898;
  assign n6900 = n6897 | n6898;
  assign n6901 = ~n6899 & n6900;
  assign n6902 = n6702 & n6901;
  assign n6903 = n6702 | n6901;
  assign n6904 = ~n6902 & n6903;
  assign n6905 = x48 & x106;
  assign n6906 = n6904 & n6905;
  assign n6907 = n6904 | n6905;
  assign n6908 = ~n6906 & n6907;
  assign n17725 = n6701 | n6898;
  assign n17726 = (n6700 & n6898) | (n6700 & n17725) | (n6898 & n17725);
  assign n16226 = (n6702 & n6897) | (n6702 & n17726) | (n6897 & n17726);
  assign n13051 = (n6899 & n6901) | (n6899 & n16226) | (n6901 & n16226);
  assign n13052 = n6892 | n12973;
  assign n13053 = (n6892 & n6894) | (n6892 & n13052) | (n6894 & n13052);
  assign n13054 = n6885 | n12975;
  assign n13055 = (n6885 & n6887) | (n6885 & n13054) | (n6887 & n13054);
  assign n13056 = n6878 | n12977;
  assign n13057 = (n6878 & n6880) | (n6878 & n13056) | (n6880 & n13056);
  assign n16227 = n6871 | n16177;
  assign n16228 = (n6871 & n6873) | (n6871 & n16227) | (n6873 & n16227);
  assign n6914 = n6864 | n6867;
  assign n13058 = n6857 | n6859;
  assign n13059 = (n6710 & n6857) | (n6710 & n13058) | (n6857 & n13058);
  assign n13060 = n6850 | n6852;
  assign n13061 = (n6850 & n12979) | (n6850 & n13060) | (n12979 & n13060);
  assign n13062 = n6843 | n6845;
  assign n13063 = (n6843 & n12981) | (n6843 & n13062) | (n12981 & n13062);
  assign n13064 = n6836 | n6838;
  assign n13065 = (n6836 & n12983) | (n6836 & n13064) | (n12983 & n13064);
  assign n13066 = n6829 | n6831;
  assign n13067 = (n6829 & n12985) | (n6829 & n13066) | (n12985 & n13066);
  assign n13068 = n6822 | n6824;
  assign n13069 = (n6822 & n12987) | (n6822 & n13068) | (n12987 & n13068);
  assign n13070 = n6815 | n6817;
  assign n13071 = (n6815 & n12989) | (n6815 & n13070) | (n12989 & n13070);
  assign n12993 = (n6604 & n12928) | (n6604 & n12992) | (n12928 & n12992);
  assign n12995 = (n6597 & n12930) | (n6597 & n12994) | (n12930 & n12994);
  assign n13081 = n6773 | n6775;
  assign n16229 = n6576 | n6773;
  assign n16230 = (n6773 & n6775) | (n6773 & n16229) | (n6775 & n16229);
  assign n16231 = (n12963 & n13081) | (n12963 & n16230) | (n13081 & n16230);
  assign n16232 = (n12962 & n13081) | (n12962 & n16230) | (n13081 & n16230);
  assign n16233 = (n16069 & n16231) | (n16069 & n16232) | (n16231 & n16232);
  assign n16234 = n6752 | n6754;
  assign n16235 = (n6752 & n13006) | (n6752 & n16234) | (n13006 & n16234);
  assign n16236 = n6555 | n6752;
  assign n16237 = (n6752 & n6754) | (n6752 & n16236) | (n6754 & n16236);
  assign n16238 = (n12939 & n16235) | (n12939 & n16237) | (n16235 & n16237);
  assign n16239 = (n16130 & n16235) | (n16130 & n16237) | (n16235 & n16237);
  assign n16240 = (n12799 & n16238) | (n12799 & n16239) | (n16238 & n16239);
  assign n13088 = n6745 | n13022;
  assign n13089 = n6745 | n13023;
  assign n16241 = (n12879 & n13088) | (n12879 & n13089) | (n13088 & n13089);
  assign n16242 = (n12880 & n13088) | (n12880 & n13089) | (n13088 & n13089);
  assign n16243 = (n12722 & n16241) | (n12722 & n16242) | (n16241 & n16242);
  assign n6934 = x75 & x80;
  assign n6935 = x74 & x81;
  assign n6936 = n6934 & n6935;
  assign n6937 = n6934 | n6935;
  assign n6938 = ~n6936 & n6937;
  assign n16244 = n6731 | n6733;
  assign n16245 = (n6731 & n13014) | (n6731 & n16244) | (n13014 & n16244);
  assign n13096 = n6938 & n16245;
  assign n16246 = n6534 | n6731;
  assign n16247 = (n6731 & n6733) | (n6731 & n16246) | (n6733 & n16246);
  assign n13097 = n6938 & n16247;
  assign n13098 = (n16133 & n13096) | (n16133 & n13097) | (n13096 & n13097);
  assign n13099 = n6938 | n16245;
  assign n13100 = n6938 | n16247;
  assign n13101 = (n16133 & n13099) | (n16133 & n13100) | (n13099 & n13100);
  assign n6941 = ~n13098 & n13101;
  assign n6942 = x73 & x82;
  assign n6943 = n6941 & n6942;
  assign n6944 = n6941 | n6942;
  assign n6945 = ~n6943 & n6944;
  assign n13091 = n6738 | n6740;
  assign n13102 = n6945 & n13091;
  assign n13103 = n6738 & n6945;
  assign n13104 = (n16192 & n13102) | (n16192 & n13103) | (n13102 & n13103);
  assign n13105 = n6945 | n13091;
  assign n13106 = n6738 | n6945;
  assign n13107 = (n16192 & n13105) | (n16192 & n13106) | (n13105 & n13106);
  assign n6948 = ~n13104 & n13107;
  assign n6949 = x72 & x83;
  assign n6950 = n6948 & n6949;
  assign n6951 = n6948 | n6949;
  assign n6952 = ~n6950 & n6951;
  assign n6953 = n16243 & n6952;
  assign n6954 = n16243 | n6952;
  assign n6955 = ~n6953 & n6954;
  assign n6956 = x71 & x84;
  assign n6957 = n6955 & n6956;
  assign n6958 = n6955 | n6956;
  assign n6959 = ~n6957 & n6958;
  assign n6960 = n16240 & n6959;
  assign n6961 = n16240 | n6959;
  assign n6962 = ~n6960 & n6961;
  assign n6963 = x70 & x85;
  assign n6964 = n6962 & n6963;
  assign n6965 = n6962 | n6963;
  assign n6966 = ~n6964 & n6965;
  assign n13083 = n6759 | n6761;
  assign n13108 = n6966 & n13083;
  assign n13109 = n6759 & n6966;
  assign n13110 = (n16187 & n13108) | (n16187 & n13109) | (n13108 & n13109);
  assign n13111 = n6966 | n13083;
  assign n13112 = n6759 | n6966;
  assign n13113 = (n16187 & n13111) | (n16187 & n13112) | (n13111 & n13112);
  assign n6969 = ~n13110 & n13113;
  assign n6970 = x69 & x86;
  assign n6971 = n6969 & n6970;
  assign n6972 = n6969 | n6970;
  assign n6973 = ~n6971 & n6972;
  assign n13114 = n6766 & n6973;
  assign n16248 = (n6973 & n13035) | (n6973 & n13114) | (n13035 & n13114);
  assign n16249 = (n6973 & n13034) | (n6973 & n13114) | (n13034 & n13114);
  assign n16250 = (n16128 & n16248) | (n16128 & n16249) | (n16248 & n16249);
  assign n13116 = n6766 | n6973;
  assign n16251 = n13035 | n13116;
  assign n16252 = n13034 | n13116;
  assign n16253 = (n16128 & n16251) | (n16128 & n16252) | (n16251 & n16252);
  assign n6976 = ~n16250 & n16253;
  assign n6977 = x68 & x87;
  assign n6978 = n6976 & n6977;
  assign n6979 = n6976 | n6977;
  assign n6980 = ~n6978 & n6979;
  assign n6981 = n16233 & n6980;
  assign n6982 = n16233 | n6980;
  assign n6983 = ~n6981 & n6982;
  assign n6984 = x67 & x88;
  assign n6985 = n6983 & n6984;
  assign n6986 = n6983 | n6984;
  assign n6987 = ~n6985 & n6986;
  assign n13078 = n6780 | n6782;
  assign n13118 = n6987 & n13078;
  assign n13119 = n6780 & n6987;
  assign n13120 = (n16182 & n13118) | (n16182 & n13119) | (n13118 & n13119);
  assign n13121 = n6987 | n13078;
  assign n13122 = n6780 | n6987;
  assign n13123 = (n16182 & n13121) | (n16182 & n13122) | (n13121 & n13122);
  assign n6990 = ~n13120 & n13123;
  assign n6991 = x66 & x89;
  assign n6992 = n6990 & n6991;
  assign n6993 = n6990 | n6991;
  assign n6994 = ~n6992 & n6993;
  assign n13124 = n6787 & n6994;
  assign n16254 = (n6994 & n13045) | (n6994 & n13124) | (n13045 & n13124);
  assign n16255 = (n6994 & n13044) | (n6994 & n13124) | (n13044 & n13124);
  assign n16256 = (n16123 & n16254) | (n16123 & n16255) | (n16254 & n16255);
  assign n13126 = n6787 | n6994;
  assign n16257 = n13045 | n13126;
  assign n16258 = n13044 | n13126;
  assign n16259 = (n16123 & n16257) | (n16123 & n16258) | (n16257 & n16258);
  assign n6997 = ~n16256 & n16259;
  assign n6998 = x65 & x90;
  assign n6999 = n6997 & n6998;
  assign n7000 = n6997 | n6998;
  assign n7001 = ~n6999 & n7000;
  assign n13076 = n6794 | n6796;
  assign n13128 = n7001 & n13076;
  assign n13129 = n6794 & n7001;
  assign n13130 = (n12995 & n13128) | (n12995 & n13129) | (n13128 & n13129);
  assign n13131 = n7001 | n13076;
  assign n13132 = n6794 | n7001;
  assign n13133 = (n12995 & n13131) | (n12995 & n13132) | (n13131 & n13132);
  assign n7004 = ~n13130 & n13133;
  assign n7005 = x64 & x91;
  assign n7006 = n7004 & n7005;
  assign n7007 = n7004 | n7005;
  assign n7008 = ~n7006 & n7007;
  assign n13074 = n6801 | n6803;
  assign n16260 = n7008 & n13074;
  assign n16261 = n6801 & n7008;
  assign n16262 = (n12993 & n16260) | (n12993 & n16261) | (n16260 & n16261);
  assign n16263 = n7008 | n13074;
  assign n16264 = n6801 | n7008;
  assign n16265 = (n12993 & n16263) | (n12993 & n16264) | (n16263 & n16264);
  assign n7011 = ~n16262 & n16265;
  assign n7012 = x63 & x92;
  assign n7013 = n7011 & n7012;
  assign n7014 = n7011 | n7012;
  assign n7015 = ~n7013 & n7014;
  assign n13072 = n6808 | n6810;
  assign n16266 = n7015 & n13072;
  assign n16267 = n6808 & n7015;
  assign n16268 = (n12991 & n16266) | (n12991 & n16267) | (n16266 & n16267);
  assign n16269 = n7015 | n13072;
  assign n16270 = n6808 | n7015;
  assign n16271 = (n12991 & n16269) | (n12991 & n16270) | (n16269 & n16270);
  assign n7018 = ~n16268 & n16271;
  assign n7019 = x62 & x93;
  assign n7020 = n7018 & n7019;
  assign n7021 = n7018 | n7019;
  assign n7022 = ~n7020 & n7021;
  assign n7023 = n13071 & n7022;
  assign n7024 = n13071 | n7022;
  assign n7025 = ~n7023 & n7024;
  assign n7026 = x61 & x94;
  assign n7027 = n7025 & n7026;
  assign n7028 = n7025 | n7026;
  assign n7029 = ~n7027 & n7028;
  assign n7030 = n13069 & n7029;
  assign n7031 = n13069 | n7029;
  assign n7032 = ~n7030 & n7031;
  assign n7033 = x60 & x95;
  assign n7034 = n7032 & n7033;
  assign n7035 = n7032 | n7033;
  assign n7036 = ~n7034 & n7035;
  assign n7037 = n13067 & n7036;
  assign n7038 = n13067 | n7036;
  assign n7039 = ~n7037 & n7038;
  assign n7040 = x59 & x96;
  assign n7041 = n7039 & n7040;
  assign n7042 = n7039 | n7040;
  assign n7043 = ~n7041 & n7042;
  assign n7044 = n13065 & n7043;
  assign n7045 = n13065 | n7043;
  assign n7046 = ~n7044 & n7045;
  assign n7047 = x58 & x97;
  assign n7048 = n7046 & n7047;
  assign n7049 = n7046 | n7047;
  assign n7050 = ~n7048 & n7049;
  assign n7051 = n13063 & n7050;
  assign n7052 = n13063 | n7050;
  assign n7053 = ~n7051 & n7052;
  assign n7054 = x57 & x98;
  assign n7055 = n7053 & n7054;
  assign n7056 = n7053 | n7054;
  assign n7057 = ~n7055 & n7056;
  assign n7058 = n13061 & n7057;
  assign n7059 = n13061 | n7057;
  assign n7060 = ~n7058 & n7059;
  assign n7061 = x56 & x99;
  assign n7062 = n7060 & n7061;
  assign n7063 = n7060 | n7061;
  assign n7064 = ~n7062 & n7063;
  assign n7065 = n13059 & n7064;
  assign n7066 = n13059 | n7064;
  assign n7067 = ~n7065 & n7066;
  assign n7068 = x55 & x100;
  assign n7069 = n7067 & n7068;
  assign n7070 = n7067 | n7068;
  assign n7071 = ~n7069 & n7070;
  assign n7072 = n6914 & n7071;
  assign n7073 = n6914 | n7071;
  assign n7074 = ~n7072 & n7073;
  assign n7075 = x54 & x101;
  assign n7076 = n7074 & n7075;
  assign n7077 = n7074 | n7075;
  assign n7078 = ~n7076 & n7077;
  assign n7079 = n16228 & n7078;
  assign n7080 = n16228 | n7078;
  assign n7081 = ~n7079 & n7080;
  assign n7082 = x53 & x102;
  assign n7083 = n7081 & n7082;
  assign n7084 = n7081 | n7082;
  assign n7085 = ~n7083 & n7084;
  assign n7086 = n13057 & n7085;
  assign n7087 = n13057 | n7085;
  assign n7088 = ~n7086 & n7087;
  assign n7089 = x52 & x103;
  assign n7090 = n7088 & n7089;
  assign n7091 = n7088 | n7089;
  assign n7092 = ~n7090 & n7091;
  assign n7093 = n13055 & n7092;
  assign n7094 = n13055 | n7092;
  assign n7095 = ~n7093 & n7094;
  assign n7096 = x51 & x104;
  assign n7097 = n7095 & n7096;
  assign n7098 = n7095 | n7096;
  assign n7099 = ~n7097 & n7098;
  assign n7100 = n13053 & n7099;
  assign n7101 = n13053 | n7099;
  assign n7102 = ~n7100 & n7101;
  assign n7103 = x50 & x105;
  assign n7104 = n7102 & n7103;
  assign n7105 = n7102 | n7103;
  assign n7106 = ~n7104 & n7105;
  assign n7107 = n13051 & n7106;
  assign n7108 = n13051 | n7106;
  assign n7109 = ~n7107 & n7108;
  assign n7110 = x49 & x106;
  assign n7111 = n7109 & n7110;
  assign n7112 = n7109 | n7110;
  assign n7113 = ~n7111 & n7112;
  assign n7114 = n6906 & n7113;
  assign n7115 = n6906 | n7113;
  assign n7116 = ~n7114 & n7115;
  assign n7117 = x48 & x107;
  assign n7118 = n7116 & n7117;
  assign n7119 = n7116 | n7117;
  assign n7120 = ~n7118 & n7119;
  assign n17727 = n6905 | n7110;
  assign n17728 = (n6904 & n7110) | (n6904 & n17727) | (n7110 & n17727);
  assign n16273 = (n6906 & n7109) | (n6906 & n17728) | (n7109 & n17728);
  assign n13135 = (n7111 & n7113) | (n7111 & n16273) | (n7113 & n16273);
  assign n13136 = n7104 | n13051;
  assign n13137 = (n7104 & n7106) | (n7104 & n13136) | (n7106 & n13136);
  assign n13138 = n7097 | n13053;
  assign n13139 = (n7097 & n7099) | (n7097 & n13138) | (n7099 & n13138);
  assign n13140 = n7090 | n13055;
  assign n13141 = (n7090 & n7092) | (n7090 & n13140) | (n7092 & n13140);
  assign n13142 = n7083 | n13057;
  assign n13143 = (n7083 & n7085) | (n7083 & n13142) | (n7085 & n13142);
  assign n16274 = n7076 | n16228;
  assign n16275 = (n7076 & n7078) | (n7076 & n16274) | (n7078 & n16274);
  assign n13144 = n7069 | n7071;
  assign n13145 = (n6914 & n7069) | (n6914 & n13144) | (n7069 & n13144);
  assign n13146 = n7062 | n7064;
  assign n13147 = (n7062 & n13059) | (n7062 & n13146) | (n13059 & n13146);
  assign n13148 = n7055 | n7057;
  assign n13149 = (n7055 & n13061) | (n7055 & n13148) | (n13061 & n13148);
  assign n13150 = n7048 | n7050;
  assign n13151 = (n7048 & n13063) | (n7048 & n13150) | (n13063 & n13150);
  assign n13152 = n7041 | n7043;
  assign n13153 = (n7041 & n13065) | (n7041 & n13152) | (n13065 & n13152);
  assign n13154 = n7034 | n7036;
  assign n13155 = (n7034 & n13067) | (n7034 & n13154) | (n13067 & n13154);
  assign n13156 = n7027 | n7029;
  assign n13157 = (n7027 & n13069) | (n7027 & n13156) | (n13069 & n13156);
  assign n13073 = (n6808 & n12991) | (n6808 & n13072) | (n12991 & n13072);
  assign n13075 = (n6801 & n12993) | (n6801 & n13074) | (n12993 & n13074);
  assign n13165 = n6992 | n6994;
  assign n16276 = n6787 | n6992;
  assign n16277 = (n6992 & n6994) | (n6992 & n16276) | (n6994 & n16276);
  assign n16278 = (n13045 & n13165) | (n13045 & n16277) | (n13165 & n16277);
  assign n16279 = (n13044 & n13165) | (n13044 & n16277) | (n13165 & n16277);
  assign n16280 = (n16123 & n16278) | (n16123 & n16279) | (n16278 & n16279);
  assign n13170 = n6971 | n6973;
  assign n16281 = n6766 | n6971;
  assign n16282 = (n6971 & n6973) | (n6971 & n16281) | (n6973 & n16281);
  assign n16283 = (n13035 & n13170) | (n13035 & n16282) | (n13170 & n16282);
  assign n16284 = (n13034 & n13170) | (n13034 & n16282) | (n13170 & n16282);
  assign n16285 = (n16128 & n16283) | (n16128 & n16284) | (n16283 & n16284);
  assign n16286 = n6759 | n6964;
  assign n16287 = (n6964 & n6966) | (n6964 & n16286) | (n6966 & n16286);
  assign n13173 = n6964 | n13108;
  assign n13174 = (n16187 & n16287) | (n16187 & n13173) | (n16287 & n13173);
  assign n7147 = x76 & x80;
  assign n7148 = x75 & x81;
  assign n7149 = n7147 & n7148;
  assign n7150 = n7147 | n7148;
  assign n7151 = ~n7149 & n7150;
  assign n16288 = n6936 | n6938;
  assign n16290 = n7151 & n16288;
  assign n16291 = n6936 & n7151;
  assign n16292 = (n16245 & n16290) | (n16245 & n16291) | (n16290 & n16291);
  assign n16293 = (n6936 & n16247) | (n6936 & n16288) | (n16247 & n16288);
  assign n13186 = n7151 & n16293;
  assign n13187 = (n16133 & n16292) | (n16133 & n13186) | (n16292 & n13186);
  assign n16294 = n7151 | n16288;
  assign n16295 = n6936 | n7151;
  assign n16296 = (n16245 & n16294) | (n16245 & n16295) | (n16294 & n16295);
  assign n13189 = n7151 | n16293;
  assign n13190 = (n16133 & n16296) | (n16133 & n13189) | (n16296 & n13189);
  assign n7154 = ~n13187 & n13190;
  assign n7155 = x74 & x82;
  assign n7156 = n7154 & n7155;
  assign n7157 = n7154 | n7155;
  assign n7158 = ~n7156 & n7157;
  assign n16297 = n6943 | n6945;
  assign n16298 = (n6943 & n13091) | (n6943 & n16297) | (n13091 & n16297);
  assign n13191 = n7158 & n16298;
  assign n16299 = n6738 | n6943;
  assign n16300 = (n6943 & n6945) | (n6943 & n16299) | (n6945 & n16299);
  assign n13192 = n7158 & n16300;
  assign n13193 = (n16192 & n13191) | (n16192 & n13192) | (n13191 & n13192);
  assign n13194 = n7158 | n16298;
  assign n13195 = n7158 | n16300;
  assign n13196 = (n16192 & n13194) | (n16192 & n13195) | (n13194 & n13195);
  assign n7161 = ~n13193 & n13196;
  assign n7162 = x73 & x83;
  assign n7163 = n7161 & n7162;
  assign n7164 = n7161 | n7162;
  assign n7165 = ~n7163 & n7164;
  assign n13177 = n6950 | n6952;
  assign n13197 = n7165 & n13177;
  assign n13198 = n6950 & n7165;
  assign n13199 = (n16243 & n13197) | (n16243 & n13198) | (n13197 & n13198);
  assign n13200 = n7165 | n13177;
  assign n13201 = n6950 | n7165;
  assign n13202 = (n16243 & n13200) | (n16243 & n13201) | (n13200 & n13201);
  assign n7168 = ~n13199 & n13202;
  assign n7169 = x72 & x84;
  assign n7170 = n7168 & n7169;
  assign n7171 = n7168 | n7169;
  assign n7172 = ~n7170 & n7171;
  assign n13175 = n6957 | n6959;
  assign n13203 = n7172 & n13175;
  assign n13204 = n6957 & n7172;
  assign n13205 = (n16240 & n13203) | (n16240 & n13204) | (n13203 & n13204);
  assign n13206 = n7172 | n13175;
  assign n13207 = n6957 | n7172;
  assign n13208 = (n16240 & n13206) | (n16240 & n13207) | (n13206 & n13207);
  assign n7175 = ~n13205 & n13208;
  assign n7176 = x71 & x85;
  assign n7177 = n7175 & n7176;
  assign n7178 = n7175 | n7176;
  assign n7179 = ~n7177 & n7178;
  assign n7180 = n13174 & n7179;
  assign n7181 = n13174 | n7179;
  assign n7182 = ~n7180 & n7181;
  assign n7183 = x70 & x86;
  assign n7184 = n7182 & n7183;
  assign n7185 = n7182 | n7183;
  assign n7186 = ~n7184 & n7185;
  assign n7187 = n16285 & n7186;
  assign n7188 = n16285 | n7186;
  assign n7189 = ~n7187 & n7188;
  assign n7190 = x69 & x87;
  assign n7191 = n7189 & n7190;
  assign n7192 = n7189 | n7190;
  assign n7193 = ~n7191 & n7192;
  assign n13167 = n6978 | n6980;
  assign n13209 = n7193 & n13167;
  assign n13210 = n6978 & n7193;
  assign n13211 = (n16233 & n13209) | (n16233 & n13210) | (n13209 & n13210);
  assign n13212 = n7193 | n13167;
  assign n13213 = n6978 | n7193;
  assign n13214 = (n16233 & n13212) | (n16233 & n13213) | (n13212 & n13213);
  assign n7196 = ~n13211 & n13214;
  assign n7197 = x68 & x88;
  assign n7198 = n7196 & n7197;
  assign n7199 = n7196 | n7197;
  assign n7200 = ~n7198 & n7199;
  assign n13215 = n6985 & n7200;
  assign n16301 = (n7200 & n13119) | (n7200 & n13215) | (n13119 & n13215);
  assign n16302 = (n7200 & n13118) | (n7200 & n13215) | (n13118 & n13215);
  assign n16303 = (n16182 & n16301) | (n16182 & n16302) | (n16301 & n16302);
  assign n13217 = n6985 | n7200;
  assign n16304 = n13119 | n13217;
  assign n16305 = n13118 | n13217;
  assign n16306 = (n16182 & n16304) | (n16182 & n16305) | (n16304 & n16305);
  assign n7203 = ~n16303 & n16306;
  assign n7204 = x67 & x89;
  assign n7205 = n7203 & n7204;
  assign n7206 = n7203 | n7204;
  assign n7207 = ~n7205 & n7206;
  assign n7208 = n16280 & n7207;
  assign n7209 = n16280 | n7207;
  assign n7210 = ~n7208 & n7209;
  assign n7211 = x66 & x90;
  assign n7212 = n7210 & n7211;
  assign n7213 = n7210 | n7211;
  assign n7214 = ~n7212 & n7213;
  assign n13219 = n6999 & n7214;
  assign n16307 = (n7214 & n13128) | (n7214 & n13219) | (n13128 & n13219);
  assign n16308 = (n7214 & n13129) | (n7214 & n13219) | (n13129 & n13219);
  assign n16309 = (n12995 & n16307) | (n12995 & n16308) | (n16307 & n16308);
  assign n13221 = n6999 | n7214;
  assign n16310 = n13128 | n13221;
  assign n16311 = n13129 | n13221;
  assign n16312 = (n12995 & n16310) | (n12995 & n16311) | (n16310 & n16311);
  assign n7217 = ~n16309 & n16312;
  assign n7218 = x65 & x91;
  assign n7219 = n7217 & n7218;
  assign n7220 = n7217 | n7218;
  assign n7221 = ~n7219 & n7220;
  assign n13162 = n7006 | n7008;
  assign n13223 = n7221 & n13162;
  assign n13224 = n7006 & n7221;
  assign n13225 = (n13075 & n13223) | (n13075 & n13224) | (n13223 & n13224);
  assign n13226 = n7221 | n13162;
  assign n13227 = n7006 | n7221;
  assign n13228 = (n13075 & n13226) | (n13075 & n13227) | (n13226 & n13227);
  assign n7224 = ~n13225 & n13228;
  assign n7225 = x64 & x92;
  assign n7226 = n7224 & n7225;
  assign n7227 = n7224 | n7225;
  assign n7228 = ~n7226 & n7227;
  assign n13160 = n7013 | n7015;
  assign n16313 = n7228 & n13160;
  assign n16314 = n7013 & n7228;
  assign n16315 = (n13073 & n16313) | (n13073 & n16314) | (n16313 & n16314);
  assign n16316 = n7228 | n13160;
  assign n16317 = n7013 | n7228;
  assign n16318 = (n13073 & n16316) | (n13073 & n16317) | (n16316 & n16317);
  assign n7231 = ~n16315 & n16318;
  assign n7232 = x63 & x93;
  assign n7233 = n7231 & n7232;
  assign n7234 = n7231 | n7232;
  assign n7235 = ~n7233 & n7234;
  assign n13158 = n7020 | n7022;
  assign n16319 = n7235 & n13158;
  assign n16320 = n7020 & n7235;
  assign n16321 = (n13071 & n16319) | (n13071 & n16320) | (n16319 & n16320);
  assign n16322 = n7235 | n13158;
  assign n16323 = n7020 | n7235;
  assign n16324 = (n13071 & n16322) | (n13071 & n16323) | (n16322 & n16323);
  assign n7238 = ~n16321 & n16324;
  assign n7239 = x62 & x94;
  assign n7240 = n7238 & n7239;
  assign n7241 = n7238 | n7239;
  assign n7242 = ~n7240 & n7241;
  assign n7243 = n13157 & n7242;
  assign n7244 = n13157 | n7242;
  assign n7245 = ~n7243 & n7244;
  assign n7246 = x61 & x95;
  assign n7247 = n7245 & n7246;
  assign n7248 = n7245 | n7246;
  assign n7249 = ~n7247 & n7248;
  assign n7250 = n13155 & n7249;
  assign n7251 = n13155 | n7249;
  assign n7252 = ~n7250 & n7251;
  assign n7253 = x60 & x96;
  assign n7254 = n7252 & n7253;
  assign n7255 = n7252 | n7253;
  assign n7256 = ~n7254 & n7255;
  assign n7257 = n13153 & n7256;
  assign n7258 = n13153 | n7256;
  assign n7259 = ~n7257 & n7258;
  assign n7260 = x59 & x97;
  assign n7261 = n7259 & n7260;
  assign n7262 = n7259 | n7260;
  assign n7263 = ~n7261 & n7262;
  assign n7264 = n13151 & n7263;
  assign n7265 = n13151 | n7263;
  assign n7266 = ~n7264 & n7265;
  assign n7267 = x58 & x98;
  assign n7268 = n7266 & n7267;
  assign n7269 = n7266 | n7267;
  assign n7270 = ~n7268 & n7269;
  assign n7271 = n13149 & n7270;
  assign n7272 = n13149 | n7270;
  assign n7273 = ~n7271 & n7272;
  assign n7274 = x57 & x99;
  assign n7275 = n7273 & n7274;
  assign n7276 = n7273 | n7274;
  assign n7277 = ~n7275 & n7276;
  assign n7278 = n13147 & n7277;
  assign n7279 = n13147 | n7277;
  assign n7280 = ~n7278 & n7279;
  assign n7281 = x56 & x100;
  assign n7282 = n7280 & n7281;
  assign n7283 = n7280 | n7281;
  assign n7284 = ~n7282 & n7283;
  assign n7285 = n13145 & n7284;
  assign n7286 = n13145 | n7284;
  assign n7287 = ~n7285 & n7286;
  assign n7288 = x55 & x101;
  assign n7289 = n7287 & n7288;
  assign n7290 = n7287 | n7288;
  assign n7291 = ~n7289 & n7290;
  assign n7292 = n16275 & n7291;
  assign n7293 = n16275 | n7291;
  assign n7294 = ~n7292 & n7293;
  assign n7295 = x54 & x102;
  assign n7296 = n7294 & n7295;
  assign n7297 = n7294 | n7295;
  assign n7298 = ~n7296 & n7297;
  assign n7299 = n13143 & n7298;
  assign n7300 = n13143 | n7298;
  assign n7301 = ~n7299 & n7300;
  assign n7302 = x53 & x103;
  assign n7303 = n7301 & n7302;
  assign n7304 = n7301 | n7302;
  assign n7305 = ~n7303 & n7304;
  assign n7306 = n13141 & n7305;
  assign n7307 = n13141 | n7305;
  assign n7308 = ~n7306 & n7307;
  assign n7309 = x52 & x104;
  assign n7310 = n7308 & n7309;
  assign n7311 = n7308 | n7309;
  assign n7312 = ~n7310 & n7311;
  assign n7313 = n13139 & n7312;
  assign n7314 = n13139 | n7312;
  assign n7315 = ~n7313 & n7314;
  assign n7316 = x51 & x105;
  assign n7317 = n7315 & n7316;
  assign n7318 = n7315 | n7316;
  assign n7319 = ~n7317 & n7318;
  assign n7320 = n13137 & n7319;
  assign n7321 = n13137 | n7319;
  assign n7322 = ~n7320 & n7321;
  assign n7323 = x50 & x106;
  assign n7324 = n7322 & n7323;
  assign n7325 = n7322 | n7323;
  assign n7326 = ~n7324 & n7325;
  assign n7327 = n13135 & n7326;
  assign n7328 = n13135 | n7326;
  assign n7329 = ~n7327 & n7328;
  assign n7330 = x49 & x107;
  assign n7331 = n7329 & n7330;
  assign n7332 = n7329 | n7330;
  assign n7333 = ~n7331 & n7332;
  assign n7334 = n7118 & n7333;
  assign n7335 = n7118 | n7333;
  assign n7336 = ~n7334 & n7335;
  assign n7337 = x48 & x108;
  assign n7338 = n7336 & n7337;
  assign n7339 = n7336 | n7337;
  assign n7340 = ~n7338 & n7339;
  assign n13229 = n7118 | n7331;
  assign n13230 = (n7331 & n7333) | (n7331 & n13229) | (n7333 & n13229);
  assign n13231 = n7324 | n13135;
  assign n13232 = (n7324 & n7326) | (n7324 & n13231) | (n7326 & n13231);
  assign n13233 = n7317 | n13137;
  assign n13234 = (n7317 & n7319) | (n7317 & n13233) | (n7319 & n13233);
  assign n13235 = n7310 | n13139;
  assign n13236 = (n7310 & n7312) | (n7310 & n13235) | (n7312 & n13235);
  assign n13237 = n7303 | n13141;
  assign n13238 = (n7303 & n7305) | (n7303 & n13237) | (n7305 & n13237);
  assign n13239 = n7296 | n13143;
  assign n13240 = (n7296 & n7298) | (n7296 & n13239) | (n7298 & n13239);
  assign n13241 = n7289 | n7291;
  assign n13242 = (n16275 & n7289) | (n16275 & n13241) | (n7289 & n13241);
  assign n13243 = n7282 | n7284;
  assign n13244 = (n7282 & n13145) | (n7282 & n13243) | (n13145 & n13243);
  assign n13245 = n7275 | n7277;
  assign n13246 = (n7275 & n13147) | (n7275 & n13245) | (n13147 & n13245);
  assign n13247 = n7268 | n7270;
  assign n13248 = (n7268 & n13149) | (n7268 & n13247) | (n13149 & n13247);
  assign n13249 = n7261 | n7263;
  assign n13250 = (n7261 & n13151) | (n7261 & n13249) | (n13151 & n13249);
  assign n13251 = n7254 | n7256;
  assign n13252 = (n7254 & n13153) | (n7254 & n13251) | (n13153 & n13251);
  assign n13253 = n7247 | n7249;
  assign n13254 = (n7247 & n13155) | (n7247 & n13253) | (n13155 & n13253);
  assign n13159 = (n7020 & n13071) | (n7020 & n13158) | (n13071 & n13158);
  assign n13161 = (n7013 & n13073) | (n7013 & n13160) | (n13073 & n13160);
  assign n13264 = n7198 | n7200;
  assign n16325 = n6985 | n7198;
  assign n16326 = (n7198 & n7200) | (n7198 & n16325) | (n7200 & n16325);
  assign n16327 = (n13119 & n13264) | (n13119 & n16326) | (n13264 & n16326);
  assign n16328 = (n13118 & n13264) | (n13118 & n16326) | (n13264 & n16326);
  assign n16329 = (n16182 & n16327) | (n16182 & n16328) | (n16327 & n16328);
  assign n7368 = x77 & x80;
  assign n7369 = x76 & x81;
  assign n7370 = n7368 & n7369;
  assign n7371 = n7368 | n7369;
  assign n7372 = ~n7370 & n7371;
  assign n16337 = n7149 & n7372;
  assign n16338 = (n7372 & n16292) | (n7372 & n16337) | (n16292 & n16337);
  assign n16339 = n7149 | n7151;
  assign n16341 = n7372 & n16339;
  assign n16342 = (n16293 & n16337) | (n16293 & n16341) | (n16337 & n16341);
  assign n13284 = (n16133 & n16338) | (n16133 & n16342) | (n16338 & n16342);
  assign n16343 = n7149 | n7372;
  assign n16344 = n16292 | n16343;
  assign n16345 = n7372 | n16339;
  assign n16346 = (n16293 & n16343) | (n16293 & n16345) | (n16343 & n16345);
  assign n13287 = (n16133 & n16344) | (n16133 & n16346) | (n16344 & n16346);
  assign n7375 = ~n13284 & n13287;
  assign n7376 = x75 & x82;
  assign n7377 = n7375 & n7376;
  assign n7378 = n7375 | n7376;
  assign n7379 = ~n7377 & n7378;
  assign n16334 = n7156 | n7158;
  assign n17729 = n7379 & n16334;
  assign n17730 = n7156 & n7379;
  assign n17731 = (n16298 & n17729) | (n16298 & n17730) | (n17729 & n17730);
  assign n16336 = (n7156 & n16300) | (n7156 & n16334) | (n16300 & n16334);
  assign n16348 = n7379 & n16336;
  assign n16349 = (n16192 & n17731) | (n16192 & n16348) | (n17731 & n16348);
  assign n17732 = n7379 | n16334;
  assign n17733 = n7156 | n7379;
  assign n17734 = (n16298 & n17732) | (n16298 & n17733) | (n17732 & n17733);
  assign n16351 = n7379 | n16336;
  assign n16352 = (n16192 & n17734) | (n16192 & n16351) | (n17734 & n16351);
  assign n7382 = ~n16349 & n16352;
  assign n7383 = x74 & x83;
  assign n7384 = n7382 & n7383;
  assign n7385 = n7382 | n7383;
  assign n7386 = ~n7384 & n7385;
  assign n16353 = n7163 | n7165;
  assign n16354 = (n7163 & n13177) | (n7163 & n16353) | (n13177 & n16353);
  assign n13288 = n7386 & n16354;
  assign n16355 = n6950 | n7163;
  assign n16356 = (n7163 & n7165) | (n7163 & n16355) | (n7165 & n16355);
  assign n13289 = n7386 & n16356;
  assign n13290 = (n16243 & n13288) | (n16243 & n13289) | (n13288 & n13289);
  assign n13291 = n7386 | n16354;
  assign n13292 = n7386 | n16356;
  assign n13293 = (n16243 & n13291) | (n16243 & n13292) | (n13291 & n13292);
  assign n7389 = ~n13290 & n13293;
  assign n7390 = x73 & x84;
  assign n7391 = n7389 & n7390;
  assign n7392 = n7389 | n7390;
  assign n7393 = ~n7391 & n7392;
  assign n16330 = n7170 | n7172;
  assign n16331 = (n7170 & n13175) | (n7170 & n16330) | (n13175 & n16330);
  assign n16357 = n7393 & n16331;
  assign n16332 = n6957 | n7170;
  assign n16333 = (n7170 & n7172) | (n7170 & n16332) | (n7172 & n16332);
  assign n16358 = n7393 & n16333;
  assign n16359 = (n16240 & n16357) | (n16240 & n16358) | (n16357 & n16358);
  assign n16360 = n7393 | n16331;
  assign n16361 = n7393 | n16333;
  assign n16362 = (n16240 & n16360) | (n16240 & n16361) | (n16360 & n16361);
  assign n7396 = ~n16359 & n16362;
  assign n7397 = x72 & x85;
  assign n7398 = n7396 & n7397;
  assign n7399 = n7396 | n7397;
  assign n7400 = ~n7398 & n7399;
  assign n13268 = n7177 | n7179;
  assign n13294 = n7400 & n13268;
  assign n13295 = n7177 & n7400;
  assign n13296 = (n13174 & n13294) | (n13174 & n13295) | (n13294 & n13295);
  assign n13297 = n7400 | n13268;
  assign n13298 = n7177 | n7400;
  assign n13299 = (n13174 & n13297) | (n13174 & n13298) | (n13297 & n13298);
  assign n7403 = ~n13296 & n13299;
  assign n7404 = x71 & x86;
  assign n7405 = n7403 & n7404;
  assign n7406 = n7403 | n7404;
  assign n7407 = ~n7405 & n7406;
  assign n13266 = n7184 | n7186;
  assign n13300 = n7407 & n13266;
  assign n13301 = n7184 & n7407;
  assign n13302 = (n16285 & n13300) | (n16285 & n13301) | (n13300 & n13301);
  assign n13303 = n7407 | n13266;
  assign n13304 = n7184 | n7407;
  assign n13305 = (n16285 & n13303) | (n16285 & n13304) | (n13303 & n13304);
  assign n7410 = ~n13302 & n13305;
  assign n7411 = x70 & x87;
  assign n7412 = n7410 & n7411;
  assign n7413 = n7410 | n7411;
  assign n7414 = ~n7412 & n7413;
  assign n13306 = n7191 & n7414;
  assign n16363 = (n7414 & n13210) | (n7414 & n13306) | (n13210 & n13306);
  assign n16364 = (n7414 & n13209) | (n7414 & n13306) | (n13209 & n13306);
  assign n16365 = (n16233 & n16363) | (n16233 & n16364) | (n16363 & n16364);
  assign n13308 = n7191 | n7414;
  assign n16366 = n13210 | n13308;
  assign n16367 = n13209 | n13308;
  assign n16368 = (n16233 & n16366) | (n16233 & n16367) | (n16366 & n16367);
  assign n7417 = ~n16365 & n16368;
  assign n7418 = x69 & x88;
  assign n7419 = n7417 & n7418;
  assign n7420 = n7417 | n7418;
  assign n7421 = ~n7419 & n7420;
  assign n7422 = n16329 & n7421;
  assign n7423 = n16329 | n7421;
  assign n7424 = ~n7422 & n7423;
  assign n7425 = x68 & x89;
  assign n7426 = n7424 & n7425;
  assign n7427 = n7424 | n7425;
  assign n7428 = ~n7426 & n7427;
  assign n13261 = n7205 | n7207;
  assign n13310 = n7428 & n13261;
  assign n13311 = n7205 & n7428;
  assign n13312 = (n16280 & n13310) | (n16280 & n13311) | (n13310 & n13311);
  assign n13313 = n7428 | n13261;
  assign n13314 = n7205 | n7428;
  assign n13315 = (n16280 & n13313) | (n16280 & n13314) | (n13313 & n13314);
  assign n7431 = ~n13312 & n13315;
  assign n7432 = x67 & x90;
  assign n7433 = n7431 & n7432;
  assign n7434 = n7431 | n7432;
  assign n7435 = ~n7433 & n7434;
  assign n13316 = n7212 & n7435;
  assign n13317 = (n7435 & n16309) | (n7435 & n13316) | (n16309 & n13316);
  assign n13318 = n7212 | n7435;
  assign n13319 = n16309 | n13318;
  assign n7438 = ~n13317 & n13319;
  assign n7439 = x66 & x91;
  assign n7440 = n7438 & n7439;
  assign n7441 = n7438 | n7439;
  assign n7442 = ~n7440 & n7441;
  assign n13320 = n7219 & n7442;
  assign n13321 = (n7442 & n13225) | (n7442 & n13320) | (n13225 & n13320);
  assign n13322 = n7219 | n7442;
  assign n13323 = n13225 | n13322;
  assign n7445 = ~n13321 & n13323;
  assign n7446 = x65 & x92;
  assign n7447 = n7445 & n7446;
  assign n7448 = n7445 | n7446;
  assign n7449 = ~n7447 & n7448;
  assign n13259 = n7226 | n7228;
  assign n13324 = n7449 & n13259;
  assign n13325 = n7226 & n7449;
  assign n13326 = (n13161 & n13324) | (n13161 & n13325) | (n13324 & n13325);
  assign n13327 = n7449 | n13259;
  assign n13328 = n7226 | n7449;
  assign n13329 = (n13161 & n13327) | (n13161 & n13328) | (n13327 & n13328);
  assign n7452 = ~n13326 & n13329;
  assign n7453 = x64 & x93;
  assign n7454 = n7452 & n7453;
  assign n7455 = n7452 | n7453;
  assign n7456 = ~n7454 & n7455;
  assign n13257 = n7233 | n7235;
  assign n16369 = n7456 & n13257;
  assign n16370 = n7233 & n7456;
  assign n16371 = (n13159 & n16369) | (n13159 & n16370) | (n16369 & n16370);
  assign n16372 = n7456 | n13257;
  assign n16373 = n7233 | n7456;
  assign n16374 = (n13159 & n16372) | (n13159 & n16373) | (n16372 & n16373);
  assign n7459 = ~n16371 & n16374;
  assign n7460 = x63 & x94;
  assign n7461 = n7459 & n7460;
  assign n7462 = n7459 | n7460;
  assign n7463 = ~n7461 & n7462;
  assign n13255 = n7240 | n7242;
  assign n16375 = n7463 & n13255;
  assign n16376 = n7240 & n7463;
  assign n16377 = (n13157 & n16375) | (n13157 & n16376) | (n16375 & n16376);
  assign n16378 = n7463 | n13255;
  assign n16379 = n7240 | n7463;
  assign n16380 = (n13157 & n16378) | (n13157 & n16379) | (n16378 & n16379);
  assign n7466 = ~n16377 & n16380;
  assign n7467 = x62 & x95;
  assign n7468 = n7466 & n7467;
  assign n7469 = n7466 | n7467;
  assign n7470 = ~n7468 & n7469;
  assign n7471 = n13254 & n7470;
  assign n7472 = n13254 | n7470;
  assign n7473 = ~n7471 & n7472;
  assign n7474 = x61 & x96;
  assign n7475 = n7473 & n7474;
  assign n7476 = n7473 | n7474;
  assign n7477 = ~n7475 & n7476;
  assign n7478 = n13252 & n7477;
  assign n7479 = n13252 | n7477;
  assign n7480 = ~n7478 & n7479;
  assign n7481 = x60 & x97;
  assign n7482 = n7480 & n7481;
  assign n7483 = n7480 | n7481;
  assign n7484 = ~n7482 & n7483;
  assign n7485 = n13250 & n7484;
  assign n7486 = n13250 | n7484;
  assign n7487 = ~n7485 & n7486;
  assign n7488 = x59 & x98;
  assign n7489 = n7487 & n7488;
  assign n7490 = n7487 | n7488;
  assign n7491 = ~n7489 & n7490;
  assign n7492 = n13248 & n7491;
  assign n7493 = n13248 | n7491;
  assign n7494 = ~n7492 & n7493;
  assign n7495 = x58 & x99;
  assign n7496 = n7494 & n7495;
  assign n7497 = n7494 | n7495;
  assign n7498 = ~n7496 & n7497;
  assign n7499 = n13246 & n7498;
  assign n7500 = n13246 | n7498;
  assign n7501 = ~n7499 & n7500;
  assign n7502 = x57 & x100;
  assign n7503 = n7501 & n7502;
  assign n7504 = n7501 | n7502;
  assign n7505 = ~n7503 & n7504;
  assign n7506 = n13244 & n7505;
  assign n7507 = n13244 | n7505;
  assign n7508 = ~n7506 & n7507;
  assign n7509 = x56 & x101;
  assign n7510 = n7508 & n7509;
  assign n7511 = n7508 | n7509;
  assign n7512 = ~n7510 & n7511;
  assign n7513 = n13242 & n7512;
  assign n7514 = n13242 | n7512;
  assign n7515 = ~n7513 & n7514;
  assign n7516 = x55 & x102;
  assign n7517 = n7515 & n7516;
  assign n7518 = n7515 | n7516;
  assign n7519 = ~n7517 & n7518;
  assign n7520 = n13240 & n7519;
  assign n7521 = n13240 | n7519;
  assign n7522 = ~n7520 & n7521;
  assign n7523 = x54 & x103;
  assign n7524 = n7522 & n7523;
  assign n7525 = n7522 | n7523;
  assign n7526 = ~n7524 & n7525;
  assign n7527 = n13238 & n7526;
  assign n7528 = n13238 | n7526;
  assign n7529 = ~n7527 & n7528;
  assign n7530 = x53 & x104;
  assign n7531 = n7529 & n7530;
  assign n7532 = n7529 | n7530;
  assign n7533 = ~n7531 & n7532;
  assign n7534 = n13236 & n7533;
  assign n7535 = n13236 | n7533;
  assign n7536 = ~n7534 & n7535;
  assign n7537 = x52 & x105;
  assign n7538 = n7536 & n7537;
  assign n7539 = n7536 | n7537;
  assign n7540 = ~n7538 & n7539;
  assign n7541 = n13234 & n7540;
  assign n7542 = n13234 | n7540;
  assign n7543 = ~n7541 & n7542;
  assign n7544 = x51 & x106;
  assign n7545 = n7543 & n7544;
  assign n7546 = n7543 | n7544;
  assign n7547 = ~n7545 & n7546;
  assign n7548 = n13232 & n7547;
  assign n7549 = n13232 | n7547;
  assign n7550 = ~n7548 & n7549;
  assign n7551 = x50 & x107;
  assign n7552 = n7550 & n7551;
  assign n7553 = n7550 | n7551;
  assign n7554 = ~n7552 & n7553;
  assign n7555 = n13230 & n7554;
  assign n7556 = n13230 | n7554;
  assign n7557 = ~n7555 & n7556;
  assign n7558 = x49 & x108;
  assign n7559 = n7557 & n7558;
  assign n7560 = n7557 | n7558;
  assign n7561 = ~n7559 & n7560;
  assign n7562 = n7338 & n7561;
  assign n7563 = n7338 | n7561;
  assign n7564 = ~n7562 & n7563;
  assign n7565 = x48 & x109;
  assign n7566 = n7564 & n7565;
  assign n7567 = n7564 | n7565;
  assign n7568 = ~n7566 & n7567;
  assign n17735 = n7337 | n7558;
  assign n17736 = (n7336 & n7558) | (n7336 & n17735) | (n7558 & n17735);
  assign n16382 = (n7338 & n7557) | (n7338 & n17736) | (n7557 & n17736);
  assign n13331 = (n7559 & n7561) | (n7559 & n16382) | (n7561 & n16382);
  assign n16383 = n7552 | n13230;
  assign n16384 = (n7552 & n7554) | (n7552 & n16383) | (n7554 & n16383);
  assign n7571 = n7545 | n7548;
  assign n7572 = n7538 | n7541;
  assign n7573 = n7531 | n7534;
  assign n7574 = n7524 | n7527;
  assign n7575 = n7517 | n7520;
  assign n13332 = n7510 | n7512;
  assign n13333 = (n7510 & n13242) | (n7510 & n13332) | (n13242 & n13332);
  assign n13334 = n7503 | n7505;
  assign n13335 = (n7503 & n13244) | (n7503 & n13334) | (n13244 & n13334);
  assign n13336 = n7496 | n7498;
  assign n13337 = (n7496 & n13246) | (n7496 & n13336) | (n13246 & n13336);
  assign n13338 = n7489 | n7491;
  assign n13339 = (n7489 & n13248) | (n7489 & n13338) | (n13248 & n13338);
  assign n13340 = n7482 | n7484;
  assign n13341 = (n7482 & n13250) | (n7482 & n13340) | (n13250 & n13340);
  assign n13342 = n7475 | n7477;
  assign n13343 = (n7475 & n13252) | (n7475 & n13342) | (n13252 & n13342);
  assign n13256 = (n7240 & n13157) | (n7240 & n13255) | (n13157 & n13255);
  assign n13258 = (n7233 & n13159) | (n7233 & n13257) | (n13159 & n13257);
  assign n13356 = n7412 | n7414;
  assign n16387 = n7191 | n7412;
  assign n16388 = (n7412 & n7414) | (n7412 & n16387) | (n7414 & n16387);
  assign n16389 = (n13210 & n13356) | (n13210 & n16388) | (n13356 & n16388);
  assign n16390 = (n13209 & n13356) | (n13209 & n16388) | (n13356 & n16388);
  assign n16391 = (n16233 & n16389) | (n16233 & n16390) | (n16389 & n16390);
  assign n7597 = x78 & x80;
  assign n7598 = x77 & x81;
  assign n7599 = n7597 & n7598;
  assign n7600 = n7597 | n7598;
  assign n7601 = ~n7599 & n7600;
  assign n17737 = n7370 & n7601;
  assign n17738 = (n7601 & n16342) | (n7601 & n17737) | (n16342 & n17737);
  assign n16397 = n7370 | n7372;
  assign n17741 = n7601 & n16397;
  assign n17739 = n7149 | n7370;
  assign n17740 = (n7370 & n7372) | (n7370 & n17739) | (n7372 & n17739);
  assign n17742 = n7601 & n17740;
  assign n17743 = (n16292 & n17741) | (n16292 & n17742) | (n17741 & n17742);
  assign n16401 = (n16133 & n17738) | (n16133 & n17743) | (n17738 & n17743);
  assign n17744 = n7370 | n7601;
  assign n17745 = n16342 | n17744;
  assign n17746 = n7601 | n16397;
  assign n17747 = n7601 | n17740;
  assign n17748 = (n16292 & n17746) | (n16292 & n17747) | (n17746 & n17747);
  assign n16404 = (n16133 & n17745) | (n16133 & n17748) | (n17745 & n17748);
  assign n7604 = ~n16401 & n16404;
  assign n7605 = x76 & x82;
  assign n7606 = n7604 & n7605;
  assign n7607 = n7604 | n7605;
  assign n7608 = ~n7606 & n7607;
  assign n13363 = n7377 | n7379;
  assign n13368 = n7608 & n13363;
  assign n13369 = n7377 & n7608;
  assign n16335 = (n7156 & n16298) | (n7156 & n16334) | (n16298 & n16334);
  assign n16405 = (n13368 & n13369) | (n13368 & n16335) | (n13369 & n16335);
  assign n16406 = (n13368 & n13369) | (n13368 & n16336) | (n13369 & n16336);
  assign n16407 = (n16192 & n16405) | (n16192 & n16406) | (n16405 & n16406);
  assign n13371 = n7608 | n13363;
  assign n13372 = n7377 | n7608;
  assign n16408 = (n13371 & n13372) | (n13371 & n16335) | (n13372 & n16335);
  assign n16409 = (n13371 & n13372) | (n13371 & n16336) | (n13372 & n16336);
  assign n16410 = (n16192 & n16408) | (n16192 & n16409) | (n16408 & n16409);
  assign n7611 = ~n16407 & n16410;
  assign n7612 = x75 & x83;
  assign n7613 = n7611 & n7612;
  assign n7614 = n7611 | n7612;
  assign n7615 = ~n7613 & n7614;
  assign n13374 = n7384 & n7615;
  assign n17749 = (n7386 & n7615) | (n7386 & n13374) | (n7615 & n13374);
  assign n17750 = n7615 & n13374;
  assign n17751 = (n16354 & n17749) | (n16354 & n17750) | (n17749 & n17750);
  assign n16412 = (n7615 & n13289) | (n7615 & n13374) | (n13289 & n13374);
  assign n16413 = (n16243 & n17751) | (n16243 & n16412) | (n17751 & n16412);
  assign n13376 = n7384 | n7615;
  assign n17752 = n7386 | n13376;
  assign n17753 = (n13376 & n16354) | (n13376 & n17752) | (n16354 & n17752);
  assign n16415 = n13289 | n13376;
  assign n16416 = (n16243 & n17753) | (n16243 & n16415) | (n17753 & n16415);
  assign n7618 = ~n16413 & n16416;
  assign n7619 = x74 & x84;
  assign n7620 = n7618 & n7619;
  assign n7621 = n7618 | n7619;
  assign n7622 = ~n7620 & n7621;
  assign n13361 = n7391 | n7393;
  assign n13378 = n7622 & n13361;
  assign n13379 = n7391 & n7622;
  assign n16417 = (n13378 & n13379) | (n13378 & n16331) | (n13379 & n16331);
  assign n16418 = (n13378 & n13379) | (n13378 & n16333) | (n13379 & n16333);
  assign n16419 = (n16240 & n16417) | (n16240 & n16418) | (n16417 & n16418);
  assign n13381 = n7622 | n13361;
  assign n13382 = n7391 | n7622;
  assign n16420 = (n13381 & n13382) | (n13381 & n16331) | (n13382 & n16331);
  assign n16421 = (n13381 & n13382) | (n13381 & n16333) | (n13382 & n16333);
  assign n16422 = (n16240 & n16420) | (n16240 & n16421) | (n16420 & n16421);
  assign n7625 = ~n16419 & n16422;
  assign n7626 = x73 & x85;
  assign n7627 = n7625 & n7626;
  assign n7628 = n7625 | n7626;
  assign n7629 = ~n7627 & n7628;
  assign n16394 = n7398 | n7400;
  assign n16395 = (n7398 & n13268) | (n7398 & n16394) | (n13268 & n16394);
  assign n16423 = n7629 & n16395;
  assign n16392 = n7177 | n7398;
  assign n16393 = (n7398 & n7400) | (n7398 & n16392) | (n7400 & n16392);
  assign n16424 = n7629 & n16393;
  assign n16425 = (n13174 & n16423) | (n13174 & n16424) | (n16423 & n16424);
  assign n16426 = n7629 | n16395;
  assign n16427 = n7629 | n16393;
  assign n16428 = (n13174 & n16426) | (n13174 & n16427) | (n16426 & n16427);
  assign n7632 = ~n16425 & n16428;
  assign n7633 = x72 & x86;
  assign n7634 = n7632 & n7633;
  assign n7635 = n7632 | n7633;
  assign n7636 = ~n7634 & n7635;
  assign n13384 = n7405 & n7636;
  assign n13385 = (n7636 & n13302) | (n7636 & n13384) | (n13302 & n13384);
  assign n13386 = n7405 | n7636;
  assign n13387 = n13302 | n13386;
  assign n7639 = ~n13385 & n13387;
  assign n7640 = x71 & x87;
  assign n7641 = n7639 & n7640;
  assign n7642 = n7639 | n7640;
  assign n7643 = ~n7641 & n7642;
  assign n7644 = n16391 & n7643;
  assign n7645 = n16391 | n7643;
  assign n7646 = ~n7644 & n7645;
  assign n7647 = x70 & x88;
  assign n7648 = n7646 & n7647;
  assign n7649 = n7646 | n7647;
  assign n7650 = ~n7648 & n7649;
  assign n13353 = n7419 | n7421;
  assign n13388 = n7650 & n13353;
  assign n13389 = n7419 & n7650;
  assign n13390 = (n16329 & n13388) | (n16329 & n13389) | (n13388 & n13389);
  assign n13391 = n7650 | n13353;
  assign n13392 = n7419 | n7650;
  assign n13393 = (n16329 & n13391) | (n16329 & n13392) | (n13391 & n13392);
  assign n7653 = ~n13390 & n13393;
  assign n7654 = x69 & x89;
  assign n7655 = n7653 & n7654;
  assign n7656 = n7653 | n7654;
  assign n7657 = ~n7655 & n7656;
  assign n13394 = n7426 & n7657;
  assign n16429 = (n7657 & n13311) | (n7657 & n13394) | (n13311 & n13394);
  assign n16430 = (n7657 & n13310) | (n7657 & n13394) | (n13310 & n13394);
  assign n16431 = (n16280 & n16429) | (n16280 & n16430) | (n16429 & n16430);
  assign n13396 = n7426 | n7657;
  assign n16432 = n13311 | n13396;
  assign n16433 = n13310 | n13396;
  assign n16434 = (n16280 & n16432) | (n16280 & n16433) | (n16432 & n16433);
  assign n7660 = ~n16431 & n16434;
  assign n7661 = x68 & x90;
  assign n7662 = n7660 & n7661;
  assign n7663 = n7660 | n7661;
  assign n7664 = ~n7662 & n7663;
  assign n13351 = n7433 | n7435;
  assign n16435 = n7664 & n13351;
  assign n16385 = n7212 | n7433;
  assign n16386 = (n7433 & n7435) | (n7433 & n16385) | (n7435 & n16385);
  assign n16436 = n7664 & n16386;
  assign n16437 = (n16309 & n16435) | (n16309 & n16436) | (n16435 & n16436);
  assign n16438 = n7664 | n13351;
  assign n16439 = n7664 | n16386;
  assign n16440 = (n16309 & n16438) | (n16309 & n16439) | (n16438 & n16439);
  assign n7667 = ~n16437 & n16440;
  assign n7668 = x67 & x91;
  assign n7669 = n7667 & n7668;
  assign n7670 = n7667 | n7668;
  assign n7671 = ~n7669 & n7670;
  assign n13398 = n7440 & n7671;
  assign n16441 = (n7671 & n13320) | (n7671 & n13398) | (n13320 & n13398);
  assign n16442 = (n7442 & n7671) | (n7442 & n13398) | (n7671 & n13398);
  assign n16443 = (n13225 & n16441) | (n13225 & n16442) | (n16441 & n16442);
  assign n13400 = n7440 | n7671;
  assign n16444 = n13320 | n13400;
  assign n16445 = n7442 | n13400;
  assign n16446 = (n13225 & n16444) | (n13225 & n16445) | (n16444 & n16445);
  assign n7674 = ~n16443 & n16446;
  assign n7675 = x66 & x92;
  assign n7676 = n7674 & n7675;
  assign n7677 = n7674 | n7675;
  assign n7678 = ~n7676 & n7677;
  assign n13402 = n7447 & n7678;
  assign n13403 = (n7678 & n13326) | (n7678 & n13402) | (n13326 & n13402);
  assign n13404 = n7447 | n7678;
  assign n13405 = n13326 | n13404;
  assign n7681 = ~n13403 & n13405;
  assign n7682 = x65 & x93;
  assign n7683 = n7681 & n7682;
  assign n7684 = n7681 | n7682;
  assign n7685 = ~n7683 & n7684;
  assign n13348 = n7454 | n7456;
  assign n13406 = n7685 & n13348;
  assign n13407 = n7454 & n7685;
  assign n13408 = (n13258 & n13406) | (n13258 & n13407) | (n13406 & n13407);
  assign n13409 = n7685 | n13348;
  assign n13410 = n7454 | n7685;
  assign n13411 = (n13258 & n13409) | (n13258 & n13410) | (n13409 & n13410);
  assign n7688 = ~n13408 & n13411;
  assign n7689 = x64 & x94;
  assign n7690 = n7688 & n7689;
  assign n7691 = n7688 | n7689;
  assign n7692 = ~n7690 & n7691;
  assign n13346 = n7461 | n7463;
  assign n16447 = n7692 & n13346;
  assign n16448 = n7461 & n7692;
  assign n16449 = (n13256 & n16447) | (n13256 & n16448) | (n16447 & n16448);
  assign n16450 = n7692 | n13346;
  assign n16451 = n7461 | n7692;
  assign n16452 = (n13256 & n16450) | (n13256 & n16451) | (n16450 & n16451);
  assign n7695 = ~n16449 & n16452;
  assign n7696 = x63 & x95;
  assign n7697 = n7695 & n7696;
  assign n7698 = n7695 | n7696;
  assign n7699 = ~n7697 & n7698;
  assign n13344 = n7468 | n7470;
  assign n16453 = n7699 & n13344;
  assign n16454 = n7468 & n7699;
  assign n16455 = (n13254 & n16453) | (n13254 & n16454) | (n16453 & n16454);
  assign n16456 = n7699 | n13344;
  assign n16457 = n7468 | n7699;
  assign n16458 = (n13254 & n16456) | (n13254 & n16457) | (n16456 & n16457);
  assign n7702 = ~n16455 & n16458;
  assign n7703 = x62 & x96;
  assign n7704 = n7702 & n7703;
  assign n7705 = n7702 | n7703;
  assign n7706 = ~n7704 & n7705;
  assign n7707 = n13343 & n7706;
  assign n7708 = n13343 | n7706;
  assign n7709 = ~n7707 & n7708;
  assign n7710 = x61 & x97;
  assign n7711 = n7709 & n7710;
  assign n7712 = n7709 | n7710;
  assign n7713 = ~n7711 & n7712;
  assign n7714 = n13341 & n7713;
  assign n7715 = n13341 | n7713;
  assign n7716 = ~n7714 & n7715;
  assign n7717 = x60 & x98;
  assign n7718 = n7716 & n7717;
  assign n7719 = n7716 | n7717;
  assign n7720 = ~n7718 & n7719;
  assign n7721 = n13339 & n7720;
  assign n7722 = n13339 | n7720;
  assign n7723 = ~n7721 & n7722;
  assign n7724 = x59 & x99;
  assign n7725 = n7723 & n7724;
  assign n7726 = n7723 | n7724;
  assign n7727 = ~n7725 & n7726;
  assign n7728 = n13337 & n7727;
  assign n7729 = n13337 | n7727;
  assign n7730 = ~n7728 & n7729;
  assign n7731 = x58 & x100;
  assign n7732 = n7730 & n7731;
  assign n7733 = n7730 | n7731;
  assign n7734 = ~n7732 & n7733;
  assign n7735 = n13335 & n7734;
  assign n7736 = n13335 | n7734;
  assign n7737 = ~n7735 & n7736;
  assign n7738 = x57 & x101;
  assign n7739 = n7737 & n7738;
  assign n7740 = n7737 | n7738;
  assign n7741 = ~n7739 & n7740;
  assign n7742 = n13333 & n7741;
  assign n7743 = n13333 | n7741;
  assign n7744 = ~n7742 & n7743;
  assign n7745 = x56 & x102;
  assign n7746 = n7744 & n7745;
  assign n7747 = n7744 | n7745;
  assign n7748 = ~n7746 & n7747;
  assign n7749 = n7575 & n7748;
  assign n7750 = n7575 | n7748;
  assign n7751 = ~n7749 & n7750;
  assign n7752 = x55 & x103;
  assign n7753 = n7751 & n7752;
  assign n7754 = n7751 | n7752;
  assign n7755 = ~n7753 & n7754;
  assign n7756 = n7574 & n7755;
  assign n7757 = n7574 | n7755;
  assign n7758 = ~n7756 & n7757;
  assign n7759 = x54 & x104;
  assign n7760 = n7758 & n7759;
  assign n7761 = n7758 | n7759;
  assign n7762 = ~n7760 & n7761;
  assign n7763 = n7573 & n7762;
  assign n7764 = n7573 | n7762;
  assign n7765 = ~n7763 & n7764;
  assign n7766 = x53 & x105;
  assign n7767 = n7765 & n7766;
  assign n7768 = n7765 | n7766;
  assign n7769 = ~n7767 & n7768;
  assign n7770 = n7572 & n7769;
  assign n7771 = n7572 | n7769;
  assign n7772 = ~n7770 & n7771;
  assign n7773 = x52 & x106;
  assign n7774 = n7772 & n7773;
  assign n7775 = n7772 | n7773;
  assign n7776 = ~n7774 & n7775;
  assign n7777 = n7571 & n7776;
  assign n7778 = n7571 | n7776;
  assign n7779 = ~n7777 & n7778;
  assign n7780 = x51 & x107;
  assign n7781 = n7779 & n7780;
  assign n7782 = n7779 | n7780;
  assign n7783 = ~n7781 & n7782;
  assign n7784 = n16384 & n7783;
  assign n7785 = n16384 | n7783;
  assign n7786 = ~n7784 & n7785;
  assign n7787 = x50 & x108;
  assign n7788 = n7786 & n7787;
  assign n7789 = n7786 | n7787;
  assign n7790 = ~n7788 & n7789;
  assign n7791 = n13331 & n7790;
  assign n7792 = n13331 | n7790;
  assign n7793 = ~n7791 & n7792;
  assign n7794 = x49 & x109;
  assign n7795 = n7793 & n7794;
  assign n7796 = n7793 | n7794;
  assign n7797 = ~n7795 & n7796;
  assign n7798 = n7566 & n7797;
  assign n7799 = n7566 | n7797;
  assign n7800 = ~n7798 & n7799;
  assign n7801 = x48 & x110;
  assign n7802 = n7800 & n7801;
  assign n7803 = n7800 | n7801;
  assign n7804 = ~n7802 & n7803;
  assign n17754 = n7565 | n7794;
  assign n17755 = (n7564 & n7794) | (n7564 & n17754) | (n7794 & n17754);
  assign n16460 = (n7566 & n7793) | (n7566 & n17755) | (n7793 & n17755);
  assign n13413 = (n7795 & n7797) | (n7795 & n16460) | (n7797 & n16460);
  assign n13414 = n7788 | n13331;
  assign n13415 = (n7788 & n7790) | (n7788 & n13414) | (n7790 & n13414);
  assign n16461 = n7781 | n16384;
  assign n16462 = (n7781 & n7783) | (n7781 & n16461) | (n7783 & n16461);
  assign n7808 = n7774 | n7777;
  assign n7809 = n7767 | n7770;
  assign n7810 = n7760 | n7763;
  assign n7811 = n7753 | n7756;
  assign n13416 = n7746 | n7748;
  assign n13417 = (n7575 & n7746) | (n7575 & n13416) | (n7746 & n13416);
  assign n13418 = n7739 | n7741;
  assign n13419 = (n7739 & n13333) | (n7739 & n13418) | (n13333 & n13418);
  assign n13420 = n7732 | n7734;
  assign n13421 = (n7732 & n13335) | (n7732 & n13420) | (n13335 & n13420);
  assign n13422 = n7725 | n7727;
  assign n13423 = (n7725 & n13337) | (n7725 & n13422) | (n13337 & n13422);
  assign n13424 = n7718 | n7720;
  assign n13425 = (n7718 & n13339) | (n7718 & n13424) | (n13339 & n13424);
  assign n13426 = n7711 | n7713;
  assign n13427 = (n7711 & n13341) | (n7711 & n13426) | (n13341 & n13426);
  assign n13345 = (n7468 & n13254) | (n7468 & n13344) | (n13254 & n13344);
  assign n13347 = (n7461 & n13256) | (n7461 & n13346) | (n13256 & n13346);
  assign n13437 = n7655 | n7657;
  assign n16463 = n7426 | n7655;
  assign n16464 = (n7655 & n7657) | (n7655 & n16463) | (n7657 & n16463);
  assign n16465 = (n13311 & n13437) | (n13311 & n16464) | (n13437 & n16464);
  assign n16466 = (n13310 & n13437) | (n13310 & n16464) | (n13437 & n16464);
  assign n16467 = (n16280 & n16465) | (n16280 & n16466) | (n16465 & n16466);
  assign n13272 = (n16240 & n16331) | (n16240 & n16333) | (n16331 & n16333);
  assign n7834 = x79 & x80;
  assign n7835 = x78 & x81;
  assign n7836 = n7834 & n7835;
  assign n7837 = n7834 | n7835;
  assign n7838 = ~n7836 & n7837;
  assign n13455 = n7599 | n7601;
  assign n13457 = n7838 & n13455;
  assign n13458 = n7599 & n7838;
  assign n17756 = (n7370 & n13457) | (n7370 & n13458) | (n13457 & n13458);
  assign n17757 = n13457 | n13458;
  assign n17758 = (n16342 & n17756) | (n16342 & n17757) | (n17756 & n17757);
  assign n17759 = (n13457 & n13458) | (n13457 & n16397) | (n13458 & n16397);
  assign n17760 = (n13457 & n13458) | (n13457 & n17740) | (n13458 & n17740);
  assign n17761 = (n16292 & n17759) | (n16292 & n17760) | (n17759 & n17760);
  assign n16472 = (n16133 & n17758) | (n16133 & n17761) | (n17758 & n17761);
  assign n13460 = n7838 | n13455;
  assign n13461 = n7599 | n7838;
  assign n17762 = (n7370 & n13460) | (n7370 & n13461) | (n13460 & n13461);
  assign n17763 = n13460 | n13461;
  assign n17764 = (n16342 & n17762) | (n16342 & n17763) | (n17762 & n17763);
  assign n17765 = (n13460 & n13461) | (n13460 & n16397) | (n13461 & n16397);
  assign n17766 = (n13460 & n13461) | (n13460 & n17740) | (n13461 & n17740);
  assign n17767 = (n16292 & n17765) | (n16292 & n17766) | (n17765 & n17766);
  assign n16475 = (n16133 & n17764) | (n16133 & n17767) | (n17764 & n17767);
  assign n7841 = ~n16472 & n16475;
  assign n7842 = x77 & x82;
  assign n7843 = n7841 & n7842;
  assign n7844 = n7841 | n7842;
  assign n7845 = ~n7843 & n7844;
  assign n16476 = n7606 | n7608;
  assign n16477 = (n7606 & n13363) | (n7606 & n16476) | (n13363 & n16476);
  assign n13463 = n7845 & n16477;
  assign n16478 = n7377 | n7606;
  assign n16479 = (n7606 & n7608) | (n7606 & n16478) | (n7608 & n16478);
  assign n13464 = n7845 & n16479;
  assign n16480 = (n13463 & n13464) | (n13463 & n16335) | (n13464 & n16335);
  assign n16481 = (n13463 & n13464) | (n13463 & n16336) | (n13464 & n16336);
  assign n16482 = (n16192 & n16480) | (n16192 & n16481) | (n16480 & n16481);
  assign n13466 = n7845 | n16477;
  assign n13467 = n7845 | n16479;
  assign n16483 = (n13466 & n13467) | (n13466 & n16335) | (n13467 & n16335);
  assign n16484 = (n13466 & n13467) | (n13466 & n16336) | (n13467 & n16336);
  assign n16485 = (n16192 & n16483) | (n16192 & n16484) | (n16483 & n16484);
  assign n7848 = ~n16482 & n16485;
  assign n7849 = x76 & x83;
  assign n7850 = n7848 & n7849;
  assign n7851 = n7848 | n7849;
  assign n7852 = ~n7850 & n7851;
  assign n16486 = n7384 | n7613;
  assign n16487 = (n7613 & n7615) | (n7613 & n16486) | (n7615 & n16486);
  assign n13469 = n7852 & n16487;
  assign n13450 = n7613 | n7615;
  assign n13470 = n7852 & n13450;
  assign n16488 = (n13288 & n13469) | (n13288 & n13470) | (n13469 & n13470);
  assign n16489 = (n13289 & n13469) | (n13289 & n13470) | (n13469 & n13470);
  assign n16490 = (n16243 & n16488) | (n16243 & n16489) | (n16488 & n16489);
  assign n13472 = n7852 | n16487;
  assign n13473 = n7852 | n13450;
  assign n16491 = (n13288 & n13472) | (n13288 & n13473) | (n13472 & n13473);
  assign n16492 = (n13289 & n13472) | (n13289 & n13473) | (n13472 & n13473);
  assign n16493 = (n16243 & n16491) | (n16243 & n16492) | (n16491 & n16492);
  assign n7855 = ~n16490 & n16493;
  assign n7856 = x75 & x84;
  assign n7857 = n7855 & n7856;
  assign n7858 = n7855 | n7856;
  assign n7859 = ~n7857 & n7858;
  assign n16494 = n7620 | n7622;
  assign n16495 = (n7620 & n13361) | (n7620 & n16494) | (n13361 & n16494);
  assign n13475 = n7859 & n16495;
  assign n16496 = n7391 | n7620;
  assign n16497 = (n7620 & n7622) | (n7620 & n16496) | (n7622 & n16496);
  assign n13476 = n7859 & n16497;
  assign n13477 = (n13272 & n13475) | (n13272 & n13476) | (n13475 & n13476);
  assign n13478 = n7859 | n16495;
  assign n13479 = n7859 | n16497;
  assign n13480 = (n13272 & n13478) | (n13272 & n13479) | (n13478 & n13479);
  assign n7862 = ~n13477 & n13480;
  assign n7863 = x74 & x85;
  assign n7864 = n7862 & n7863;
  assign n7865 = n7862 | n7863;
  assign n7866 = ~n7864 & n7865;
  assign n13444 = n7627 | n7629;
  assign n13481 = n7866 & n13444;
  assign n13482 = n7627 & n7866;
  assign n16498 = (n13481 & n13482) | (n13481 & n16395) | (n13482 & n16395);
  assign n16499 = (n13481 & n13482) | (n13481 & n16393) | (n13482 & n16393);
  assign n16500 = (n13174 & n16498) | (n13174 & n16499) | (n16498 & n16499);
  assign n13484 = n7866 | n13444;
  assign n13485 = n7627 | n7866;
  assign n16501 = (n13484 & n13485) | (n13484 & n16395) | (n13485 & n16395);
  assign n16502 = (n13484 & n13485) | (n13484 & n16393) | (n13485 & n16393);
  assign n16503 = (n13174 & n16501) | (n13174 & n16502) | (n16501 & n16502);
  assign n7869 = ~n16500 & n16503;
  assign n7870 = x73 & x86;
  assign n7871 = n7869 & n7870;
  assign n7872 = n7869 | n7870;
  assign n7873 = ~n7871 & n7872;
  assign n13442 = n7634 | n7636;
  assign n16504 = n7873 & n13442;
  assign n16468 = n7405 | n7634;
  assign n16469 = (n7634 & n7636) | (n7634 & n16468) | (n7636 & n16468);
  assign n16505 = n7873 & n16469;
  assign n16506 = (n13302 & n16504) | (n13302 & n16505) | (n16504 & n16505);
  assign n16507 = n7873 | n13442;
  assign n16508 = n7873 | n16469;
  assign n16509 = (n13302 & n16507) | (n13302 & n16508) | (n16507 & n16508);
  assign n7876 = ~n16506 & n16509;
  assign n7877 = x72 & x87;
  assign n7878 = n7876 & n7877;
  assign n7879 = n7876 | n7877;
  assign n7880 = ~n7878 & n7879;
  assign n13439 = n7641 | n7643;
  assign n13487 = n7880 & n13439;
  assign n13488 = n7641 & n7880;
  assign n13489 = (n16391 & n13487) | (n16391 & n13488) | (n13487 & n13488);
  assign n13490 = n7880 | n13439;
  assign n13491 = n7641 | n7880;
  assign n13492 = (n16391 & n13490) | (n16391 & n13491) | (n13490 & n13491);
  assign n7883 = ~n13489 & n13492;
  assign n7884 = x71 & x88;
  assign n7885 = n7883 & n7884;
  assign n7886 = n7883 | n7884;
  assign n7887 = ~n7885 & n7886;
  assign n13493 = n7648 & n7887;
  assign n16510 = (n7887 & n13389) | (n7887 & n13493) | (n13389 & n13493);
  assign n16511 = (n7887 & n13388) | (n7887 & n13493) | (n13388 & n13493);
  assign n16512 = (n16329 & n16510) | (n16329 & n16511) | (n16510 & n16511);
  assign n13495 = n7648 | n7887;
  assign n16513 = n13389 | n13495;
  assign n16514 = n13388 | n13495;
  assign n16515 = (n16329 & n16513) | (n16329 & n16514) | (n16513 & n16514);
  assign n7890 = ~n16512 & n16515;
  assign n7891 = x70 & x89;
  assign n7892 = n7890 & n7891;
  assign n7893 = n7890 | n7891;
  assign n7894 = ~n7892 & n7893;
  assign n7895 = n16467 & n7894;
  assign n7896 = n16467 | n7894;
  assign n7897 = ~n7895 & n7896;
  assign n7898 = x69 & x90;
  assign n7899 = n7897 & n7898;
  assign n7900 = n7897 | n7898;
  assign n7901 = ~n7899 & n7900;
  assign n13434 = n7662 | n7664;
  assign n13497 = n7901 & n13434;
  assign n13498 = n7662 & n7901;
  assign n16516 = (n13351 & n13497) | (n13351 & n13498) | (n13497 & n13498);
  assign n16517 = (n13497 & n13498) | (n13497 & n16386) | (n13498 & n16386);
  assign n16518 = (n16309 & n16516) | (n16309 & n16517) | (n16516 & n16517);
  assign n13500 = n7901 | n13434;
  assign n13501 = n7662 | n7901;
  assign n16519 = (n13351 & n13500) | (n13351 & n13501) | (n13500 & n13501);
  assign n16520 = (n13500 & n13501) | (n13500 & n16386) | (n13501 & n16386);
  assign n16521 = (n16309 & n16519) | (n16309 & n16520) | (n16519 & n16520);
  assign n7904 = ~n16518 & n16521;
  assign n7905 = x68 & x91;
  assign n7906 = n7904 & n7905;
  assign n7907 = n7904 | n7905;
  assign n7908 = ~n7906 & n7907;
  assign n13503 = n7669 & n7908;
  assign n13504 = (n7908 & n16443) | (n7908 & n13503) | (n16443 & n13503);
  assign n13505 = n7669 | n7908;
  assign n13506 = n16443 | n13505;
  assign n7911 = ~n13504 & n13506;
  assign n7912 = x67 & x92;
  assign n7913 = n7911 & n7912;
  assign n7914 = n7911 | n7912;
  assign n7915 = ~n7913 & n7914;
  assign n13507 = n7676 & n7915;
  assign n13508 = (n7915 & n13403) | (n7915 & n13507) | (n13403 & n13507);
  assign n13509 = n7676 | n7915;
  assign n13510 = n13403 | n13509;
  assign n7918 = ~n13508 & n13510;
  assign n7919 = x66 & x93;
  assign n7920 = n7918 & n7919;
  assign n7921 = n7918 | n7919;
  assign n7922 = ~n7920 & n7921;
  assign n13511 = n7683 & n7922;
  assign n13512 = (n7922 & n13408) | (n7922 & n13511) | (n13408 & n13511);
  assign n13513 = n7683 | n7922;
  assign n13514 = n13408 | n13513;
  assign n7925 = ~n13512 & n13514;
  assign n7926 = x65 & x94;
  assign n7927 = n7925 & n7926;
  assign n7928 = n7925 | n7926;
  assign n7929 = ~n7927 & n7928;
  assign n13432 = n7690 | n7692;
  assign n13515 = n7929 & n13432;
  assign n13516 = n7690 & n7929;
  assign n13517 = (n13347 & n13515) | (n13347 & n13516) | (n13515 & n13516);
  assign n13518 = n7929 | n13432;
  assign n13519 = n7690 | n7929;
  assign n13520 = (n13347 & n13518) | (n13347 & n13519) | (n13518 & n13519);
  assign n7932 = ~n13517 & n13520;
  assign n7933 = x64 & x95;
  assign n7934 = n7932 & n7933;
  assign n7935 = n7932 | n7933;
  assign n7936 = ~n7934 & n7935;
  assign n13430 = n7697 | n7699;
  assign n16522 = n7936 & n13430;
  assign n16523 = n7697 & n7936;
  assign n16524 = (n13345 & n16522) | (n13345 & n16523) | (n16522 & n16523);
  assign n16525 = n7936 | n13430;
  assign n16526 = n7697 | n7936;
  assign n16527 = (n13345 & n16525) | (n13345 & n16526) | (n16525 & n16526);
  assign n7939 = ~n16524 & n16527;
  assign n7940 = x63 & x96;
  assign n7941 = n7939 & n7940;
  assign n7942 = n7939 | n7940;
  assign n7943 = ~n7941 & n7942;
  assign n13428 = n7704 | n7706;
  assign n16528 = n7943 & n13428;
  assign n16529 = n7704 & n7943;
  assign n16530 = (n13343 & n16528) | (n13343 & n16529) | (n16528 & n16529);
  assign n16531 = n7943 | n13428;
  assign n16532 = n7704 | n7943;
  assign n16533 = (n13343 & n16531) | (n13343 & n16532) | (n16531 & n16532);
  assign n7946 = ~n16530 & n16533;
  assign n7947 = x62 & x97;
  assign n7948 = n7946 & n7947;
  assign n7949 = n7946 | n7947;
  assign n7950 = ~n7948 & n7949;
  assign n7951 = n13427 & n7950;
  assign n7952 = n13427 | n7950;
  assign n7953 = ~n7951 & n7952;
  assign n7954 = x61 & x98;
  assign n7955 = n7953 & n7954;
  assign n7956 = n7953 | n7954;
  assign n7957 = ~n7955 & n7956;
  assign n7958 = n13425 & n7957;
  assign n7959 = n13425 | n7957;
  assign n7960 = ~n7958 & n7959;
  assign n7961 = x60 & x99;
  assign n7962 = n7960 & n7961;
  assign n7963 = n7960 | n7961;
  assign n7964 = ~n7962 & n7963;
  assign n7965 = n13423 & n7964;
  assign n7966 = n13423 | n7964;
  assign n7967 = ~n7965 & n7966;
  assign n7968 = x59 & x100;
  assign n7969 = n7967 & n7968;
  assign n7970 = n7967 | n7968;
  assign n7971 = ~n7969 & n7970;
  assign n7972 = n13421 & n7971;
  assign n7973 = n13421 | n7971;
  assign n7974 = ~n7972 & n7973;
  assign n7975 = x58 & x101;
  assign n7976 = n7974 & n7975;
  assign n7977 = n7974 | n7975;
  assign n7978 = ~n7976 & n7977;
  assign n7979 = n13419 & n7978;
  assign n7980 = n13419 | n7978;
  assign n7981 = ~n7979 & n7980;
  assign n7982 = x57 & x102;
  assign n7983 = n7981 & n7982;
  assign n7984 = n7981 | n7982;
  assign n7985 = ~n7983 & n7984;
  assign n7986 = n13417 & n7985;
  assign n7987 = n13417 | n7985;
  assign n7988 = ~n7986 & n7987;
  assign n7989 = x56 & x103;
  assign n7990 = n7988 & n7989;
  assign n7991 = n7988 | n7989;
  assign n7992 = ~n7990 & n7991;
  assign n7993 = n7811 & n7992;
  assign n7994 = n7811 | n7992;
  assign n7995 = ~n7993 & n7994;
  assign n7996 = x55 & x104;
  assign n7997 = n7995 & n7996;
  assign n7998 = n7995 | n7996;
  assign n7999 = ~n7997 & n7998;
  assign n8000 = n7810 & n7999;
  assign n8001 = n7810 | n7999;
  assign n8002 = ~n8000 & n8001;
  assign n8003 = x54 & x105;
  assign n8004 = n8002 & n8003;
  assign n8005 = n8002 | n8003;
  assign n8006 = ~n8004 & n8005;
  assign n8007 = n7809 & n8006;
  assign n8008 = n7809 | n8006;
  assign n8009 = ~n8007 & n8008;
  assign n8010 = x53 & x106;
  assign n8011 = n8009 & n8010;
  assign n8012 = n8009 | n8010;
  assign n8013 = ~n8011 & n8012;
  assign n8014 = n7808 & n8013;
  assign n8015 = n7808 | n8013;
  assign n8016 = ~n8014 & n8015;
  assign n8017 = x52 & x107;
  assign n8018 = n8016 & n8017;
  assign n8019 = n8016 | n8017;
  assign n8020 = ~n8018 & n8019;
  assign n8021 = n16462 & n8020;
  assign n8022 = n16462 | n8020;
  assign n8023 = ~n8021 & n8022;
  assign n8024 = x51 & x108;
  assign n8025 = n8023 & n8024;
  assign n8026 = n8023 | n8024;
  assign n8027 = ~n8025 & n8026;
  assign n8028 = n13415 & n8027;
  assign n8029 = n13415 | n8027;
  assign n8030 = ~n8028 & n8029;
  assign n8031 = x50 & x109;
  assign n8032 = n8030 & n8031;
  assign n8033 = n8030 | n8031;
  assign n8034 = ~n8032 & n8033;
  assign n8035 = n13413 & n8034;
  assign n8036 = n13413 | n8034;
  assign n8037 = ~n8035 & n8036;
  assign n8038 = x49 & x110;
  assign n8039 = n8037 & n8038;
  assign n8040 = n8037 | n8038;
  assign n8041 = ~n8039 & n8040;
  assign n8042 = n7802 & n8041;
  assign n8043 = n7802 | n8041;
  assign n8044 = ~n8042 & n8043;
  assign n8045 = x48 & x111;
  assign n8046 = n8044 & n8045;
  assign n8047 = n8044 | n8045;
  assign n8048 = ~n8046 & n8047;
  assign n17768 = n7801 | n8038;
  assign n17769 = (n7800 & n8038) | (n7800 & n17768) | (n8038 & n17768);
  assign n16535 = (n7802 & n8037) | (n7802 & n17769) | (n8037 & n17769);
  assign n13522 = (n8039 & n8041) | (n8039 & n16535) | (n8041 & n16535);
  assign n13523 = n8032 | n13413;
  assign n13524 = (n8032 & n8034) | (n8032 & n13523) | (n8034 & n13523);
  assign n13525 = n8025 | n13415;
  assign n13526 = (n8025 & n8027) | (n8025 & n13525) | (n8027 & n13525);
  assign n16536 = n8018 | n16462;
  assign n16537 = (n8018 & n8020) | (n8018 & n16536) | (n8020 & n16536);
  assign n8053 = n8011 | n8014;
  assign n8054 = n8004 | n8007;
  assign n8055 = n7997 | n8000;
  assign n13527 = n7990 | n7992;
  assign n13528 = (n7811 & n7990) | (n7811 & n13527) | (n7990 & n13527);
  assign n13529 = n7983 | n7985;
  assign n13530 = (n7983 & n13417) | (n7983 & n13529) | (n13417 & n13529);
  assign n13531 = n7976 | n7978;
  assign n13532 = (n7976 & n13419) | (n7976 & n13531) | (n13419 & n13531);
  assign n13533 = n7969 | n7971;
  assign n13534 = (n7969 & n13421) | (n7969 & n13533) | (n13421 & n13533);
  assign n13535 = n7962 | n7964;
  assign n13536 = (n7962 & n13423) | (n7962 & n13535) | (n13423 & n13535);
  assign n13537 = n7955 | n7957;
  assign n13538 = (n7955 & n13425) | (n7955 & n13537) | (n13425 & n13537);
  assign n13429 = (n7704 & n13343) | (n7704 & n13428) | (n13343 & n13428);
  assign n13431 = (n7697 & n13345) | (n7697 & n13430) | (n13345 & n13430);
  assign n13551 = n7885 | n7887;
  assign n16540 = n7648 | n7885;
  assign n16541 = (n7885 & n7887) | (n7885 & n16540) | (n7887 & n16540);
  assign n16542 = (n13389 & n13551) | (n13389 & n16541) | (n13551 & n16541);
  assign n16543 = (n13388 & n13551) | (n13388 & n16541) | (n13551 & n16541);
  assign n16544 = (n16329 & n16542) | (n16329 & n16543) | (n16542 & n16543);
  assign n13360 = (n13174 & n16393) | (n13174 & n16395) | (n16393 & n16395);
  assign n16547 = n7850 | n7852;
  assign n16548 = (n7850 & n16487) | (n7850 & n16547) | (n16487 & n16547);
  assign n16549 = (n7850 & n13450) | (n7850 & n16547) | (n13450 & n16547);
  assign n16550 = (n13288 & n16548) | (n13288 & n16549) | (n16548 & n16549);
  assign n16551 = (n13289 & n16548) | (n13289 & n16549) | (n16548 & n16549);
  assign n16552 = (n16243 & n16550) | (n16243 & n16551) | (n16550 & n16551);
  assign n13366 = n7370 | n16342;
  assign n8079 = x79 & x81;
  assign n16553 = n7836 | n7838;
  assign n16554 = (n7836 & n13455) | (n7836 & n16553) | (n13455 & n16553);
  assign n13567 = n8079 & n16554;
  assign n16555 = n7599 | n7836;
  assign n16556 = (n7836 & n7838) | (n7836 & n16555) | (n7838 & n16555);
  assign n13568 = n8079 & n16556;
  assign n16557 = (n13366 & n13567) | (n13366 & n13568) | (n13567 & n13568);
  assign n16398 = (n16292 & n17740) | (n16292 & n16397) | (n17740 & n16397);
  assign n16558 = (n13567 & n13568) | (n13567 & n16398) | (n13568 & n16398);
  assign n16559 = (n16133 & n16557) | (n16133 & n16558) | (n16557 & n16558);
  assign n13570 = n8079 | n16554;
  assign n13571 = n8079 | n16556;
  assign n16560 = (n13366 & n13570) | (n13366 & n13571) | (n13570 & n13571);
  assign n16561 = (n13570 & n13571) | (n13570 & n16398) | (n13571 & n16398);
  assign n16562 = (n16133 & n16560) | (n16133 & n16561) | (n16560 & n16561);
  assign n8082 = ~n16559 & n16562;
  assign n8083 = x78 & x82;
  assign n8084 = n8082 & n8083;
  assign n8085 = n8082 | n8083;
  assign n8086 = ~n8084 & n8085;
  assign n16563 = n7843 | n7845;
  assign n16568 = (n7843 & n16479) | (n7843 & n16563) | (n16479 & n16563);
  assign n13574 = n8086 & n16568;
  assign n16565 = n8086 & n16563;
  assign n16566 = n7843 & n8086;
  assign n16567 = (n16477 & n16565) | (n16477 & n16566) | (n16565 & n16566);
  assign n16569 = (n13574 & n16335) | (n13574 & n16567) | (n16335 & n16567);
  assign n16570 = (n13574 & n16336) | (n13574 & n16567) | (n16336 & n16567);
  assign n16571 = (n16192 & n16569) | (n16192 & n16570) | (n16569 & n16570);
  assign n13577 = n8086 | n16568;
  assign n16572 = n8086 | n16563;
  assign n16573 = n7843 | n8086;
  assign n16574 = (n16477 & n16572) | (n16477 & n16573) | (n16572 & n16573);
  assign n16575 = (n13577 & n16335) | (n13577 & n16574) | (n16335 & n16574);
  assign n16576 = (n13577 & n16336) | (n13577 & n16574) | (n16336 & n16574);
  assign n16577 = (n16192 & n16575) | (n16192 & n16576) | (n16575 & n16576);
  assign n8089 = ~n16571 & n16577;
  assign n8090 = x77 & x83;
  assign n8091 = n8089 & n8090;
  assign n8092 = n8089 | n8090;
  assign n8093 = ~n8091 & n8092;
  assign n8094 = n16552 & n8093;
  assign n8095 = n16552 | n8093;
  assign n8096 = ~n8094 & n8095;
  assign n8097 = x76 & x84;
  assign n8098 = n8096 & n8097;
  assign n8099 = n8096 | n8097;
  assign n8100 = ~n8098 & n8099;
  assign n13579 = n7857 & n8100;
  assign n16578 = (n8100 & n13475) | (n8100 & n13579) | (n13475 & n13579);
  assign n16579 = (n8100 & n13476) | (n8100 & n13579) | (n13476 & n13579);
  assign n16580 = (n13272 & n16578) | (n13272 & n16579) | (n16578 & n16579);
  assign n13581 = n7857 | n8100;
  assign n16581 = n13475 | n13581;
  assign n16582 = n13476 | n13581;
  assign n16583 = (n13272 & n16581) | (n13272 & n16582) | (n16581 & n16582);
  assign n8103 = ~n16580 & n16583;
  assign n8104 = x75 & x85;
  assign n8105 = n8103 & n8104;
  assign n8106 = n8103 | n8104;
  assign n8107 = ~n8105 & n8106;
  assign n17770 = n7864 & n8107;
  assign n17771 = (n8107 & n13481) | (n8107 & n17770) | (n13481 & n17770);
  assign n16545 = n7627 | n7864;
  assign n16546 = (n7864 & n7866) | (n7864 & n16545) | (n7866 & n16545);
  assign n16585 = n8107 & n16546;
  assign n16586 = (n13360 & n17771) | (n13360 & n16585) | (n17771 & n16585);
  assign n17772 = n7864 | n8107;
  assign n17773 = n13481 | n17772;
  assign n16588 = n8107 | n16546;
  assign n16589 = (n13360 & n17773) | (n13360 & n16588) | (n17773 & n16588);
  assign n8110 = ~n16586 & n16589;
  assign n8111 = x74 & x86;
  assign n8112 = n8110 & n8111;
  assign n8113 = n8110 | n8111;
  assign n8114 = ~n8112 & n8113;
  assign n13553 = n7871 | n7873;
  assign n13583 = n8114 & n13553;
  assign n13584 = n7871 & n8114;
  assign n16590 = (n13442 & n13583) | (n13442 & n13584) | (n13583 & n13584);
  assign n16591 = (n13583 & n13584) | (n13583 & n16469) | (n13584 & n16469);
  assign n16592 = (n13302 & n16590) | (n13302 & n16591) | (n16590 & n16591);
  assign n13586 = n8114 | n13553;
  assign n13587 = n7871 | n8114;
  assign n16593 = (n13442 & n13586) | (n13442 & n13587) | (n13586 & n13587);
  assign n16594 = (n13586 & n13587) | (n13586 & n16469) | (n13587 & n16469);
  assign n16595 = (n13302 & n16593) | (n13302 & n16594) | (n16593 & n16594);
  assign n8117 = ~n16592 & n16595;
  assign n8118 = x73 & x87;
  assign n8119 = n8117 & n8118;
  assign n8120 = n8117 | n8118;
  assign n8121 = ~n8119 & n8120;
  assign n13589 = n7878 & n8121;
  assign n13590 = (n8121 & n13489) | (n8121 & n13589) | (n13489 & n13589);
  assign n13591 = n7878 | n8121;
  assign n13592 = n13489 | n13591;
  assign n8124 = ~n13590 & n13592;
  assign n8125 = x72 & x88;
  assign n8126 = n8124 & n8125;
  assign n8127 = n8124 | n8125;
  assign n8128 = ~n8126 & n8127;
  assign n8129 = n16544 & n8128;
  assign n8130 = n16544 | n8128;
  assign n8131 = ~n8129 & n8130;
  assign n8132 = x71 & x89;
  assign n8133 = n8131 & n8132;
  assign n8134 = n8131 | n8132;
  assign n8135 = ~n8133 & n8134;
  assign n13548 = n7892 | n7894;
  assign n13593 = n8135 & n13548;
  assign n13594 = n7892 & n8135;
  assign n13595 = (n16467 & n13593) | (n16467 & n13594) | (n13593 & n13594);
  assign n13596 = n8135 | n13548;
  assign n13597 = n7892 | n8135;
  assign n13598 = (n16467 & n13596) | (n16467 & n13597) | (n13596 & n13597);
  assign n8138 = ~n13595 & n13598;
  assign n8139 = x70 & x90;
  assign n8140 = n8138 & n8139;
  assign n8141 = n8138 | n8139;
  assign n8142 = ~n8140 & n8141;
  assign n13599 = n7899 & n8142;
  assign n13600 = (n8142 & n16518) | (n8142 & n13599) | (n16518 & n13599);
  assign n13601 = n7899 | n8142;
  assign n13602 = n16518 | n13601;
  assign n8145 = ~n13600 & n13602;
  assign n8146 = x69 & x91;
  assign n8147 = n8145 & n8146;
  assign n8148 = n8145 | n8146;
  assign n8149 = ~n8147 & n8148;
  assign n13546 = n7906 | n7908;
  assign n16596 = n8149 & n13546;
  assign n16538 = n7669 | n7906;
  assign n16539 = (n7906 & n7908) | (n7906 & n16538) | (n7908 & n16538);
  assign n16597 = n8149 & n16539;
  assign n16598 = (n16443 & n16596) | (n16443 & n16597) | (n16596 & n16597);
  assign n16599 = n8149 | n13546;
  assign n16600 = n8149 | n16539;
  assign n16601 = (n16443 & n16599) | (n16443 & n16600) | (n16599 & n16600);
  assign n8152 = ~n16598 & n16601;
  assign n8153 = x68 & x92;
  assign n8154 = n8152 & n8153;
  assign n8155 = n8152 | n8153;
  assign n8156 = ~n8154 & n8155;
  assign n13603 = n7913 & n8156;
  assign n16602 = (n8156 & n13507) | (n8156 & n13603) | (n13507 & n13603);
  assign n16603 = (n7915 & n8156) | (n7915 & n13603) | (n8156 & n13603);
  assign n16604 = (n13403 & n16602) | (n13403 & n16603) | (n16602 & n16603);
  assign n13605 = n7913 | n8156;
  assign n16605 = n13507 | n13605;
  assign n16606 = n7915 | n13605;
  assign n16607 = (n13403 & n16605) | (n13403 & n16606) | (n16605 & n16606);
  assign n8159 = ~n16604 & n16607;
  assign n8160 = x67 & x93;
  assign n8161 = n8159 & n8160;
  assign n8162 = n8159 | n8160;
  assign n8163 = ~n8161 & n8162;
  assign n13607 = n7920 & n8163;
  assign n13608 = (n8163 & n13512) | (n8163 & n13607) | (n13512 & n13607);
  assign n13609 = n7920 | n8163;
  assign n13610 = n13512 | n13609;
  assign n8166 = ~n13608 & n13610;
  assign n8167 = x66 & x94;
  assign n8168 = n8166 & n8167;
  assign n8169 = n8166 | n8167;
  assign n8170 = ~n8168 & n8169;
  assign n13611 = n7927 & n8170;
  assign n13612 = (n8170 & n13517) | (n8170 & n13611) | (n13517 & n13611);
  assign n13613 = n7927 | n8170;
  assign n13614 = n13517 | n13613;
  assign n8173 = ~n13612 & n13614;
  assign n8174 = x65 & x95;
  assign n8175 = n8173 & n8174;
  assign n8176 = n8173 | n8174;
  assign n8177 = ~n8175 & n8176;
  assign n13543 = n7934 | n7936;
  assign n13615 = n8177 & n13543;
  assign n13616 = n7934 & n8177;
  assign n13617 = (n13431 & n13615) | (n13431 & n13616) | (n13615 & n13616);
  assign n13618 = n8177 | n13543;
  assign n13619 = n7934 | n8177;
  assign n13620 = (n13431 & n13618) | (n13431 & n13619) | (n13618 & n13619);
  assign n8180 = ~n13617 & n13620;
  assign n8181 = x64 & x96;
  assign n8182 = n8180 & n8181;
  assign n8183 = n8180 | n8181;
  assign n8184 = ~n8182 & n8183;
  assign n13541 = n7941 | n7943;
  assign n16608 = n8184 & n13541;
  assign n16609 = n7941 & n8184;
  assign n16610 = (n13429 & n16608) | (n13429 & n16609) | (n16608 & n16609);
  assign n16611 = n8184 | n13541;
  assign n16612 = n7941 | n8184;
  assign n16613 = (n13429 & n16611) | (n13429 & n16612) | (n16611 & n16612);
  assign n8187 = ~n16610 & n16613;
  assign n8188 = x63 & x97;
  assign n8189 = n8187 & n8188;
  assign n8190 = n8187 | n8188;
  assign n8191 = ~n8189 & n8190;
  assign n13539 = n7948 | n7950;
  assign n16614 = n8191 & n13539;
  assign n16615 = n7948 & n8191;
  assign n16616 = (n13427 & n16614) | (n13427 & n16615) | (n16614 & n16615);
  assign n16617 = n8191 | n13539;
  assign n16618 = n7948 | n8191;
  assign n16619 = (n13427 & n16617) | (n13427 & n16618) | (n16617 & n16618);
  assign n8194 = ~n16616 & n16619;
  assign n8195 = x62 & x98;
  assign n8196 = n8194 & n8195;
  assign n8197 = n8194 | n8195;
  assign n8198 = ~n8196 & n8197;
  assign n8199 = n13538 & n8198;
  assign n8200 = n13538 | n8198;
  assign n8201 = ~n8199 & n8200;
  assign n8202 = x61 & x99;
  assign n8203 = n8201 & n8202;
  assign n8204 = n8201 | n8202;
  assign n8205 = ~n8203 & n8204;
  assign n8206 = n13536 & n8205;
  assign n8207 = n13536 | n8205;
  assign n8208 = ~n8206 & n8207;
  assign n8209 = x60 & x100;
  assign n8210 = n8208 & n8209;
  assign n8211 = n8208 | n8209;
  assign n8212 = ~n8210 & n8211;
  assign n8213 = n13534 & n8212;
  assign n8214 = n13534 | n8212;
  assign n8215 = ~n8213 & n8214;
  assign n8216 = x59 & x101;
  assign n8217 = n8215 & n8216;
  assign n8218 = n8215 | n8216;
  assign n8219 = ~n8217 & n8218;
  assign n8220 = n13532 & n8219;
  assign n8221 = n13532 | n8219;
  assign n8222 = ~n8220 & n8221;
  assign n8223 = x58 & x102;
  assign n8224 = n8222 & n8223;
  assign n8225 = n8222 | n8223;
  assign n8226 = ~n8224 & n8225;
  assign n8227 = n13530 & n8226;
  assign n8228 = n13530 | n8226;
  assign n8229 = ~n8227 & n8228;
  assign n8230 = x57 & x103;
  assign n8231 = n8229 & n8230;
  assign n8232 = n8229 | n8230;
  assign n8233 = ~n8231 & n8232;
  assign n8234 = n13528 & n8233;
  assign n8235 = n13528 | n8233;
  assign n8236 = ~n8234 & n8235;
  assign n8237 = x56 & x104;
  assign n8238 = n8236 & n8237;
  assign n8239 = n8236 | n8237;
  assign n8240 = ~n8238 & n8239;
  assign n8241 = n8055 & n8240;
  assign n8242 = n8055 | n8240;
  assign n8243 = ~n8241 & n8242;
  assign n8244 = x55 & x105;
  assign n8245 = n8243 & n8244;
  assign n8246 = n8243 | n8244;
  assign n8247 = ~n8245 & n8246;
  assign n8248 = n8054 & n8247;
  assign n8249 = n8054 | n8247;
  assign n8250 = ~n8248 & n8249;
  assign n8251 = x54 & x106;
  assign n8252 = n8250 & n8251;
  assign n8253 = n8250 | n8251;
  assign n8254 = ~n8252 & n8253;
  assign n8255 = n8053 & n8254;
  assign n8256 = n8053 | n8254;
  assign n8257 = ~n8255 & n8256;
  assign n8258 = x53 & x107;
  assign n8259 = n8257 & n8258;
  assign n8260 = n8257 | n8258;
  assign n8261 = ~n8259 & n8260;
  assign n8262 = n16537 & n8261;
  assign n8263 = n16537 | n8261;
  assign n8264 = ~n8262 & n8263;
  assign n8265 = x52 & x108;
  assign n8266 = n8264 & n8265;
  assign n8267 = n8264 | n8265;
  assign n8268 = ~n8266 & n8267;
  assign n8269 = n13526 & n8268;
  assign n8270 = n13526 | n8268;
  assign n8271 = ~n8269 & n8270;
  assign n8272 = x51 & x109;
  assign n8273 = n8271 & n8272;
  assign n8274 = n8271 | n8272;
  assign n8275 = ~n8273 & n8274;
  assign n8276 = n13524 & n8275;
  assign n8277 = n13524 | n8275;
  assign n8278 = ~n8276 & n8277;
  assign n8279 = x50 & x110;
  assign n8280 = n8278 & n8279;
  assign n8281 = n8278 | n8279;
  assign n8282 = ~n8280 & n8281;
  assign n8283 = n13522 & n8282;
  assign n8284 = n13522 | n8282;
  assign n8285 = ~n8283 & n8284;
  assign n8286 = x49 & x111;
  assign n8287 = n8285 & n8286;
  assign n8288 = n8285 | n8286;
  assign n8289 = ~n8287 & n8288;
  assign n8290 = n8046 & n8289;
  assign n8291 = n8046 | n8289;
  assign n8292 = ~n8290 & n8291;
  assign n17774 = n8045 | n8286;
  assign n17775 = (n8044 & n8286) | (n8044 & n17774) | (n8286 & n17774);
  assign n16621 = (n8046 & n8285) | (n8046 & n17775) | (n8285 & n17775);
  assign n13622 = (n8287 & n8289) | (n8287 & n16621) | (n8289 & n16621);
  assign n13623 = n8280 | n13522;
  assign n13624 = (n8280 & n8282) | (n8280 & n13623) | (n8282 & n13623);
  assign n13625 = n8273 | n13524;
  assign n13626 = (n8273 & n8275) | (n8273 & n13625) | (n8275 & n13625);
  assign n13627 = n8266 | n13526;
  assign n13628 = (n8266 & n8268) | (n8266 & n13627) | (n8268 & n13627);
  assign n16622 = n8259 | n16537;
  assign n16623 = (n8259 & n8261) | (n8259 & n16622) | (n8261 & n16622);
  assign n8298 = n8252 | n8255;
  assign n8299 = n8245 | n8248;
  assign n13629 = n8238 | n8240;
  assign n13630 = (n8055 & n8238) | (n8055 & n13629) | (n8238 & n13629);
  assign n13631 = n8231 | n8233;
  assign n13632 = (n8231 & n13528) | (n8231 & n13631) | (n13528 & n13631);
  assign n13633 = n8224 | n8226;
  assign n13634 = (n8224 & n13530) | (n8224 & n13633) | (n13530 & n13633);
  assign n13635 = n8217 | n8219;
  assign n13636 = (n8217 & n13532) | (n8217 & n13635) | (n13532 & n13635);
  assign n13637 = n8210 | n8212;
  assign n13638 = (n8210 & n13534) | (n8210 & n13637) | (n13534 & n13637);
  assign n13639 = n8203 | n8205;
  assign n13640 = (n8203 & n13536) | (n8203 & n13639) | (n13536 & n13639);
  assign n13540 = (n7948 & n13427) | (n7948 & n13539) | (n13427 & n13539);
  assign n13542 = (n7941 & n13429) | (n7941 & n13541) | (n13429 & n13541);
  assign n13547 = (n16443 & n16539) | (n16443 & n13546) | (n16539 & n13546);
  assign n13443 = (n13302 & n16469) | (n13302 & n13442) | (n16469 & n13442);
  assign n13555 = n7864 | n13481;
  assign n8323 = x79 & x82;
  assign n16630 = n8079 & n8323;
  assign n16631 = n16554 & n16630;
  assign n16632 = n16556 & n16630;
  assign n16633 = (n13366 & n16631) | (n13366 & n16632) | (n16631 & n16632);
  assign n16634 = (n16398 & n16631) | (n16398 & n16632) | (n16631 & n16632);
  assign n16635 = (n16133 & n16633) | (n16133 & n16634) | (n16633 & n16634);
  assign n16636 = n8079 | n8323;
  assign n16637 = (n8323 & n16554) | (n8323 & n16636) | (n16554 & n16636);
  assign n16638 = (n8323 & n16556) | (n8323 & n16636) | (n16556 & n16636);
  assign n16639 = (n13366 & n16637) | (n13366 & n16638) | (n16637 & n16638);
  assign n16640 = (n16398 & n16637) | (n16398 & n16638) | (n16637 & n16638);
  assign n16641 = (n16133 & n16639) | (n16133 & n16640) | (n16639 & n16640);
  assign n8326 = ~n16635 & n16641;
  assign n13673 = n8084 & n8326;
  assign n13674 = (n8326 & n16571) | (n8326 & n13673) | (n16571 & n13673);
  assign n13675 = n8084 | n8326;
  assign n13676 = n16571 | n13675;
  assign n8329 = ~n13674 & n13676;
  assign n8330 = x78 & x83;
  assign n8331 = n8329 & n8330;
  assign n8332 = n8329 | n8330;
  assign n8333 = ~n8331 & n8332;
  assign n13665 = n8091 | n8093;
  assign n13677 = n8333 & n13665;
  assign n13678 = n8091 & n8333;
  assign n13679 = (n16552 & n13677) | (n16552 & n13678) | (n13677 & n13678);
  assign n13680 = n8333 | n13665;
  assign n13681 = n8091 | n8333;
  assign n13682 = (n16552 & n13680) | (n16552 & n13681) | (n13680 & n13681);
  assign n8336 = ~n13679 & n13682;
  assign n8337 = x77 & x84;
  assign n8338 = n8336 & n8337;
  assign n8339 = n8336 | n8337;
  assign n8340 = ~n8338 & n8339;
  assign n16642 = n7857 | n8098;
  assign n16643 = (n8098 & n8100) | (n8098 & n16642) | (n8100 & n16642);
  assign n13683 = n8340 & n16643;
  assign n13663 = n8098 | n8100;
  assign n13684 = n8340 & n13663;
  assign n16644 = (n13475 & n13683) | (n13475 & n13684) | (n13683 & n13684);
  assign n16645 = (n13476 & n13683) | (n13476 & n13684) | (n13683 & n13684);
  assign n16646 = (n13272 & n16644) | (n13272 & n16645) | (n16644 & n16645);
  assign n13686 = n8340 | n16643;
  assign n13687 = n8340 | n13663;
  assign n16647 = (n13475 & n13686) | (n13475 & n13687) | (n13686 & n13687);
  assign n16648 = (n13476 & n13686) | (n13476 & n13687) | (n13686 & n13687);
  assign n16649 = (n13272 & n16647) | (n13272 & n16648) | (n16647 & n16648);
  assign n8343 = ~n16646 & n16649;
  assign n8344 = x76 & x85;
  assign n8345 = n8343 & n8344;
  assign n8346 = n8343 | n8344;
  assign n8347 = ~n8345 & n8346;
  assign n13660 = n8105 | n8107;
  assign n13689 = n8347 & n13660;
  assign n13690 = n8105 & n8347;
  assign n16650 = (n13555 & n13689) | (n13555 & n13690) | (n13689 & n13690);
  assign n16651 = (n13689 & n13690) | (n13689 & n16546) | (n13690 & n16546);
  assign n16652 = (n13360 & n16650) | (n13360 & n16651) | (n16650 & n16651);
  assign n13692 = n8347 | n13660;
  assign n13693 = n8105 | n8347;
  assign n16653 = (n13555 & n13692) | (n13555 & n13693) | (n13692 & n13693);
  assign n16654 = (n13692 & n13693) | (n13692 & n16546) | (n13693 & n16546);
  assign n16655 = (n13360 & n16653) | (n13360 & n16654) | (n16653 & n16654);
  assign n8350 = ~n16652 & n16655;
  assign n8351 = x75 & x86;
  assign n8352 = n8350 & n8351;
  assign n8353 = n8350 | n8351;
  assign n8354 = ~n8352 & n8353;
  assign n17776 = n8112 & n8354;
  assign n17777 = (n8354 & n13583) | (n8354 & n17776) | (n13583 & n17776);
  assign n16628 = n7871 | n8112;
  assign n16629 = (n8112 & n8114) | (n8112 & n16628) | (n8114 & n16628);
  assign n16657 = n8354 & n16629;
  assign n16658 = (n13443 & n17777) | (n13443 & n16657) | (n17777 & n16657);
  assign n17778 = n8112 | n8354;
  assign n17779 = n13583 | n17778;
  assign n16660 = n8354 | n16629;
  assign n16661 = (n13443 & n17779) | (n13443 & n16660) | (n17779 & n16660);
  assign n8357 = ~n16658 & n16661;
  assign n8358 = x74 & x87;
  assign n8359 = n8357 & n8358;
  assign n8360 = n8357 | n8358;
  assign n8361 = ~n8359 & n8360;
  assign n13655 = n8119 | n8121;
  assign n16662 = n8361 & n13655;
  assign n16626 = n7878 | n8119;
  assign n16627 = (n8119 & n8121) | (n8119 & n16626) | (n8121 & n16626);
  assign n16663 = n8361 & n16627;
  assign n16664 = (n13489 & n16662) | (n13489 & n16663) | (n16662 & n16663);
  assign n16665 = n8361 | n13655;
  assign n16666 = n8361 | n16627;
  assign n16667 = (n13489 & n16665) | (n13489 & n16666) | (n16665 & n16666);
  assign n8364 = ~n16664 & n16667;
  assign n8365 = x73 & x88;
  assign n8366 = n8364 & n8365;
  assign n8367 = n8364 | n8365;
  assign n8368 = ~n8366 & n8367;
  assign n13652 = n8126 | n8128;
  assign n13695 = n8368 & n13652;
  assign n13696 = n8126 & n8368;
  assign n13697 = (n16544 & n13695) | (n16544 & n13696) | (n13695 & n13696);
  assign n13698 = n8368 | n13652;
  assign n13699 = n8126 | n8368;
  assign n13700 = (n16544 & n13698) | (n16544 & n13699) | (n13698 & n13699);
  assign n8371 = ~n13697 & n13700;
  assign n8372 = x72 & x89;
  assign n8373 = n8371 & n8372;
  assign n8374 = n8371 | n8372;
  assign n8375 = ~n8373 & n8374;
  assign n13701 = n8133 & n8375;
  assign n16668 = (n8375 & n13594) | (n8375 & n13701) | (n13594 & n13701);
  assign n16669 = (n8375 & n13593) | (n8375 & n13701) | (n13593 & n13701);
  assign n16670 = (n16467 & n16668) | (n16467 & n16669) | (n16668 & n16669);
  assign n13703 = n8133 | n8375;
  assign n16671 = n13594 | n13703;
  assign n16672 = n13593 | n13703;
  assign n16673 = (n16467 & n16671) | (n16467 & n16672) | (n16671 & n16672);
  assign n8378 = ~n16670 & n16673;
  assign n8379 = x71 & x90;
  assign n8380 = n8378 & n8379;
  assign n8381 = n8378 | n8379;
  assign n8382 = ~n8380 & n8381;
  assign n13650 = n8140 | n8142;
  assign n16674 = n8382 & n13650;
  assign n16624 = n7899 | n8140;
  assign n16625 = (n8140 & n8142) | (n8140 & n16624) | (n8142 & n16624);
  assign n16675 = n8382 & n16625;
  assign n16676 = (n16518 & n16674) | (n16518 & n16675) | (n16674 & n16675);
  assign n16677 = n8382 | n13650;
  assign n16678 = n8382 | n16625;
  assign n16679 = (n16518 & n16677) | (n16518 & n16678) | (n16677 & n16678);
  assign n8385 = ~n16676 & n16679;
  assign n8386 = x70 & x91;
  assign n8387 = n8385 & n8386;
  assign n8388 = n8385 | n8386;
  assign n8389 = ~n8387 & n8388;
  assign n13647 = n8147 | n8149;
  assign n13705 = n8389 & n13647;
  assign n13706 = n8147 & n8389;
  assign n13707 = (n13547 & n13705) | (n13547 & n13706) | (n13705 & n13706);
  assign n13708 = n8389 | n13647;
  assign n13709 = n8147 | n8389;
  assign n13710 = (n13547 & n13708) | (n13547 & n13709) | (n13708 & n13709);
  assign n8392 = ~n13707 & n13710;
  assign n8393 = x69 & x92;
  assign n8394 = n8392 & n8393;
  assign n8395 = n8392 | n8393;
  assign n8396 = ~n8394 & n8395;
  assign n13711 = n8154 & n8396;
  assign n13712 = (n8396 & n16604) | (n8396 & n13711) | (n16604 & n13711);
  assign n13713 = n8154 | n8396;
  assign n13714 = n16604 | n13713;
  assign n8399 = ~n13712 & n13714;
  assign n8400 = x68 & x93;
  assign n8401 = n8399 & n8400;
  assign n8402 = n8399 | n8400;
  assign n8403 = ~n8401 & n8402;
  assign n13715 = n8161 & n8403;
  assign n13716 = (n8403 & n13608) | (n8403 & n13715) | (n13608 & n13715);
  assign n13717 = n8161 | n8403;
  assign n13718 = n13608 | n13717;
  assign n8406 = ~n13716 & n13718;
  assign n8407 = x67 & x94;
  assign n8408 = n8406 & n8407;
  assign n8409 = n8406 | n8407;
  assign n8410 = ~n8408 & n8409;
  assign n13719 = n8168 & n8410;
  assign n13720 = (n8410 & n13612) | (n8410 & n13719) | (n13612 & n13719);
  assign n13721 = n8168 | n8410;
  assign n13722 = n13612 | n13721;
  assign n8413 = ~n13720 & n13722;
  assign n8414 = x66 & x95;
  assign n8415 = n8413 & n8414;
  assign n8416 = n8413 | n8414;
  assign n8417 = ~n8415 & n8416;
  assign n13723 = n8175 & n8417;
  assign n13724 = (n8417 & n13617) | (n8417 & n13723) | (n13617 & n13723);
  assign n13725 = n8175 | n8417;
  assign n13726 = n13617 | n13725;
  assign n8420 = ~n13724 & n13726;
  assign n8421 = x65 & x96;
  assign n8422 = n8420 & n8421;
  assign n8423 = n8420 | n8421;
  assign n8424 = ~n8422 & n8423;
  assign n13645 = n8182 | n8184;
  assign n13727 = n8424 & n13645;
  assign n13728 = n8182 & n8424;
  assign n13729 = (n13542 & n13727) | (n13542 & n13728) | (n13727 & n13728);
  assign n13730 = n8424 | n13645;
  assign n13731 = n8182 | n8424;
  assign n13732 = (n13542 & n13730) | (n13542 & n13731) | (n13730 & n13731);
  assign n8427 = ~n13729 & n13732;
  assign n8428 = x64 & x97;
  assign n8429 = n8427 & n8428;
  assign n8430 = n8427 | n8428;
  assign n8431 = ~n8429 & n8430;
  assign n13643 = n8189 | n8191;
  assign n16680 = n8431 & n13643;
  assign n16681 = n8189 & n8431;
  assign n16682 = (n13540 & n16680) | (n13540 & n16681) | (n16680 & n16681);
  assign n16683 = n8431 | n13643;
  assign n16684 = n8189 | n8431;
  assign n16685 = (n13540 & n16683) | (n13540 & n16684) | (n16683 & n16684);
  assign n8434 = ~n16682 & n16685;
  assign n8435 = x63 & x98;
  assign n8436 = n8434 & n8435;
  assign n8437 = n8434 | n8435;
  assign n8438 = ~n8436 & n8437;
  assign n13641 = n8196 | n8198;
  assign n16686 = n8438 & n13641;
  assign n16687 = n8196 & n8438;
  assign n16688 = (n13538 & n16686) | (n13538 & n16687) | (n16686 & n16687);
  assign n16689 = n8438 | n13641;
  assign n16690 = n8196 | n8438;
  assign n16691 = (n13538 & n16689) | (n13538 & n16690) | (n16689 & n16690);
  assign n8441 = ~n16688 & n16691;
  assign n8442 = x62 & x99;
  assign n8443 = n8441 & n8442;
  assign n8444 = n8441 | n8442;
  assign n8445 = ~n8443 & n8444;
  assign n8446 = n13640 & n8445;
  assign n8447 = n13640 | n8445;
  assign n8448 = ~n8446 & n8447;
  assign n8449 = x61 & x100;
  assign n8450 = n8448 & n8449;
  assign n8451 = n8448 | n8449;
  assign n8452 = ~n8450 & n8451;
  assign n8453 = n13638 & n8452;
  assign n8454 = n13638 | n8452;
  assign n8455 = ~n8453 & n8454;
  assign n8456 = x60 & x101;
  assign n8457 = n8455 & n8456;
  assign n8458 = n8455 | n8456;
  assign n8459 = ~n8457 & n8458;
  assign n8460 = n13636 & n8459;
  assign n8461 = n13636 | n8459;
  assign n8462 = ~n8460 & n8461;
  assign n8463 = x59 & x102;
  assign n8464 = n8462 & n8463;
  assign n8465 = n8462 | n8463;
  assign n8466 = ~n8464 & n8465;
  assign n8467 = n13634 & n8466;
  assign n8468 = n13634 | n8466;
  assign n8469 = ~n8467 & n8468;
  assign n8470 = x58 & x103;
  assign n8471 = n8469 & n8470;
  assign n8472 = n8469 | n8470;
  assign n8473 = ~n8471 & n8472;
  assign n8474 = n13632 & n8473;
  assign n8475 = n13632 | n8473;
  assign n8476 = ~n8474 & n8475;
  assign n8477 = x57 & x104;
  assign n8478 = n8476 & n8477;
  assign n8479 = n8476 | n8477;
  assign n8480 = ~n8478 & n8479;
  assign n8481 = n13630 & n8480;
  assign n8482 = n13630 | n8480;
  assign n8483 = ~n8481 & n8482;
  assign n8484 = x56 & x105;
  assign n8485 = n8483 & n8484;
  assign n8486 = n8483 | n8484;
  assign n8487 = ~n8485 & n8486;
  assign n8488 = n8299 & n8487;
  assign n8489 = n8299 | n8487;
  assign n8490 = ~n8488 & n8489;
  assign n8491 = x55 & x106;
  assign n8492 = n8490 & n8491;
  assign n8493 = n8490 | n8491;
  assign n8494 = ~n8492 & n8493;
  assign n8495 = n8298 & n8494;
  assign n8496 = n8298 | n8494;
  assign n8497 = ~n8495 & n8496;
  assign n8498 = x54 & x107;
  assign n8499 = n8497 & n8498;
  assign n8500 = n8497 | n8498;
  assign n8501 = ~n8499 & n8500;
  assign n8502 = n16623 & n8501;
  assign n8503 = n16623 | n8501;
  assign n8504 = ~n8502 & n8503;
  assign n8505 = x53 & x108;
  assign n8506 = n8504 & n8505;
  assign n8507 = n8504 | n8505;
  assign n8508 = ~n8506 & n8507;
  assign n8509 = n13628 & n8508;
  assign n8510 = n13628 | n8508;
  assign n8511 = ~n8509 & n8510;
  assign n8512 = x52 & x109;
  assign n8513 = n8511 & n8512;
  assign n8514 = n8511 | n8512;
  assign n8515 = ~n8513 & n8514;
  assign n8516 = n13626 & n8515;
  assign n8517 = n13626 | n8515;
  assign n8518 = ~n8516 & n8517;
  assign n8519 = x51 & x110;
  assign n8520 = n8518 & n8519;
  assign n8521 = n8518 | n8519;
  assign n8522 = ~n8520 & n8521;
  assign n8523 = n13624 & n8522;
  assign n8524 = n13624 | n8522;
  assign n8525 = ~n8523 & n8524;
  assign n8526 = x50 & x111;
  assign n8527 = n8525 & n8526;
  assign n8528 = n8525 | n8526;
  assign n8529 = ~n8527 & n8528;
  assign n8530 = n13622 & n8529;
  assign n8531 = n13622 | n8529;
  assign n8532 = ~n8530 & n8531;
  assign n13733 = n8527 | n13622;
  assign n13734 = (n8527 & n8529) | (n8527 & n13733) | (n8529 & n13733);
  assign n13735 = n8520 | n13624;
  assign n13736 = (n8520 & n8522) | (n8520 & n13735) | (n8522 & n13735);
  assign n13737 = n8513 | n13626;
  assign n13738 = (n8513 & n8515) | (n8513 & n13737) | (n8515 & n13737);
  assign n13739 = n8506 | n13628;
  assign n13740 = (n8506 & n8508) | (n8506 & n13739) | (n8508 & n13739);
  assign n16692 = n8499 | n16623;
  assign n16693 = (n8499 & n8501) | (n8499 & n16692) | (n8501 & n16692);
  assign n8538 = n8492 | n8495;
  assign n13741 = n8485 | n8487;
  assign n13742 = (n8299 & n8485) | (n8299 & n13741) | (n8485 & n13741);
  assign n13743 = n8478 | n8480;
  assign n13744 = (n8478 & n13630) | (n8478 & n13743) | (n13630 & n13743);
  assign n13745 = n8471 | n8473;
  assign n13746 = (n8471 & n13632) | (n8471 & n13745) | (n13632 & n13745);
  assign n13747 = n8464 | n8466;
  assign n13748 = (n8464 & n13634) | (n8464 & n13747) | (n13634 & n13747);
  assign n13749 = n8457 | n8459;
  assign n13750 = (n8457 & n13636) | (n8457 & n13749) | (n13636 & n13749);
  assign n13751 = n8450 | n8452;
  assign n13752 = (n8450 & n13638) | (n8450 & n13751) | (n13638 & n13751);
  assign n13642 = (n8196 & n13538) | (n8196 & n13641) | (n13538 & n13641);
  assign n13644 = (n8189 & n13540) | (n8189 & n13643) | (n13540 & n13643);
  assign n13765 = n8373 | n8375;
  assign n16696 = n8133 | n8373;
  assign n16697 = (n8373 & n8375) | (n8373 & n16696) | (n8375 & n16696);
  assign n16698 = (n13594 & n13765) | (n13594 & n16697) | (n13765 & n16697);
  assign n16699 = (n13593 & n13765) | (n13593 & n16697) | (n13765 & n16697);
  assign n16700 = (n16467 & n16698) | (n16467 & n16699) | (n16698 & n16699);
  assign n13656 = (n13489 & n16627) | (n13489 & n13655) | (n16627 & n13655);
  assign n13658 = n8112 | n13583;
  assign n16701 = n8345 | n8347;
  assign n16702 = (n8345 & n13660) | (n8345 & n16701) | (n13660 & n16701);
  assign n16703 = n8105 | n8345;
  assign n16704 = (n8345 & n8347) | (n8345 & n16703) | (n8347 & n16703);
  assign n16705 = (n13555 & n16702) | (n13555 & n16704) | (n16702 & n16704);
  assign n16706 = (n16546 & n16702) | (n16546 & n16704) | (n16702 & n16704);
  assign n16707 = (n13360 & n16705) | (n13360 & n16706) | (n16705 & n16706);
  assign n8563 = x79 & x83;
  assign n16708 = n8326 | n16635;
  assign n16709 = (n8084 & n16635) | (n8084 & n16708) | (n16635 & n16708);
  assign n13780 = n8563 & n16709;
  assign n18043 = n8563 & n16630;
  assign n18044 = n16554 & n18043;
  assign n18045 = n16556 & n18043;
  assign n17933 = (n16398 & n18044) | (n16398 & n18045) | (n18044 & n18045);
  assign n17934 = (n13366 & n18044) | (n13366 & n18045) | (n18044 & n18045);
  assign n17782 = (n16133 & n17933) | (n16133 & n17934) | (n17933 & n17934);
  assign n16711 = (n8326 & n8563) | (n8326 & n17782) | (n8563 & n17782);
  assign n13782 = (n16571 & n13780) | (n16571 & n16711) | (n13780 & n16711);
  assign n13783 = n8563 | n16709;
  assign n18046 = n8563 | n16630;
  assign n18047 = (n8563 & n16554) | (n8563 & n18046) | (n16554 & n18046);
  assign n18048 = (n8563 & n16556) | (n8563 & n18046) | (n16556 & n18046);
  assign n17937 = (n16398 & n18047) | (n16398 & n18048) | (n18047 & n18048);
  assign n17938 = (n13366 & n18047) | (n13366 & n18048) | (n18047 & n18048);
  assign n17785 = (n16133 & n17937) | (n16133 & n17938) | (n17937 & n17938);
  assign n16713 = n8326 | n17785;
  assign n13785 = (n16571 & n13783) | (n16571 & n16713) | (n13783 & n16713);
  assign n8566 = ~n13782 & n13785;
  assign n16714 = n8331 & n8566;
  assign n16715 = (n8566 & n13677) | (n8566 & n16714) | (n13677 & n16714);
  assign n16716 = n8091 | n8331;
  assign n16717 = (n8331 & n8333) | (n8331 & n16716) | (n8333 & n16716);
  assign n13787 = n8566 & n16717;
  assign n13788 = (n16552 & n16715) | (n16552 & n13787) | (n16715 & n13787);
  assign n16718 = n8331 | n8566;
  assign n16719 = n13677 | n16718;
  assign n13790 = n8566 | n16717;
  assign n13791 = (n16552 & n16719) | (n16552 & n13790) | (n16719 & n13790);
  assign n8569 = ~n13788 & n13791;
  assign n8570 = x78 & x84;
  assign n8571 = n8569 & n8570;
  assign n8572 = n8569 | n8570;
  assign n8573 = ~n8571 & n8572;
  assign n13792 = n8338 & n8573;
  assign n13793 = (n8573 & n16646) | (n8573 & n13792) | (n16646 & n13792);
  assign n13794 = n8338 | n8573;
  assign n13795 = n16646 | n13794;
  assign n8576 = ~n13793 & n13795;
  assign n8577 = x77 & x85;
  assign n8578 = n8576 & n8577;
  assign n8579 = n8576 | n8577;
  assign n8580 = ~n8578 & n8579;
  assign n8581 = n16707 & n8580;
  assign n8582 = n16707 | n8580;
  assign n8583 = ~n8581 & n8582;
  assign n8584 = x76 & x86;
  assign n8585 = n8583 & n8584;
  assign n8586 = n8583 | n8584;
  assign n8587 = ~n8585 & n8586;
  assign n13769 = n8352 | n8354;
  assign n13796 = n8587 & n13769;
  assign n13797 = n8352 & n8587;
  assign n16720 = (n13658 & n13796) | (n13658 & n13797) | (n13796 & n13797);
  assign n16721 = (n13796 & n13797) | (n13796 & n16629) | (n13797 & n16629);
  assign n16722 = (n13443 & n16720) | (n13443 & n16721) | (n16720 & n16721);
  assign n13799 = n8587 | n13769;
  assign n13800 = n8352 | n8587;
  assign n16723 = (n13658 & n13799) | (n13658 & n13800) | (n13799 & n13800);
  assign n16724 = (n13799 & n13800) | (n13799 & n16629) | (n13800 & n16629);
  assign n16725 = (n13443 & n16723) | (n13443 & n16724) | (n16723 & n16724);
  assign n8590 = ~n16722 & n16725;
  assign n8591 = x75 & x87;
  assign n8592 = n8590 & n8591;
  assign n8593 = n8590 | n8591;
  assign n8594 = ~n8592 & n8593;
  assign n13767 = n8359 | n8361;
  assign n13802 = n8594 & n13767;
  assign n13803 = n8359 & n8594;
  assign n13804 = (n13656 & n13802) | (n13656 & n13803) | (n13802 & n13803);
  assign n13805 = n8594 | n13767;
  assign n13806 = n8359 | n8594;
  assign n13807 = (n13656 & n13805) | (n13656 & n13806) | (n13805 & n13806);
  assign n8597 = ~n13804 & n13807;
  assign n8598 = x74 & x88;
  assign n8599 = n8597 & n8598;
  assign n8600 = n8597 | n8598;
  assign n8601 = ~n8599 & n8600;
  assign n13808 = n8366 & n8601;
  assign n13809 = (n8601 & n13697) | (n8601 & n13808) | (n13697 & n13808);
  assign n13810 = n8366 | n8601;
  assign n13811 = n13697 | n13810;
  assign n8604 = ~n13809 & n13811;
  assign n8605 = x73 & x89;
  assign n8606 = n8604 & n8605;
  assign n8607 = n8604 | n8605;
  assign n8608 = ~n8606 & n8607;
  assign n8609 = n16700 & n8608;
  assign n8610 = n16700 | n8608;
  assign n8611 = ~n8609 & n8610;
  assign n8612 = x72 & x90;
  assign n8613 = n8611 & n8612;
  assign n8614 = n8611 | n8612;
  assign n8615 = ~n8613 & n8614;
  assign n13762 = n8380 | n8382;
  assign n13812 = n8615 & n13762;
  assign n13813 = n8380 & n8615;
  assign n16726 = (n13650 & n13812) | (n13650 & n13813) | (n13812 & n13813);
  assign n16727 = (n13812 & n13813) | (n13812 & n16625) | (n13813 & n16625);
  assign n16728 = (n16518 & n16726) | (n16518 & n16727) | (n16726 & n16727);
  assign n13815 = n8615 | n13762;
  assign n13816 = n8380 | n8615;
  assign n16729 = (n13650 & n13815) | (n13650 & n13816) | (n13815 & n13816);
  assign n16730 = (n13815 & n13816) | (n13815 & n16625) | (n13816 & n16625);
  assign n16731 = (n16518 & n16729) | (n16518 & n16730) | (n16729 & n16730);
  assign n8618 = ~n16728 & n16731;
  assign n8619 = x71 & x91;
  assign n8620 = n8618 & n8619;
  assign n8621 = n8618 | n8619;
  assign n8622 = ~n8620 & n8621;
  assign n13818 = n8387 & n8622;
  assign n16732 = (n8622 & n13705) | (n8622 & n13818) | (n13705 & n13818);
  assign n16733 = (n8622 & n13706) | (n8622 & n13818) | (n13706 & n13818);
  assign n16734 = (n13547 & n16732) | (n13547 & n16733) | (n16732 & n16733);
  assign n13820 = n8387 | n8622;
  assign n16735 = n13705 | n13820;
  assign n16736 = n13706 | n13820;
  assign n16737 = (n13547 & n16735) | (n13547 & n16736) | (n16735 & n16736);
  assign n8625 = ~n16734 & n16737;
  assign n8626 = x70 & x92;
  assign n8627 = n8625 & n8626;
  assign n8628 = n8625 | n8626;
  assign n8629 = ~n8627 & n8628;
  assign n13760 = n8394 | n8396;
  assign n16738 = n8629 & n13760;
  assign n16694 = n8154 | n8394;
  assign n16695 = (n8394 & n8396) | (n8394 & n16694) | (n8396 & n16694);
  assign n16739 = n8629 & n16695;
  assign n16740 = (n16604 & n16738) | (n16604 & n16739) | (n16738 & n16739);
  assign n16741 = n8629 | n13760;
  assign n16742 = n8629 | n16695;
  assign n16743 = (n16604 & n16741) | (n16604 & n16742) | (n16741 & n16742);
  assign n8632 = ~n16740 & n16743;
  assign n8633 = x69 & x93;
  assign n8634 = n8632 & n8633;
  assign n8635 = n8632 | n8633;
  assign n8636 = ~n8634 & n8635;
  assign n13822 = n8401 & n8636;
  assign n16744 = (n8636 & n13715) | (n8636 & n13822) | (n13715 & n13822);
  assign n16745 = (n8403 & n8636) | (n8403 & n13822) | (n8636 & n13822);
  assign n16746 = (n13608 & n16744) | (n13608 & n16745) | (n16744 & n16745);
  assign n13824 = n8401 | n8636;
  assign n16747 = n13715 | n13824;
  assign n16748 = n8403 | n13824;
  assign n16749 = (n13608 & n16747) | (n13608 & n16748) | (n16747 & n16748);
  assign n8639 = ~n16746 & n16749;
  assign n8640 = x68 & x94;
  assign n8641 = n8639 & n8640;
  assign n8642 = n8639 | n8640;
  assign n8643 = ~n8641 & n8642;
  assign n13826 = n8408 & n8643;
  assign n13827 = (n8643 & n13720) | (n8643 & n13826) | (n13720 & n13826);
  assign n13828 = n8408 | n8643;
  assign n13829 = n13720 | n13828;
  assign n8646 = ~n13827 & n13829;
  assign n8647 = x67 & x95;
  assign n8648 = n8646 & n8647;
  assign n8649 = n8646 | n8647;
  assign n8650 = ~n8648 & n8649;
  assign n13830 = n8415 & n8650;
  assign n13831 = (n8650 & n13724) | (n8650 & n13830) | (n13724 & n13830);
  assign n13832 = n8415 | n8650;
  assign n13833 = n13724 | n13832;
  assign n8653 = ~n13831 & n13833;
  assign n8654 = x66 & x96;
  assign n8655 = n8653 & n8654;
  assign n8656 = n8653 | n8654;
  assign n8657 = ~n8655 & n8656;
  assign n13834 = n8422 & n8657;
  assign n13835 = (n8657 & n13729) | (n8657 & n13834) | (n13729 & n13834);
  assign n13836 = n8422 | n8657;
  assign n13837 = n13729 | n13836;
  assign n8660 = ~n13835 & n13837;
  assign n8661 = x65 & x97;
  assign n8662 = n8660 & n8661;
  assign n8663 = n8660 | n8661;
  assign n8664 = ~n8662 & n8663;
  assign n13757 = n8429 | n8431;
  assign n13838 = n8664 & n13757;
  assign n13839 = n8429 & n8664;
  assign n13840 = (n13644 & n13838) | (n13644 & n13839) | (n13838 & n13839);
  assign n13841 = n8664 | n13757;
  assign n13842 = n8429 | n8664;
  assign n13843 = (n13644 & n13841) | (n13644 & n13842) | (n13841 & n13842);
  assign n8667 = ~n13840 & n13843;
  assign n8668 = x64 & x98;
  assign n8669 = n8667 & n8668;
  assign n8670 = n8667 | n8668;
  assign n8671 = ~n8669 & n8670;
  assign n13755 = n8436 | n8438;
  assign n16750 = n8671 & n13755;
  assign n16751 = n8436 & n8671;
  assign n16752 = (n13642 & n16750) | (n13642 & n16751) | (n16750 & n16751);
  assign n16753 = n8671 | n13755;
  assign n16754 = n8436 | n8671;
  assign n16755 = (n13642 & n16753) | (n13642 & n16754) | (n16753 & n16754);
  assign n8674 = ~n16752 & n16755;
  assign n8675 = x63 & x99;
  assign n8676 = n8674 & n8675;
  assign n8677 = n8674 | n8675;
  assign n8678 = ~n8676 & n8677;
  assign n13753 = n8443 | n8445;
  assign n16756 = n8678 & n13753;
  assign n16757 = n8443 & n8678;
  assign n16758 = (n13640 & n16756) | (n13640 & n16757) | (n16756 & n16757);
  assign n16759 = n8678 | n13753;
  assign n16760 = n8443 | n8678;
  assign n16761 = (n13640 & n16759) | (n13640 & n16760) | (n16759 & n16760);
  assign n8681 = ~n16758 & n16761;
  assign n8682 = x62 & x100;
  assign n8683 = n8681 & n8682;
  assign n8684 = n8681 | n8682;
  assign n8685 = ~n8683 & n8684;
  assign n8686 = n13752 & n8685;
  assign n8687 = n13752 | n8685;
  assign n8688 = ~n8686 & n8687;
  assign n8689 = x61 & x101;
  assign n8690 = n8688 & n8689;
  assign n8691 = n8688 | n8689;
  assign n8692 = ~n8690 & n8691;
  assign n8693 = n13750 & n8692;
  assign n8694 = n13750 | n8692;
  assign n8695 = ~n8693 & n8694;
  assign n8696 = x60 & x102;
  assign n8697 = n8695 & n8696;
  assign n8698 = n8695 | n8696;
  assign n8699 = ~n8697 & n8698;
  assign n8700 = n13748 & n8699;
  assign n8701 = n13748 | n8699;
  assign n8702 = ~n8700 & n8701;
  assign n8703 = x59 & x103;
  assign n8704 = n8702 & n8703;
  assign n8705 = n8702 | n8703;
  assign n8706 = ~n8704 & n8705;
  assign n8707 = n13746 & n8706;
  assign n8708 = n13746 | n8706;
  assign n8709 = ~n8707 & n8708;
  assign n8710 = x58 & x104;
  assign n8711 = n8709 & n8710;
  assign n8712 = n8709 | n8710;
  assign n8713 = ~n8711 & n8712;
  assign n8714 = n13744 & n8713;
  assign n8715 = n13744 | n8713;
  assign n8716 = ~n8714 & n8715;
  assign n8717 = x57 & x105;
  assign n8718 = n8716 & n8717;
  assign n8719 = n8716 | n8717;
  assign n8720 = ~n8718 & n8719;
  assign n8721 = n13742 & n8720;
  assign n8722 = n13742 | n8720;
  assign n8723 = ~n8721 & n8722;
  assign n8724 = x56 & x106;
  assign n8725 = n8723 & n8724;
  assign n8726 = n8723 | n8724;
  assign n8727 = ~n8725 & n8726;
  assign n8728 = n8538 & n8727;
  assign n8729 = n8538 | n8727;
  assign n8730 = ~n8728 & n8729;
  assign n8731 = x55 & x107;
  assign n8732 = n8730 & n8731;
  assign n8733 = n8730 | n8731;
  assign n8734 = ~n8732 & n8733;
  assign n8735 = n16693 & n8734;
  assign n8736 = n16693 | n8734;
  assign n8737 = ~n8735 & n8736;
  assign n8738 = x54 & x108;
  assign n8739 = n8737 & n8738;
  assign n8740 = n8737 | n8738;
  assign n8741 = ~n8739 & n8740;
  assign n8742 = n13740 & n8741;
  assign n8743 = n13740 | n8741;
  assign n8744 = ~n8742 & n8743;
  assign n8745 = x53 & x109;
  assign n8746 = n8744 & n8745;
  assign n8747 = n8744 | n8745;
  assign n8748 = ~n8746 & n8747;
  assign n8749 = n13738 & n8748;
  assign n8750 = n13738 | n8748;
  assign n8751 = ~n8749 & n8750;
  assign n8752 = x52 & x110;
  assign n8753 = n8751 & n8752;
  assign n8754 = n8751 | n8752;
  assign n8755 = ~n8753 & n8754;
  assign n8756 = n13736 & n8755;
  assign n8757 = n13736 | n8755;
  assign n8758 = ~n8756 & n8757;
  assign n8759 = x51 & x111;
  assign n8760 = n8758 & n8759;
  assign n8761 = n8758 | n8759;
  assign n8762 = ~n8760 & n8761;
  assign n8763 = n13734 & n8762;
  assign n8764 = n13734 | n8762;
  assign n8765 = ~n8763 & n8764;
  assign n13844 = n8760 | n13734;
  assign n13845 = (n8760 & n8762) | (n8760 & n13844) | (n8762 & n13844);
  assign n13846 = n8753 | n13736;
  assign n13847 = (n8753 & n8755) | (n8753 & n13846) | (n8755 & n13846);
  assign n13848 = n8746 | n13738;
  assign n13849 = (n8746 & n8748) | (n8746 & n13848) | (n8748 & n13848);
  assign n13850 = n8739 | n13740;
  assign n13851 = (n8739 & n8741) | (n8739 & n13850) | (n8741 & n13850);
  assign n16762 = n8732 | n16693;
  assign n16763 = (n8732 & n8734) | (n8732 & n16762) | (n8734 & n16762);
  assign n13852 = n8725 | n8727;
  assign n13853 = (n8538 & n8725) | (n8538 & n13852) | (n8725 & n13852);
  assign n13854 = n8718 | n8720;
  assign n13855 = (n8718 & n13742) | (n8718 & n13854) | (n13742 & n13854);
  assign n13856 = n8711 | n8713;
  assign n13857 = (n8711 & n13744) | (n8711 & n13856) | (n13744 & n13856);
  assign n13858 = n8704 | n8706;
  assign n13859 = (n8704 & n13746) | (n8704 & n13858) | (n13746 & n13858);
  assign n13860 = n8697 | n8699;
  assign n13861 = (n8697 & n13748) | (n8697 & n13860) | (n13748 & n13860);
  assign n13862 = n8690 | n8692;
  assign n13863 = (n8690 & n13750) | (n8690 & n13862) | (n13750 & n13862);
  assign n13754 = (n8443 & n13640) | (n8443 & n13753) | (n13640 & n13753);
  assign n13756 = (n8436 & n13642) | (n8436 & n13755) | (n13642 & n13755);
  assign n13761 = (n16604 & n16695) | (n16604 & n13760) | (n16695 & n13760);
  assign n13873 = n8620 | n8622;
  assign n16764 = n8387 | n8620;
  assign n16765 = (n8620 & n8622) | (n8620 & n16764) | (n8622 & n16764);
  assign n16766 = (n13705 & n13873) | (n13705 & n16765) | (n13873 & n16765);
  assign n16767 = (n13706 & n13873) | (n13706 & n16765) | (n13873 & n16765);
  assign n16768 = (n13547 & n16766) | (n13547 & n16767) | (n16766 & n16767);
  assign n13659 = (n13443 & n16629) | (n13443 & n13658) | (n16629 & n13658);
  assign n8795 = x79 & x84;
  assign n16773 = n8566 | n13782;
  assign n17786 = (n8331 & n13782) | (n8331 & n16773) | (n13782 & n16773);
  assign n17787 = n8795 & n17786;
  assign n18049 = n8563 & n8795;
  assign n18050 = n16709 & n18049;
  assign n18243 = n16630 & n18049;
  assign n18222 = n16554 & n18243;
  assign n18223 = n16556 & n18243;
  assign n18187 = (n13366 & n18222) | (n13366 & n18223) | (n18222 & n18223);
  assign n18188 = (n16398 & n18222) | (n16398 & n18223) | (n18222 & n18223);
  assign n18136 = (n16133 & n18187) | (n16133 & n18188) | (n18187 & n18188);
  assign n18052 = (n8326 & n18049) | (n8326 & n18136) | (n18049 & n18136);
  assign n17942 = (n16571 & n18050) | (n16571 & n18052) | (n18050 & n18052);
  assign n17939 = (n8566 & n8795) | (n8566 & n17942) | (n8795 & n17942);
  assign n17789 = (n13677 & n17787) | (n13677 & n17939) | (n17787 & n17939);
  assign n17791 = (n16717 & n17939) | (n16717 & n17942) | (n17939 & n17942);
  assign n16779 = (n16552 & n17789) | (n16552 & n17791) | (n17789 & n17791);
  assign n17792 = n8795 | n17786;
  assign n18053 = n8563 | n8795;
  assign n18054 = (n8795 & n16709) | (n8795 & n18053) | (n16709 & n18053);
  assign n18244 = (n8795 & n16630) | (n8795 & n18053) | (n16630 & n18053);
  assign n18225 = (n8795 & n16554) | (n8795 & n18244) | (n16554 & n18244);
  assign n18226 = (n8795 & n16556) | (n8795 & n18244) | (n16556 & n18244);
  assign n18191 = (n13366 & n18225) | (n13366 & n18226) | (n18225 & n18226);
  assign n18192 = (n16398 & n18225) | (n16398 & n18226) | (n18225 & n18226);
  assign n18139 = (n16133 & n18191) | (n16133 & n18192) | (n18191 & n18192);
  assign n18056 = (n8326 & n18053) | (n8326 & n18139) | (n18053 & n18139);
  assign n17946 = (n16571 & n18054) | (n16571 & n18056) | (n18054 & n18056);
  assign n17943 = n8566 | n17946;
  assign n17794 = (n13677 & n17792) | (n13677 & n17943) | (n17792 & n17943);
  assign n17796 = (n16717 & n17943) | (n16717 & n17946) | (n17943 & n17946);
  assign n16782 = (n16552 & n17794) | (n16552 & n17796) | (n17794 & n17796);
  assign n8798 = ~n16779 & n16782;
  assign n16783 = n8338 | n8571;
  assign n16784 = (n8571 & n8573) | (n8571 & n16783) | (n8573 & n16783);
  assign n13891 = n8798 & n16784;
  assign n16785 = n8571 & n8798;
  assign n16786 = (n8573 & n8798) | (n8573 & n16785) | (n8798 & n16785);
  assign n13893 = (n16646 & n13891) | (n16646 & n16786) | (n13891 & n16786);
  assign n13894 = n8798 | n16784;
  assign n16787 = n8571 | n8798;
  assign n16788 = n8573 | n16787;
  assign n13896 = (n16646 & n13894) | (n16646 & n16788) | (n13894 & n16788);
  assign n8801 = ~n13893 & n13896;
  assign n8802 = x78 & x85;
  assign n8803 = n8801 & n8802;
  assign n8804 = n8801 | n8802;
  assign n8805 = ~n8803 & n8804;
  assign n13883 = n8578 | n8580;
  assign n13897 = n8805 & n13883;
  assign n13898 = n8578 & n8805;
  assign n13899 = (n16707 & n13897) | (n16707 & n13898) | (n13897 & n13898);
  assign n13900 = n8805 | n13883;
  assign n13901 = n8578 | n8805;
  assign n13902 = (n16707 & n13900) | (n16707 & n13901) | (n13900 & n13901);
  assign n8808 = ~n13899 & n13902;
  assign n8809 = x77 & x86;
  assign n8810 = n8808 & n8809;
  assign n8811 = n8808 | n8809;
  assign n8812 = ~n8810 & n8811;
  assign n17797 = n8585 & n8812;
  assign n17798 = (n8812 & n13796) | (n8812 & n17797) | (n13796 & n17797);
  assign n16771 = n8352 | n8585;
  assign n16772 = (n8585 & n8587) | (n8585 & n16771) | (n8587 & n16771);
  assign n16790 = n8812 & n16772;
  assign n16791 = (n13659 & n17798) | (n13659 & n16790) | (n17798 & n16790);
  assign n17799 = n8585 | n8812;
  assign n17800 = n13796 | n17799;
  assign n16793 = n8812 | n16772;
  assign n16794 = (n13659 & n17800) | (n13659 & n16793) | (n17800 & n16793);
  assign n8815 = ~n16791 & n16794;
  assign n8816 = x76 & x87;
  assign n8817 = n8815 & n8816;
  assign n8818 = n8815 | n8816;
  assign n8819 = ~n8817 & n8818;
  assign n13903 = n8592 & n8819;
  assign n16795 = (n8819 & n13802) | (n8819 & n13903) | (n13802 & n13903);
  assign n16796 = (n8819 & n13803) | (n8819 & n13903) | (n13803 & n13903);
  assign n16797 = (n13656 & n16795) | (n13656 & n16796) | (n16795 & n16796);
  assign n13905 = n8592 | n8819;
  assign n16798 = n13802 | n13905;
  assign n16799 = n13803 | n13905;
  assign n16800 = (n13656 & n16798) | (n13656 & n16799) | (n16798 & n16799);
  assign n8822 = ~n16797 & n16800;
  assign n8823 = x75 & x88;
  assign n8824 = n8822 & n8823;
  assign n8825 = n8822 | n8823;
  assign n8826 = ~n8824 & n8825;
  assign n13878 = n8599 | n8601;
  assign n16801 = n8826 & n13878;
  assign n16769 = n8366 | n8599;
  assign n16770 = (n8599 & n8601) | (n8599 & n16769) | (n8601 & n16769);
  assign n16802 = n8826 & n16770;
  assign n16803 = (n13697 & n16801) | (n13697 & n16802) | (n16801 & n16802);
  assign n16804 = n8826 | n13878;
  assign n16805 = n8826 | n16770;
  assign n16806 = (n13697 & n16804) | (n13697 & n16805) | (n16804 & n16805);
  assign n8829 = ~n16803 & n16806;
  assign n8830 = x74 & x89;
  assign n8831 = n8829 & n8830;
  assign n8832 = n8829 | n8830;
  assign n8833 = ~n8831 & n8832;
  assign n13875 = n8606 | n8608;
  assign n13907 = n8833 & n13875;
  assign n13908 = n8606 & n8833;
  assign n13909 = (n16700 & n13907) | (n16700 & n13908) | (n13907 & n13908);
  assign n13910 = n8833 | n13875;
  assign n13911 = n8606 | n8833;
  assign n13912 = (n16700 & n13910) | (n16700 & n13911) | (n13910 & n13911);
  assign n8836 = ~n13909 & n13912;
  assign n8837 = x73 & x90;
  assign n8838 = n8836 & n8837;
  assign n8839 = n8836 | n8837;
  assign n8840 = ~n8838 & n8839;
  assign n13913 = n8613 & n8840;
  assign n13914 = (n8840 & n16728) | (n8840 & n13913) | (n16728 & n13913);
  assign n13915 = n8613 | n8840;
  assign n13916 = n16728 | n13915;
  assign n8843 = ~n13914 & n13916;
  assign n8844 = x72 & x91;
  assign n8845 = n8843 & n8844;
  assign n8846 = n8843 | n8844;
  assign n8847 = ~n8845 & n8846;
  assign n8848 = n16768 & n8847;
  assign n8849 = n16768 | n8847;
  assign n8850 = ~n8848 & n8849;
  assign n8851 = x71 & x92;
  assign n8852 = n8850 & n8851;
  assign n8853 = n8850 | n8851;
  assign n8854 = ~n8852 & n8853;
  assign n13870 = n8627 | n8629;
  assign n13917 = n8854 & n13870;
  assign n13918 = n8627 & n8854;
  assign n13919 = (n13761 & n13917) | (n13761 & n13918) | (n13917 & n13918);
  assign n13920 = n8854 | n13870;
  assign n13921 = n8627 | n8854;
  assign n13922 = (n13761 & n13920) | (n13761 & n13921) | (n13920 & n13921);
  assign n8857 = ~n13919 & n13922;
  assign n8858 = x70 & x93;
  assign n8859 = n8857 & n8858;
  assign n8860 = n8857 | n8858;
  assign n8861 = ~n8859 & n8860;
  assign n13923 = n8634 & n8861;
  assign n13924 = (n8861 & n16746) | (n8861 & n13923) | (n16746 & n13923);
  assign n13925 = n8634 | n8861;
  assign n13926 = n16746 | n13925;
  assign n8864 = ~n13924 & n13926;
  assign n8865 = x69 & x94;
  assign n8866 = n8864 & n8865;
  assign n8867 = n8864 | n8865;
  assign n8868 = ~n8866 & n8867;
  assign n13927 = n8641 & n8868;
  assign n13928 = (n8868 & n13827) | (n8868 & n13927) | (n13827 & n13927);
  assign n13929 = n8641 | n8868;
  assign n13930 = n13827 | n13929;
  assign n8871 = ~n13928 & n13930;
  assign n8872 = x68 & x95;
  assign n8873 = n8871 & n8872;
  assign n8874 = n8871 | n8872;
  assign n8875 = ~n8873 & n8874;
  assign n13931 = n8648 & n8875;
  assign n13932 = (n8875 & n13831) | (n8875 & n13931) | (n13831 & n13931);
  assign n13933 = n8648 | n8875;
  assign n13934 = n13831 | n13933;
  assign n8878 = ~n13932 & n13934;
  assign n8879 = x67 & x96;
  assign n8880 = n8878 & n8879;
  assign n8881 = n8878 | n8879;
  assign n8882 = ~n8880 & n8881;
  assign n13935 = n8655 & n8882;
  assign n13936 = (n8882 & n13835) | (n8882 & n13935) | (n13835 & n13935);
  assign n13937 = n8655 | n8882;
  assign n13938 = n13835 | n13937;
  assign n8885 = ~n13936 & n13938;
  assign n8886 = x66 & x97;
  assign n8887 = n8885 & n8886;
  assign n8888 = n8885 | n8886;
  assign n8889 = ~n8887 & n8888;
  assign n13939 = n8662 & n8889;
  assign n13940 = (n8889 & n13840) | (n8889 & n13939) | (n13840 & n13939);
  assign n13941 = n8662 | n8889;
  assign n13942 = n13840 | n13941;
  assign n8892 = ~n13940 & n13942;
  assign n8893 = x65 & x98;
  assign n8894 = n8892 & n8893;
  assign n8895 = n8892 | n8893;
  assign n8896 = ~n8894 & n8895;
  assign n13868 = n8669 | n8671;
  assign n13943 = n8896 & n13868;
  assign n13944 = n8669 & n8896;
  assign n13945 = (n13756 & n13943) | (n13756 & n13944) | (n13943 & n13944);
  assign n13946 = n8896 | n13868;
  assign n13947 = n8669 | n8896;
  assign n13948 = (n13756 & n13946) | (n13756 & n13947) | (n13946 & n13947);
  assign n8899 = ~n13945 & n13948;
  assign n8900 = x64 & x99;
  assign n8901 = n8899 & n8900;
  assign n8902 = n8899 | n8900;
  assign n8903 = ~n8901 & n8902;
  assign n13866 = n8676 | n8678;
  assign n16807 = n8903 & n13866;
  assign n16808 = n8676 & n8903;
  assign n16809 = (n13754 & n16807) | (n13754 & n16808) | (n16807 & n16808);
  assign n16810 = n8903 | n13866;
  assign n16811 = n8676 | n8903;
  assign n16812 = (n13754 & n16810) | (n13754 & n16811) | (n16810 & n16811);
  assign n8906 = ~n16809 & n16812;
  assign n8907 = x63 & x100;
  assign n8908 = n8906 & n8907;
  assign n8909 = n8906 | n8907;
  assign n8910 = ~n8908 & n8909;
  assign n13864 = n8683 | n8685;
  assign n16813 = n8910 & n13864;
  assign n16814 = n8683 & n8910;
  assign n16815 = (n13752 & n16813) | (n13752 & n16814) | (n16813 & n16814);
  assign n16816 = n8910 | n13864;
  assign n16817 = n8683 | n8910;
  assign n16818 = (n13752 & n16816) | (n13752 & n16817) | (n16816 & n16817);
  assign n8913 = ~n16815 & n16818;
  assign n8914 = x62 & x101;
  assign n8915 = n8913 & n8914;
  assign n8916 = n8913 | n8914;
  assign n8917 = ~n8915 & n8916;
  assign n8918 = n13863 & n8917;
  assign n8919 = n13863 | n8917;
  assign n8920 = ~n8918 & n8919;
  assign n8921 = x61 & x102;
  assign n8922 = n8920 & n8921;
  assign n8923 = n8920 | n8921;
  assign n8924 = ~n8922 & n8923;
  assign n8925 = n13861 & n8924;
  assign n8926 = n13861 | n8924;
  assign n8927 = ~n8925 & n8926;
  assign n8928 = x60 & x103;
  assign n8929 = n8927 & n8928;
  assign n8930 = n8927 | n8928;
  assign n8931 = ~n8929 & n8930;
  assign n8932 = n13859 & n8931;
  assign n8933 = n13859 | n8931;
  assign n8934 = ~n8932 & n8933;
  assign n8935 = x59 & x104;
  assign n8936 = n8934 & n8935;
  assign n8937 = n8934 | n8935;
  assign n8938 = ~n8936 & n8937;
  assign n8939 = n13857 & n8938;
  assign n8940 = n13857 | n8938;
  assign n8941 = ~n8939 & n8940;
  assign n8942 = x58 & x105;
  assign n8943 = n8941 & n8942;
  assign n8944 = n8941 | n8942;
  assign n8945 = ~n8943 & n8944;
  assign n8946 = n13855 & n8945;
  assign n8947 = n13855 | n8945;
  assign n8948 = ~n8946 & n8947;
  assign n8949 = x57 & x106;
  assign n8950 = n8948 & n8949;
  assign n8951 = n8948 | n8949;
  assign n8952 = ~n8950 & n8951;
  assign n8953 = n13853 & n8952;
  assign n8954 = n13853 | n8952;
  assign n8955 = ~n8953 & n8954;
  assign n8956 = x56 & x107;
  assign n8957 = n8955 & n8956;
  assign n8958 = n8955 | n8956;
  assign n8959 = ~n8957 & n8958;
  assign n8960 = n16763 & n8959;
  assign n8961 = n16763 | n8959;
  assign n8962 = ~n8960 & n8961;
  assign n8963 = x55 & x108;
  assign n8964 = n8962 & n8963;
  assign n8965 = n8962 | n8963;
  assign n8966 = ~n8964 & n8965;
  assign n8967 = n13851 & n8966;
  assign n8968 = n13851 | n8966;
  assign n8969 = ~n8967 & n8968;
  assign n8970 = x54 & x109;
  assign n8971 = n8969 & n8970;
  assign n8972 = n8969 | n8970;
  assign n8973 = ~n8971 & n8972;
  assign n8974 = n13849 & n8973;
  assign n8975 = n13849 | n8973;
  assign n8976 = ~n8974 & n8975;
  assign n8977 = x53 & x110;
  assign n8978 = n8976 & n8977;
  assign n8979 = n8976 | n8977;
  assign n8980 = ~n8978 & n8979;
  assign n8981 = n13847 & n8980;
  assign n8982 = n13847 | n8980;
  assign n8983 = ~n8981 & n8982;
  assign n8984 = x52 & x111;
  assign n8985 = n8983 & n8984;
  assign n8986 = n8983 | n8984;
  assign n8987 = ~n8985 & n8986;
  assign n8988 = n13845 & n8987;
  assign n8989 = n13845 | n8987;
  assign n8990 = ~n8988 & n8989;
  assign n13949 = n8985 | n13845;
  assign n13950 = (n8985 & n8987) | (n8985 & n13949) | (n8987 & n13949);
  assign n13951 = n8978 | n13847;
  assign n13952 = (n8978 & n8980) | (n8978 & n13951) | (n8980 & n13951);
  assign n13953 = n8971 | n13849;
  assign n13954 = (n8971 & n8973) | (n8971 & n13953) | (n8973 & n13953);
  assign n13955 = n8964 | n13851;
  assign n13956 = (n8964 & n8966) | (n8964 & n13955) | (n8966 & n13955);
  assign n13957 = n8957 | n8959;
  assign n13958 = (n16763 & n8957) | (n16763 & n13957) | (n8957 & n13957);
  assign n13959 = n8950 | n8952;
  assign n13960 = (n8950 & n13853) | (n8950 & n13959) | (n13853 & n13959);
  assign n13961 = n8943 | n8945;
  assign n13962 = (n8943 & n13855) | (n8943 & n13961) | (n13855 & n13961);
  assign n13963 = n8936 | n8938;
  assign n13964 = (n8936 & n13857) | (n8936 & n13963) | (n13857 & n13963);
  assign n13965 = n8929 | n8931;
  assign n13966 = (n8929 & n13859) | (n8929 & n13965) | (n13859 & n13965);
  assign n13967 = n8922 | n8924;
  assign n13968 = (n8922 & n13861) | (n8922 & n13967) | (n13861 & n13967);
  assign n13865 = (n8683 & n13752) | (n8683 & n13864) | (n13752 & n13864);
  assign n13867 = (n8676 & n13754) | (n8676 & n13866) | (n13754 & n13866);
  assign n13879 = (n13697 & n16770) | (n13697 & n13878) | (n16770 & n13878);
  assign n13986 = n8817 | n8819;
  assign n16823 = n8592 | n8817;
  assign n16824 = (n8817 & n8819) | (n8817 & n16823) | (n8819 & n16823);
  assign n16825 = (n13802 & n13986) | (n13802 & n16824) | (n13986 & n16824);
  assign n16826 = (n13803 & n13986) | (n13803 & n16824) | (n13986 & n16824);
  assign n16827 = (n13656 & n16825) | (n13656 & n16826) | (n16825 & n16826);
  assign n13881 = n8585 | n13796;
  assign n9019 = x79 & x85;
  assign n18193 = n9019 & n18049;
  assign n18194 = n16709 & n18193;
  assign n18259 = n9019 & n18243;
  assign n18260 = n16554 & n18259;
  assign n18261 = n16556 & n18259;
  assign n18247 = (n16398 & n18260) | (n16398 & n18261) | (n18260 & n18261);
  assign n18248 = (n13366 & n18260) | (n13366 & n18261) | (n18260 & n18261);
  assign n18229 = (n16133 & n18247) | (n16133 & n18248) | (n18247 & n18248);
  assign n18196 = (n8326 & n18193) | (n8326 & n18229) | (n18193 & n18229);
  assign n18144 = (n16571 & n18194) | (n16571 & n18196) | (n18194 & n18196);
  assign n18140 = n8795 & n9019;
  assign n18141 = (n8566 & n18144) | (n8566 & n18140) | (n18144 & n18140);
  assign n18059 = (n16717 & n18141) | (n16717 & n18144) | (n18141 & n18144);
  assign n17948 = n9019 & n17789;
  assign n17949 = (n16552 & n18059) | (n16552 & n17948) | (n18059 & n17948);
  assign n17802 = (n9019 & n16786) | (n9019 & n17949) | (n16786 & n17949);
  assign n17950 = (n8798 & n9019) | (n8798 & n17949) | (n9019 & n17949);
  assign n17804 = (n16784 & n17949) | (n16784 & n17950) | (n17949 & n17950);
  assign n16836 = (n16646 & n17802) | (n16646 & n17804) | (n17802 & n17804);
  assign n18197 = n9019 | n18049;
  assign n18198 = (n9019 & n16709) | (n9019 & n18197) | (n16709 & n18197);
  assign n18262 = n9019 | n18243;
  assign n18263 = (n9019 & n16554) | (n9019 & n18262) | (n16554 & n18262);
  assign n18264 = (n9019 & n16556) | (n9019 & n18262) | (n16556 & n18262);
  assign n18251 = (n16398 & n18263) | (n16398 & n18264) | (n18263 & n18264);
  assign n18252 = (n13366 & n18263) | (n13366 & n18264) | (n18263 & n18264);
  assign n18232 = (n16133 & n18251) | (n16133 & n18252) | (n18251 & n18252);
  assign n18200 = (n8326 & n18197) | (n8326 & n18232) | (n18197 & n18232);
  assign n18149 = (n16571 & n18198) | (n16571 & n18200) | (n18198 & n18200);
  assign n18145 = n8795 | n9019;
  assign n18146 = (n8566 & n18149) | (n8566 & n18145) | (n18149 & n18145);
  assign n18062 = (n16717 & n18146) | (n16717 & n18149) | (n18146 & n18149);
  assign n17952 = n9019 | n17789;
  assign n17953 = (n16552 & n18062) | (n16552 & n17952) | (n18062 & n17952);
  assign n17806 = n16786 | n17953;
  assign n17954 = n8798 | n17953;
  assign n17808 = (n16784 & n17953) | (n16784 & n17954) | (n17953 & n17954);
  assign n16839 = (n16646 & n17806) | (n16646 & n17808) | (n17806 & n17808);
  assign n9022 = ~n16836 & n16839;
  assign n16828 = n8803 | n8805;
  assign n16829 = (n8803 & n13883) | (n8803 & n16828) | (n13883 & n16828);
  assign n16840 = n9022 & n16829;
  assign n16830 = n8578 | n8803;
  assign n16831 = (n8803 & n8805) | (n8803 & n16830) | (n8805 & n16830);
  assign n16841 = n9022 & n16831;
  assign n16842 = (n16707 & n16840) | (n16707 & n16841) | (n16840 & n16841);
  assign n16843 = n9022 | n16829;
  assign n16844 = n9022 | n16831;
  assign n16845 = (n16707 & n16843) | (n16707 & n16844) | (n16843 & n16844);
  assign n9025 = ~n16842 & n16845;
  assign n9026 = x78 & x86;
  assign n9027 = n9025 & n9026;
  assign n9028 = n9025 | n9026;
  assign n9029 = ~n9027 & n9028;
  assign n13988 = n8810 | n8812;
  assign n13996 = n9029 & n13988;
  assign n13997 = n8810 & n9029;
  assign n16846 = (n13881 & n13996) | (n13881 & n13997) | (n13996 & n13997);
  assign n16847 = (n13996 & n13997) | (n13996 & n16772) | (n13997 & n16772);
  assign n16848 = (n13659 & n16846) | (n13659 & n16847) | (n16846 & n16847);
  assign n13999 = n9029 | n13988;
  assign n14000 = n8810 | n9029;
  assign n16849 = (n13881 & n13999) | (n13881 & n14000) | (n13999 & n14000);
  assign n16850 = (n13999 & n14000) | (n13999 & n16772) | (n14000 & n16772);
  assign n16851 = (n13659 & n16849) | (n13659 & n16850) | (n16849 & n16850);
  assign n9032 = ~n16848 & n16851;
  assign n9033 = x77 & x87;
  assign n9034 = n9032 & n9033;
  assign n9035 = n9032 | n9033;
  assign n9036 = ~n9034 & n9035;
  assign n9037 = n16827 & n9036;
  assign n9038 = n16827 | n9036;
  assign n9039 = ~n9037 & n9038;
  assign n9040 = x76 & x88;
  assign n9041 = n9039 & n9040;
  assign n9042 = n9039 | n9040;
  assign n9043 = ~n9041 & n9042;
  assign n13983 = n8824 | n8826;
  assign n14002 = n9043 & n13983;
  assign n14003 = n8824 & n9043;
  assign n14004 = (n13879 & n14002) | (n13879 & n14003) | (n14002 & n14003);
  assign n14005 = n9043 | n13983;
  assign n14006 = n8824 | n9043;
  assign n14007 = (n13879 & n14005) | (n13879 & n14006) | (n14005 & n14006);
  assign n9046 = ~n14004 & n14007;
  assign n9047 = x75 & x89;
  assign n9048 = n9046 & n9047;
  assign n9049 = n9046 | n9047;
  assign n9050 = ~n9048 & n9049;
  assign n14008 = n8831 & n9050;
  assign n14009 = (n9050 & n13909) | (n9050 & n14008) | (n13909 & n14008);
  assign n14010 = n8831 | n9050;
  assign n14011 = n13909 | n14010;
  assign n9053 = ~n14009 & n14011;
  assign n9054 = x74 & x90;
  assign n9055 = n9053 & n9054;
  assign n9056 = n9053 | n9054;
  assign n9057 = ~n9055 & n9056;
  assign n13981 = n8838 | n8840;
  assign n16852 = n9057 & n13981;
  assign n16821 = n8613 | n8838;
  assign n16822 = (n8838 & n8840) | (n8838 & n16821) | (n8840 & n16821);
  assign n16853 = n9057 & n16822;
  assign n16854 = (n16728 & n16852) | (n16728 & n16853) | (n16852 & n16853);
  assign n16855 = n9057 | n13981;
  assign n16856 = n9057 | n16822;
  assign n16857 = (n16728 & n16855) | (n16728 & n16856) | (n16855 & n16856);
  assign n9060 = ~n16854 & n16857;
  assign n9061 = x73 & x91;
  assign n9062 = n9060 & n9061;
  assign n9063 = n9060 | n9061;
  assign n9064 = ~n9062 & n9063;
  assign n13978 = n8845 | n8847;
  assign n14012 = n9064 & n13978;
  assign n14013 = n8845 & n9064;
  assign n14014 = (n16768 & n14012) | (n16768 & n14013) | (n14012 & n14013);
  assign n14015 = n9064 | n13978;
  assign n14016 = n8845 | n9064;
  assign n14017 = (n16768 & n14015) | (n16768 & n14016) | (n14015 & n14016);
  assign n9067 = ~n14014 & n14017;
  assign n9068 = x72 & x92;
  assign n9069 = n9067 & n9068;
  assign n9070 = n9067 | n9068;
  assign n9071 = ~n9069 & n9070;
  assign n14018 = n8852 & n9071;
  assign n16858 = (n9071 & n13918) | (n9071 & n14018) | (n13918 & n14018);
  assign n16859 = (n9071 & n13917) | (n9071 & n14018) | (n13917 & n14018);
  assign n16860 = (n13761 & n16858) | (n13761 & n16859) | (n16858 & n16859);
  assign n14020 = n8852 | n9071;
  assign n16861 = n13918 | n14020;
  assign n16862 = n13917 | n14020;
  assign n16863 = (n13761 & n16861) | (n13761 & n16862) | (n16861 & n16862);
  assign n9074 = ~n16860 & n16863;
  assign n9075 = x71 & x93;
  assign n9076 = n9074 & n9075;
  assign n9077 = n9074 | n9075;
  assign n9078 = ~n9076 & n9077;
  assign n13976 = n8859 | n8861;
  assign n16864 = n9078 & n13976;
  assign n16819 = n8634 | n8859;
  assign n16820 = (n8859 & n8861) | (n8859 & n16819) | (n8861 & n16819);
  assign n16865 = n9078 & n16820;
  assign n16866 = (n16746 & n16864) | (n16746 & n16865) | (n16864 & n16865);
  assign n16867 = n9078 | n13976;
  assign n16868 = n9078 | n16820;
  assign n16869 = (n16746 & n16867) | (n16746 & n16868) | (n16867 & n16868);
  assign n9081 = ~n16866 & n16869;
  assign n9082 = x70 & x94;
  assign n9083 = n9081 & n9082;
  assign n9084 = n9081 | n9082;
  assign n9085 = ~n9083 & n9084;
  assign n14022 = n8866 & n9085;
  assign n16870 = (n9085 & n13927) | (n9085 & n14022) | (n13927 & n14022);
  assign n16871 = (n8868 & n9085) | (n8868 & n14022) | (n9085 & n14022);
  assign n16872 = (n13827 & n16870) | (n13827 & n16871) | (n16870 & n16871);
  assign n14024 = n8866 | n9085;
  assign n16873 = n13927 | n14024;
  assign n16874 = n8868 | n14024;
  assign n16875 = (n13827 & n16873) | (n13827 & n16874) | (n16873 & n16874);
  assign n9088 = ~n16872 & n16875;
  assign n9089 = x69 & x95;
  assign n9090 = n9088 & n9089;
  assign n9091 = n9088 | n9089;
  assign n9092 = ~n9090 & n9091;
  assign n14026 = n8873 & n9092;
  assign n14027 = (n9092 & n13932) | (n9092 & n14026) | (n13932 & n14026);
  assign n14028 = n8873 | n9092;
  assign n14029 = n13932 | n14028;
  assign n9095 = ~n14027 & n14029;
  assign n9096 = x68 & x96;
  assign n9097 = n9095 & n9096;
  assign n9098 = n9095 | n9096;
  assign n9099 = ~n9097 & n9098;
  assign n14030 = n8880 & n9099;
  assign n14031 = (n9099 & n13936) | (n9099 & n14030) | (n13936 & n14030);
  assign n14032 = n8880 | n9099;
  assign n14033 = n13936 | n14032;
  assign n9102 = ~n14031 & n14033;
  assign n9103 = x67 & x97;
  assign n9104 = n9102 & n9103;
  assign n9105 = n9102 | n9103;
  assign n9106 = ~n9104 & n9105;
  assign n14034 = n8887 & n9106;
  assign n14035 = (n9106 & n13940) | (n9106 & n14034) | (n13940 & n14034);
  assign n14036 = n8887 | n9106;
  assign n14037 = n13940 | n14036;
  assign n9109 = ~n14035 & n14037;
  assign n9110 = x66 & x98;
  assign n9111 = n9109 & n9110;
  assign n9112 = n9109 | n9110;
  assign n9113 = ~n9111 & n9112;
  assign n14038 = n8894 & n9113;
  assign n14039 = (n9113 & n13945) | (n9113 & n14038) | (n13945 & n14038);
  assign n14040 = n8894 | n9113;
  assign n14041 = n13945 | n14040;
  assign n9116 = ~n14039 & n14041;
  assign n9117 = x65 & x99;
  assign n9118 = n9116 & n9117;
  assign n9119 = n9116 | n9117;
  assign n9120 = ~n9118 & n9119;
  assign n13973 = n8901 | n8903;
  assign n14042 = n9120 & n13973;
  assign n14043 = n8901 & n9120;
  assign n14044 = (n13867 & n14042) | (n13867 & n14043) | (n14042 & n14043);
  assign n14045 = n9120 | n13973;
  assign n14046 = n8901 | n9120;
  assign n14047 = (n13867 & n14045) | (n13867 & n14046) | (n14045 & n14046);
  assign n9123 = ~n14044 & n14047;
  assign n9124 = x64 & x100;
  assign n9125 = n9123 & n9124;
  assign n9126 = n9123 | n9124;
  assign n9127 = ~n9125 & n9126;
  assign n13971 = n8908 | n8910;
  assign n16876 = n9127 & n13971;
  assign n16877 = n8908 & n9127;
  assign n16878 = (n13865 & n16876) | (n13865 & n16877) | (n16876 & n16877);
  assign n16879 = n9127 | n13971;
  assign n16880 = n8908 | n9127;
  assign n16881 = (n13865 & n16879) | (n13865 & n16880) | (n16879 & n16880);
  assign n9130 = ~n16878 & n16881;
  assign n9131 = x63 & x101;
  assign n9132 = n9130 & n9131;
  assign n9133 = n9130 | n9131;
  assign n9134 = ~n9132 & n9133;
  assign n13969 = n8915 | n8917;
  assign n16882 = n9134 & n13969;
  assign n16883 = n8915 & n9134;
  assign n16884 = (n13863 & n16882) | (n13863 & n16883) | (n16882 & n16883);
  assign n16885 = n9134 | n13969;
  assign n16886 = n8915 | n9134;
  assign n16887 = (n13863 & n16885) | (n13863 & n16886) | (n16885 & n16886);
  assign n9137 = ~n16884 & n16887;
  assign n9138 = x62 & x102;
  assign n9139 = n9137 & n9138;
  assign n9140 = n9137 | n9138;
  assign n9141 = ~n9139 & n9140;
  assign n9142 = n13968 & n9141;
  assign n9143 = n13968 | n9141;
  assign n9144 = ~n9142 & n9143;
  assign n9145 = x61 & x103;
  assign n9146 = n9144 & n9145;
  assign n9147 = n9144 | n9145;
  assign n9148 = ~n9146 & n9147;
  assign n9149 = n13966 & n9148;
  assign n9150 = n13966 | n9148;
  assign n9151 = ~n9149 & n9150;
  assign n9152 = x60 & x104;
  assign n9153 = n9151 & n9152;
  assign n9154 = n9151 | n9152;
  assign n9155 = ~n9153 & n9154;
  assign n9156 = n13964 & n9155;
  assign n9157 = n13964 | n9155;
  assign n9158 = ~n9156 & n9157;
  assign n9159 = x59 & x105;
  assign n9160 = n9158 & n9159;
  assign n9161 = n9158 | n9159;
  assign n9162 = ~n9160 & n9161;
  assign n9163 = n13962 & n9162;
  assign n9164 = n13962 | n9162;
  assign n9165 = ~n9163 & n9164;
  assign n9166 = x58 & x106;
  assign n9167 = n9165 & n9166;
  assign n9168 = n9165 | n9166;
  assign n9169 = ~n9167 & n9168;
  assign n9170 = n13960 & n9169;
  assign n9171 = n13960 | n9169;
  assign n9172 = ~n9170 & n9171;
  assign n9173 = x57 & x107;
  assign n9174 = n9172 & n9173;
  assign n9175 = n9172 | n9173;
  assign n9176 = ~n9174 & n9175;
  assign n9177 = n13958 & n9176;
  assign n9178 = n13958 | n9176;
  assign n9179 = ~n9177 & n9178;
  assign n9180 = x56 & x108;
  assign n9181 = n9179 & n9180;
  assign n9182 = n9179 | n9180;
  assign n9183 = ~n9181 & n9182;
  assign n9184 = n13956 & n9183;
  assign n9185 = n13956 | n9183;
  assign n9186 = ~n9184 & n9185;
  assign n9187 = x55 & x109;
  assign n9188 = n9186 & n9187;
  assign n9189 = n9186 | n9187;
  assign n9190 = ~n9188 & n9189;
  assign n9191 = n13954 & n9190;
  assign n9192 = n13954 | n9190;
  assign n9193 = ~n9191 & n9192;
  assign n9194 = x54 & x110;
  assign n9195 = n9193 & n9194;
  assign n9196 = n9193 | n9194;
  assign n9197 = ~n9195 & n9196;
  assign n9198 = n13952 & n9197;
  assign n9199 = n13952 | n9197;
  assign n9200 = ~n9198 & n9199;
  assign n9201 = x53 & x111;
  assign n9202 = n9200 & n9201;
  assign n9203 = n9200 | n9201;
  assign n9204 = ~n9202 & n9203;
  assign n9205 = n13950 & n9204;
  assign n9206 = n13950 | n9204;
  assign n9207 = ~n9205 & n9206;
  assign n9208 = n9202 | n9205;
  assign n9209 = n9195 | n9198;
  assign n9210 = n9188 | n9191;
  assign n9211 = n9181 | n9184;
  assign n14048 = n9174 | n9176;
  assign n14049 = (n9174 & n13958) | (n9174 & n14048) | (n13958 & n14048);
  assign n14050 = n9167 | n9169;
  assign n14051 = (n9167 & n13960) | (n9167 & n14050) | (n13960 & n14050);
  assign n14052 = n9160 | n9162;
  assign n14053 = (n9160 & n13962) | (n9160 & n14052) | (n13962 & n14052);
  assign n14054 = n9153 | n9155;
  assign n14055 = (n9153 & n13964) | (n9153 & n14054) | (n13964 & n14054);
  assign n14056 = n9146 | n9148;
  assign n14057 = (n9146 & n13966) | (n9146 & n14056) | (n13966 & n14056);
  assign n13970 = (n8915 & n13863) | (n8915 & n13969) | (n13863 & n13969);
  assign n13972 = (n8908 & n13865) | (n8908 & n13971) | (n13865 & n13971);
  assign n13977 = (n16746 & n16820) | (n16746 & n13976) | (n16820 & n13976);
  assign n14067 = n9069 | n9071;
  assign n16888 = n8852 | n9069;
  assign n16889 = (n9069 & n9071) | (n9069 & n16888) | (n9071 & n16888);
  assign n16890 = (n13918 & n14067) | (n13918 & n16889) | (n14067 & n16889);
  assign n16891 = (n13917 & n14067) | (n13917 & n16889) | (n14067 & n16889);
  assign n16892 = (n13761 & n16890) | (n13761 & n16891) | (n16890 & n16891);
  assign n13982 = (n16728 & n16822) | (n16728 & n13981) | (n16822 & n13981);
  assign n16895 = n8810 | n9027;
  assign n16896 = (n9027 & n9029) | (n9027 & n16895) | (n9029 & n16895);
  assign n16897 = n9027 | n9029;
  assign n16898 = (n9027 & n13988) | (n9027 & n16897) | (n13988 & n16897);
  assign n16899 = (n13881 & n16896) | (n13881 & n16898) | (n16896 & n16898);
  assign n16900 = (n16772 & n16896) | (n16772 & n16898) | (n16896 & n16898);
  assign n16901 = (n13659 & n16899) | (n13659 & n16900) | (n16899 & n16900);
  assign n9235 = x79 & x86;
  assign n17815 = n9019 & n9235;
  assign n18066 = n17789 & n17815;
  assign n18235 = n17815 & n18049;
  assign n18205 = n16709 & n18235;
  assign n34719 = n17815 & n18243;
  assign n29526 = n16554 & n34719;
  assign n18266 = n9235 & n18261;
  assign n18267 = (n13366 & n29526) | (n13366 & n18266) | (n29526 & n18266);
  assign n18268 = (n16398 & n29526) | (n16398 & n18266) | (n29526 & n18266);
  assign n18255 = (n16133 & n18267) | (n16133 & n18268) | (n18267 & n18268);
  assign n18234 = (n8326 & n18235) | (n8326 & n18255) | (n18235 & n18255);
  assign n18203 = (n16571 & n18205) | (n16571 & n18234) | (n18205 & n18234);
  assign n18153 = n9235 & n18140;
  assign n18154 = (n8566 & n18203) | (n8566 & n18153) | (n18203 & n18153);
  assign n18152 = (n16717 & n18154) | (n16717 & n18203) | (n18154 & n18203);
  assign n18065 = (n16552 & n18066) | (n16552 & n18152) | (n18066 & n18152);
  assign n18063 = (n8798 & n17815) | (n8798 & n18065) | (n17815 & n18065);
  assign n17957 = (n16784 & n18063) | (n16784 & n18065) | (n18063 & n18065);
  assign n17958 = (n16786 & n17815) | (n16786 & n18065) | (n17815 & n18065);
  assign n17811 = (n16646 & n17957) | (n16646 & n17958) | (n17957 & n17958);
  assign n16903 = (n9022 & n9235) | (n9022 & n17811) | (n9235 & n17811);
  assign n18157 = (n16571 & n18205) | (n16571 & n18234) | (n18205 & n18234);
  assign n18069 = (n16717 & n18154) | (n16717 & n18157) | (n18154 & n18157);
  assign n17961 = (n16552 & n18066) | (n16552 & n18069) | (n18066 & n18069);
  assign n17814 = (n16784 & n18063) | (n16784 & n17961) | (n18063 & n17961);
  assign n17816 = (n16786 & n17961) | (n16786 & n17815) | (n17961 & n17815);
  assign n16906 = (n16646 & n17814) | (n16646 & n17816) | (n17814 & n17816);
  assign n16907 = (n16829 & n16903) | (n16829 & n16906) | (n16903 & n16906);
  assign n16908 = (n16831 & n16903) | (n16831 & n16906) | (n16903 & n16906);
  assign n16909 = (n16707 & n16907) | (n16707 & n16908) | (n16907 & n16908);
  assign n17823 = n9019 | n9235;
  assign n18073 = (n9235 & n17789) | (n9235 & n17823) | (n17789 & n17823);
  assign n18238 = (n9235 & n17823) | (n9235 & n18049) | (n17823 & n18049);
  assign n18210 = (n9235 & n16709) | (n9235 & n18238) | (n16709 & n18238);
  assign n34720 = (n9235 & n17823) | (n9235 & n18243) | (n17823 & n18243);
  assign n29528 = (n9235 & n16554) | (n9235 & n34720) | (n16554 & n34720);
  assign n18270 = n9235 | n18261;
  assign n18271 = (n13366 & n29528) | (n13366 & n18270) | (n29528 & n18270);
  assign n18272 = (n16398 & n29528) | (n16398 & n18270) | (n29528 & n18270);
  assign n18258 = (n16133 & n18271) | (n16133 & n18272) | (n18271 & n18272);
  assign n18237 = (n8326 & n18238) | (n8326 & n18258) | (n18238 & n18258);
  assign n18208 = (n16571 & n18210) | (n16571 & n18237) | (n18210 & n18237);
  assign n18161 = n9235 | n18140;
  assign n18162 = (n8566 & n18208) | (n8566 & n18161) | (n18208 & n18161);
  assign n18160 = (n16717 & n18162) | (n16717 & n18208) | (n18162 & n18208);
  assign n18072 = (n16552 & n18073) | (n16552 & n18160) | (n18073 & n18160);
  assign n18070 = (n8798 & n17823) | (n8798 & n18072) | (n17823 & n18072);
  assign n17964 = (n16784 & n18070) | (n16784 & n18072) | (n18070 & n18072);
  assign n17965 = (n16786 & n17823) | (n16786 & n18072) | (n17823 & n18072);
  assign n17819 = (n16646 & n17964) | (n16646 & n17965) | (n17964 & n17965);
  assign n16911 = n9022 | n17819;
  assign n18165 = (n16571 & n18210) | (n16571 & n18237) | (n18210 & n18237);
  assign n18076 = (n16717 & n18162) | (n16717 & n18165) | (n18162 & n18165);
  assign n17968 = (n16552 & n18073) | (n16552 & n18076) | (n18073 & n18076);
  assign n17822 = (n16784 & n18070) | (n16784 & n17968) | (n18070 & n17968);
  assign n17824 = (n16786 & n17968) | (n16786 & n17823) | (n17968 & n17823);
  assign n16914 = (n16646 & n17822) | (n16646 & n17824) | (n17822 & n17824);
  assign n16915 = (n16829 & n16911) | (n16829 & n16914) | (n16911 & n16914);
  assign n16916 = (n16831 & n16911) | (n16831 & n16914) | (n16911 & n16914);
  assign n16917 = (n16707 & n16915) | (n16707 & n16916) | (n16915 & n16916);
  assign n9238 = ~n16909 & n16917;
  assign n9239 = n16901 & n9238;
  assign n9240 = n16901 | n9238;
  assign n9241 = ~n9239 & n9240;
  assign n9242 = x78 & x87;
  assign n9243 = n9241 & n9242;
  assign n9244 = n9241 | n9242;
  assign n9245 = ~n9243 & n9244;
  assign n14074 = n9034 | n9036;
  assign n14087 = n9245 & n14074;
  assign n14088 = n9034 & n9245;
  assign n14089 = (n16827 & n14087) | (n16827 & n14088) | (n14087 & n14088);
  assign n14090 = n9245 | n14074;
  assign n14091 = n9034 | n9245;
  assign n14092 = (n16827 & n14090) | (n16827 & n14091) | (n14090 & n14091);
  assign n9248 = ~n14089 & n14092;
  assign n9249 = x77 & x88;
  assign n9250 = n9248 & n9249;
  assign n9251 = n9248 | n9249;
  assign n9252 = ~n9250 & n9251;
  assign n14093 = n9041 & n9252;
  assign n16918 = (n9252 & n14003) | (n9252 & n14093) | (n14003 & n14093);
  assign n16919 = (n9252 & n14002) | (n9252 & n14093) | (n14002 & n14093);
  assign n16920 = (n13879 & n16918) | (n13879 & n16919) | (n16918 & n16919);
  assign n14095 = n9041 | n9252;
  assign n16921 = n14003 | n14095;
  assign n16922 = n14002 | n14095;
  assign n16923 = (n13879 & n16921) | (n13879 & n16922) | (n16921 & n16922);
  assign n9255 = ~n16920 & n16923;
  assign n9256 = x76 & x89;
  assign n9257 = n9255 & n9256;
  assign n9258 = n9255 | n9256;
  assign n9259 = ~n9257 & n9258;
  assign n14072 = n9048 | n9050;
  assign n16924 = n9259 & n14072;
  assign n16893 = n8831 | n9048;
  assign n16894 = (n9048 & n9050) | (n9048 & n16893) | (n9050 & n16893);
  assign n16925 = n9259 & n16894;
  assign n16926 = (n13909 & n16924) | (n13909 & n16925) | (n16924 & n16925);
  assign n16927 = n9259 | n14072;
  assign n16928 = n9259 | n16894;
  assign n16929 = (n13909 & n16927) | (n13909 & n16928) | (n16927 & n16928);
  assign n9262 = ~n16926 & n16929;
  assign n9263 = x75 & x90;
  assign n9264 = n9262 & n9263;
  assign n9265 = n9262 | n9263;
  assign n9266 = ~n9264 & n9265;
  assign n14069 = n9055 | n9057;
  assign n14097 = n9266 & n14069;
  assign n14098 = n9055 & n9266;
  assign n14099 = (n13982 & n14097) | (n13982 & n14098) | (n14097 & n14098);
  assign n14100 = n9266 | n14069;
  assign n14101 = n9055 | n9266;
  assign n14102 = (n13982 & n14100) | (n13982 & n14101) | (n14100 & n14101);
  assign n9269 = ~n14099 & n14102;
  assign n9270 = x74 & x91;
  assign n9271 = n9269 & n9270;
  assign n9272 = n9269 | n9270;
  assign n9273 = ~n9271 & n9272;
  assign n14103 = n9062 & n9273;
  assign n16930 = (n9273 & n14012) | (n9273 & n14103) | (n14012 & n14103);
  assign n16931 = (n9273 & n14013) | (n9273 & n14103) | (n14013 & n14103);
  assign n16932 = (n16768 & n16930) | (n16768 & n16931) | (n16930 & n16931);
  assign n14105 = n9062 | n9273;
  assign n16933 = n14012 | n14105;
  assign n16934 = n14013 | n14105;
  assign n16935 = (n16768 & n16933) | (n16768 & n16934) | (n16933 & n16934);
  assign n9276 = ~n16932 & n16935;
  assign n9277 = x73 & x92;
  assign n9278 = n9276 & n9277;
  assign n9279 = n9276 | n9277;
  assign n9280 = ~n9278 & n9279;
  assign n9281 = n16892 & n9280;
  assign n9282 = n16892 | n9280;
  assign n9283 = ~n9281 & n9282;
  assign n9284 = x72 & x93;
  assign n9285 = n9283 & n9284;
  assign n9286 = n9283 | n9284;
  assign n9287 = ~n9285 & n9286;
  assign n14064 = n9076 | n9078;
  assign n14107 = n9287 & n14064;
  assign n14108 = n9076 & n9287;
  assign n14109 = (n13977 & n14107) | (n13977 & n14108) | (n14107 & n14108);
  assign n14110 = n9287 | n14064;
  assign n14111 = n9076 | n9287;
  assign n14112 = (n13977 & n14110) | (n13977 & n14111) | (n14110 & n14111);
  assign n9290 = ~n14109 & n14112;
  assign n9291 = x71 & x94;
  assign n9292 = n9290 & n9291;
  assign n9293 = n9290 | n9291;
  assign n9294 = ~n9292 & n9293;
  assign n14113 = n9083 & n9294;
  assign n14114 = (n9294 & n16872) | (n9294 & n14113) | (n16872 & n14113);
  assign n14115 = n9083 | n9294;
  assign n14116 = n16872 | n14115;
  assign n9297 = ~n14114 & n14116;
  assign n9298 = x70 & x95;
  assign n9299 = n9297 & n9298;
  assign n9300 = n9297 | n9298;
  assign n9301 = ~n9299 & n9300;
  assign n14117 = n9090 & n9301;
  assign n14118 = (n9301 & n14027) | (n9301 & n14117) | (n14027 & n14117);
  assign n14119 = n9090 | n9301;
  assign n14120 = n14027 | n14119;
  assign n9304 = ~n14118 & n14120;
  assign n9305 = x69 & x96;
  assign n9306 = n9304 & n9305;
  assign n9307 = n9304 | n9305;
  assign n9308 = ~n9306 & n9307;
  assign n14121 = n9097 & n9308;
  assign n14122 = (n9308 & n14031) | (n9308 & n14121) | (n14031 & n14121);
  assign n14123 = n9097 | n9308;
  assign n14124 = n14031 | n14123;
  assign n9311 = ~n14122 & n14124;
  assign n9312 = x68 & x97;
  assign n9313 = n9311 & n9312;
  assign n9314 = n9311 | n9312;
  assign n9315 = ~n9313 & n9314;
  assign n14125 = n9104 & n9315;
  assign n14126 = (n9315 & n14035) | (n9315 & n14125) | (n14035 & n14125);
  assign n14127 = n9104 | n9315;
  assign n14128 = n14035 | n14127;
  assign n9318 = ~n14126 & n14128;
  assign n9319 = x67 & x98;
  assign n9320 = n9318 & n9319;
  assign n9321 = n9318 | n9319;
  assign n9322 = ~n9320 & n9321;
  assign n14129 = n9111 & n9322;
  assign n14130 = (n9322 & n14039) | (n9322 & n14129) | (n14039 & n14129);
  assign n14131 = n9111 | n9322;
  assign n14132 = n14039 | n14131;
  assign n9325 = ~n14130 & n14132;
  assign n9326 = x66 & x99;
  assign n9327 = n9325 & n9326;
  assign n9328 = n9325 | n9326;
  assign n9329 = ~n9327 & n9328;
  assign n14133 = n9118 & n9329;
  assign n14134 = (n9329 & n14044) | (n9329 & n14133) | (n14044 & n14133);
  assign n14135 = n9118 | n9329;
  assign n14136 = n14044 | n14135;
  assign n9332 = ~n14134 & n14136;
  assign n9333 = x65 & x100;
  assign n9334 = n9332 & n9333;
  assign n9335 = n9332 | n9333;
  assign n9336 = ~n9334 & n9335;
  assign n14062 = n9125 | n9127;
  assign n14137 = n9336 & n14062;
  assign n14138 = n9125 & n9336;
  assign n14139 = (n13972 & n14137) | (n13972 & n14138) | (n14137 & n14138);
  assign n14140 = n9336 | n14062;
  assign n14141 = n9125 | n9336;
  assign n14142 = (n13972 & n14140) | (n13972 & n14141) | (n14140 & n14141);
  assign n9339 = ~n14139 & n14142;
  assign n9340 = x64 & x101;
  assign n9341 = n9339 & n9340;
  assign n9342 = n9339 | n9340;
  assign n9343 = ~n9341 & n9342;
  assign n14060 = n9132 | n9134;
  assign n16936 = n9343 & n14060;
  assign n16937 = n9132 & n9343;
  assign n16938 = (n13970 & n16936) | (n13970 & n16937) | (n16936 & n16937);
  assign n16939 = n9343 | n14060;
  assign n16940 = n9132 | n9343;
  assign n16941 = (n13970 & n16939) | (n13970 & n16940) | (n16939 & n16940);
  assign n9346 = ~n16938 & n16941;
  assign n9347 = x63 & x102;
  assign n9348 = n9346 & n9347;
  assign n9349 = n9346 | n9347;
  assign n9350 = ~n9348 & n9349;
  assign n14058 = n9139 | n9141;
  assign n16942 = n9350 & n14058;
  assign n16943 = n9139 & n9350;
  assign n16944 = (n13968 & n16942) | (n13968 & n16943) | (n16942 & n16943);
  assign n16945 = n9350 | n14058;
  assign n16946 = n9139 | n9350;
  assign n16947 = (n13968 & n16945) | (n13968 & n16946) | (n16945 & n16946);
  assign n9353 = ~n16944 & n16947;
  assign n9354 = x62 & x103;
  assign n9355 = n9353 & n9354;
  assign n9356 = n9353 | n9354;
  assign n9357 = ~n9355 & n9356;
  assign n9358 = n14057 & n9357;
  assign n9359 = n14057 | n9357;
  assign n9360 = ~n9358 & n9359;
  assign n9361 = x61 & x104;
  assign n9362 = n9360 & n9361;
  assign n9363 = n9360 | n9361;
  assign n9364 = ~n9362 & n9363;
  assign n9365 = n14055 & n9364;
  assign n9366 = n14055 | n9364;
  assign n9367 = ~n9365 & n9366;
  assign n9368 = x60 & x105;
  assign n9369 = n9367 & n9368;
  assign n9370 = n9367 | n9368;
  assign n9371 = ~n9369 & n9370;
  assign n9372 = n14053 & n9371;
  assign n9373 = n14053 | n9371;
  assign n9374 = ~n9372 & n9373;
  assign n9375 = x59 & x106;
  assign n9376 = n9374 & n9375;
  assign n9377 = n9374 | n9375;
  assign n9378 = ~n9376 & n9377;
  assign n9379 = n14051 & n9378;
  assign n9380 = n14051 | n9378;
  assign n9381 = ~n9379 & n9380;
  assign n9382 = x58 & x107;
  assign n9383 = n9381 & n9382;
  assign n9384 = n9381 | n9382;
  assign n9385 = ~n9383 & n9384;
  assign n9386 = n14049 & n9385;
  assign n9387 = n14049 | n9385;
  assign n9388 = ~n9386 & n9387;
  assign n9389 = x57 & x108;
  assign n9390 = n9388 & n9389;
  assign n9391 = n9388 | n9389;
  assign n9392 = ~n9390 & n9391;
  assign n9393 = n9211 & n9392;
  assign n9394 = n9211 | n9392;
  assign n9395 = ~n9393 & n9394;
  assign n9396 = x56 & x109;
  assign n9397 = n9395 & n9396;
  assign n9398 = n9395 | n9396;
  assign n9399 = ~n9397 & n9398;
  assign n9400 = n9210 & n9399;
  assign n9401 = n9210 | n9399;
  assign n9402 = ~n9400 & n9401;
  assign n9403 = x55 & x110;
  assign n9404 = n9402 & n9403;
  assign n9405 = n9402 | n9403;
  assign n9406 = ~n9404 & n9405;
  assign n9407 = n9209 & n9406;
  assign n9408 = n9209 | n9406;
  assign n9409 = ~n9407 & n9408;
  assign n9410 = x54 & x111;
  assign n9411 = n9409 & n9410;
  assign n9412 = n9409 | n9410;
  assign n9413 = ~n9411 & n9412;
  assign n9414 = n9208 & n9413;
  assign n9415 = n9208 | n9413;
  assign n9416 = ~n9414 & n9415;
  assign n9417 = n9411 | n9414;
  assign n9418 = n9404 | n9407;
  assign n9419 = n9397 | n9400;
  assign n14143 = n9390 | n9392;
  assign n14144 = (n9211 & n9390) | (n9211 & n14143) | (n9390 & n14143);
  assign n14145 = n9383 | n9385;
  assign n14146 = (n9383 & n14049) | (n9383 & n14145) | (n14049 & n14145);
  assign n14147 = n9376 | n9378;
  assign n14148 = (n9376 & n14051) | (n9376 & n14147) | (n14051 & n14147);
  assign n14149 = n9369 | n9371;
  assign n14150 = (n9369 & n14053) | (n9369 & n14149) | (n14053 & n14149);
  assign n14151 = n9362 | n9364;
  assign n14152 = (n9362 & n14055) | (n9362 & n14151) | (n14055 & n14151);
  assign n14059 = (n9139 & n13968) | (n9139 & n14058) | (n13968 & n14058);
  assign n14061 = (n9132 & n13970) | (n9132 & n14060) | (n13970 & n14060);
  assign n14165 = n9271 | n9273;
  assign n16950 = n9062 | n9271;
  assign n16951 = (n9271 & n9273) | (n9271 & n16950) | (n9273 & n16950);
  assign n16952 = (n14012 & n14165) | (n14012 & n16951) | (n14165 & n16951);
  assign n16953 = (n14013 & n14165) | (n14013 & n16951) | (n14165 & n16951);
  assign n16954 = (n16768 & n16952) | (n16768 & n16953) | (n16952 & n16953);
  assign n14073 = (n13909 & n16894) | (n13909 & n14072) | (n16894 & n14072);
  assign n14170 = n9250 | n9252;
  assign n16955 = n9041 | n9250;
  assign n16956 = (n9250 & n9252) | (n9250 & n16955) | (n9252 & n16955);
  assign n16957 = (n14003 & n14170) | (n14003 & n16956) | (n14170 & n16956);
  assign n16958 = (n14002 & n14170) | (n14002 & n16956) | (n14170 & n16956);
  assign n16959 = (n13879 & n16957) | (n13879 & n16958) | (n16957 & n16958);
  assign n16960 = n9034 | n9243;
  assign n16961 = (n9243 & n9245) | (n9243 & n16960) | (n9245 & n16960);
  assign n14173 = n9243 | n14087;
  assign n14174 = (n16827 & n16961) | (n16827 & n14173) | (n16961 & n14173);
  assign n9443 = x79 & x87;
  assign n16962 = n9443 & n16909;
  assign n16963 = (n9238 & n9443) | (n9238 & n16962) | (n9443 & n16962);
  assign n14178 = n9443 & n16909;
  assign n14179 = (n16901 & n16963) | (n16901 & n14178) | (n16963 & n14178);
  assign n16964 = n9443 | n16909;
  assign n16965 = n9238 | n16964;
  assign n14181 = n9443 | n16909;
  assign n14182 = (n16901 & n16965) | (n16901 & n14181) | (n16965 & n14181);
  assign n9446 = ~n14179 & n14182;
  assign n9447 = n14174 & n9446;
  assign n9448 = n14174 | n9446;
  assign n9449 = ~n9447 & n9448;
  assign n9450 = x78 & x88;
  assign n9451 = n9449 & n9450;
  assign n9452 = n9449 | n9450;
  assign n9453 = ~n9451 & n9452;
  assign n9454 = n16959 & n9453;
  assign n9455 = n16959 | n9453;
  assign n9456 = ~n9454 & n9455;
  assign n9457 = x77 & x89;
  assign n9458 = n9456 & n9457;
  assign n9459 = n9456 | n9457;
  assign n9460 = ~n9458 & n9459;
  assign n14167 = n9257 | n9259;
  assign n14183 = n9460 & n14167;
  assign n14184 = n9257 & n9460;
  assign n14185 = (n14073 & n14183) | (n14073 & n14184) | (n14183 & n14184);
  assign n14186 = n9460 | n14167;
  assign n14187 = n9257 | n9460;
  assign n14188 = (n14073 & n14186) | (n14073 & n14187) | (n14186 & n14187);
  assign n9463 = ~n14185 & n14188;
  assign n9464 = x76 & x90;
  assign n9465 = n9463 & n9464;
  assign n9466 = n9463 | n9464;
  assign n9467 = ~n9465 & n9466;
  assign n14189 = n9264 & n9467;
  assign n16966 = (n9467 & n14097) | (n9467 & n14189) | (n14097 & n14189);
  assign n16967 = (n9467 & n14098) | (n9467 & n14189) | (n14098 & n14189);
  assign n16968 = (n13982 & n16966) | (n13982 & n16967) | (n16966 & n16967);
  assign n14191 = n9264 | n9467;
  assign n16969 = n14097 | n14191;
  assign n16970 = n14098 | n14191;
  assign n16971 = (n13982 & n16969) | (n13982 & n16970) | (n16969 & n16970);
  assign n9470 = ~n16968 & n16971;
  assign n9471 = x75 & x91;
  assign n9472 = n9470 & n9471;
  assign n9473 = n9470 | n9471;
  assign n9474 = ~n9472 & n9473;
  assign n9475 = n16954 & n9474;
  assign n9476 = n16954 | n9474;
  assign n9477 = ~n9475 & n9476;
  assign n9478 = x74 & x92;
  assign n9479 = n9477 & n9478;
  assign n9480 = n9477 | n9478;
  assign n9481 = ~n9479 & n9480;
  assign n14162 = n9278 | n9280;
  assign n14193 = n9481 & n14162;
  assign n14194 = n9278 & n9481;
  assign n14195 = (n16892 & n14193) | (n16892 & n14194) | (n14193 & n14194);
  assign n14196 = n9481 | n14162;
  assign n14197 = n9278 | n9481;
  assign n14198 = (n16892 & n14196) | (n16892 & n14197) | (n14196 & n14197);
  assign n9484 = ~n14195 & n14198;
  assign n9485 = x73 & x93;
  assign n9486 = n9484 & n9485;
  assign n9487 = n9484 | n9485;
  assign n9488 = ~n9486 & n9487;
  assign n14199 = n9285 & n9488;
  assign n16972 = (n9488 & n14108) | (n9488 & n14199) | (n14108 & n14199);
  assign n16973 = (n9488 & n14107) | (n9488 & n14199) | (n14107 & n14199);
  assign n16974 = (n13977 & n16972) | (n13977 & n16973) | (n16972 & n16973);
  assign n14201 = n9285 | n9488;
  assign n16975 = n14108 | n14201;
  assign n16976 = n14107 | n14201;
  assign n16977 = (n13977 & n16975) | (n13977 & n16976) | (n16975 & n16976);
  assign n9491 = ~n16974 & n16977;
  assign n9492 = x72 & x94;
  assign n9493 = n9491 & n9492;
  assign n9494 = n9491 | n9492;
  assign n9495 = ~n9493 & n9494;
  assign n14160 = n9292 | n9294;
  assign n16978 = n9495 & n14160;
  assign n16948 = n9083 | n9292;
  assign n16949 = (n9292 & n9294) | (n9292 & n16948) | (n9294 & n16948);
  assign n16979 = n9495 & n16949;
  assign n16980 = (n16872 & n16978) | (n16872 & n16979) | (n16978 & n16979);
  assign n16981 = n9495 | n14160;
  assign n16982 = n9495 | n16949;
  assign n16983 = (n16872 & n16981) | (n16872 & n16982) | (n16981 & n16982);
  assign n9498 = ~n16980 & n16983;
  assign n9499 = x71 & x95;
  assign n9500 = n9498 & n9499;
  assign n9501 = n9498 | n9499;
  assign n9502 = ~n9500 & n9501;
  assign n14203 = n9299 & n9502;
  assign n16984 = (n9502 & n14117) | (n9502 & n14203) | (n14117 & n14203);
  assign n16985 = (n9301 & n9502) | (n9301 & n14203) | (n9502 & n14203);
  assign n16986 = (n14027 & n16984) | (n14027 & n16985) | (n16984 & n16985);
  assign n14205 = n9299 | n9502;
  assign n16987 = n14117 | n14205;
  assign n16988 = n9301 | n14205;
  assign n16989 = (n14027 & n16987) | (n14027 & n16988) | (n16987 & n16988);
  assign n9505 = ~n16986 & n16989;
  assign n9506 = x70 & x96;
  assign n9507 = n9505 & n9506;
  assign n9508 = n9505 | n9506;
  assign n9509 = ~n9507 & n9508;
  assign n14207 = n9306 & n9509;
  assign n14208 = (n9509 & n14122) | (n9509 & n14207) | (n14122 & n14207);
  assign n14209 = n9306 | n9509;
  assign n14210 = n14122 | n14209;
  assign n9512 = ~n14208 & n14210;
  assign n9513 = x69 & x97;
  assign n9514 = n9512 & n9513;
  assign n9515 = n9512 | n9513;
  assign n9516 = ~n9514 & n9515;
  assign n14211 = n9313 & n9516;
  assign n14212 = (n9516 & n14126) | (n9516 & n14211) | (n14126 & n14211);
  assign n14213 = n9313 | n9516;
  assign n14214 = n14126 | n14213;
  assign n9519 = ~n14212 & n14214;
  assign n9520 = x68 & x98;
  assign n9521 = n9519 & n9520;
  assign n9522 = n9519 | n9520;
  assign n9523 = ~n9521 & n9522;
  assign n14215 = n9320 & n9523;
  assign n14216 = (n9523 & n14130) | (n9523 & n14215) | (n14130 & n14215);
  assign n14217 = n9320 | n9523;
  assign n14218 = n14130 | n14217;
  assign n9526 = ~n14216 & n14218;
  assign n9527 = x67 & x99;
  assign n9528 = n9526 & n9527;
  assign n9529 = n9526 | n9527;
  assign n9530 = ~n9528 & n9529;
  assign n14219 = n9327 & n9530;
  assign n14220 = (n9530 & n14134) | (n9530 & n14219) | (n14134 & n14219);
  assign n14221 = n9327 | n9530;
  assign n14222 = n14134 | n14221;
  assign n9533 = ~n14220 & n14222;
  assign n9534 = x66 & x100;
  assign n9535 = n9533 & n9534;
  assign n9536 = n9533 | n9534;
  assign n9537 = ~n9535 & n9536;
  assign n14223 = n9334 & n9537;
  assign n14224 = (n9537 & n14139) | (n9537 & n14223) | (n14139 & n14223);
  assign n14225 = n9334 | n9537;
  assign n14226 = n14139 | n14225;
  assign n9540 = ~n14224 & n14226;
  assign n9541 = x65 & x101;
  assign n9542 = n9540 & n9541;
  assign n9543 = n9540 | n9541;
  assign n9544 = ~n9542 & n9543;
  assign n14157 = n9341 | n9343;
  assign n14227 = n9544 & n14157;
  assign n14228 = n9341 & n9544;
  assign n14229 = (n14061 & n14227) | (n14061 & n14228) | (n14227 & n14228);
  assign n14230 = n9544 | n14157;
  assign n14231 = n9341 | n9544;
  assign n14232 = (n14061 & n14230) | (n14061 & n14231) | (n14230 & n14231);
  assign n9547 = ~n14229 & n14232;
  assign n9548 = x64 & x102;
  assign n9549 = n9547 & n9548;
  assign n9550 = n9547 | n9548;
  assign n9551 = ~n9549 & n9550;
  assign n14155 = n9348 | n9350;
  assign n16990 = n9551 & n14155;
  assign n16991 = n9348 & n9551;
  assign n16992 = (n14059 & n16990) | (n14059 & n16991) | (n16990 & n16991);
  assign n16993 = n9551 | n14155;
  assign n16994 = n9348 | n9551;
  assign n16995 = (n14059 & n16993) | (n14059 & n16994) | (n16993 & n16994);
  assign n9554 = ~n16992 & n16995;
  assign n9555 = x63 & x103;
  assign n9556 = n9554 & n9555;
  assign n9557 = n9554 | n9555;
  assign n9558 = ~n9556 & n9557;
  assign n14153 = n9355 | n9357;
  assign n16996 = n9558 & n14153;
  assign n16997 = n9355 & n9558;
  assign n16998 = (n14057 & n16996) | (n14057 & n16997) | (n16996 & n16997);
  assign n16999 = n9558 | n14153;
  assign n17000 = n9355 | n9558;
  assign n17001 = (n14057 & n16999) | (n14057 & n17000) | (n16999 & n17000);
  assign n9561 = ~n16998 & n17001;
  assign n9562 = x62 & x104;
  assign n9563 = n9561 & n9562;
  assign n9564 = n9561 | n9562;
  assign n9565 = ~n9563 & n9564;
  assign n9566 = n14152 & n9565;
  assign n9567 = n14152 | n9565;
  assign n9568 = ~n9566 & n9567;
  assign n9569 = x61 & x105;
  assign n9570 = n9568 & n9569;
  assign n9571 = n9568 | n9569;
  assign n9572 = ~n9570 & n9571;
  assign n9573 = n14150 & n9572;
  assign n9574 = n14150 | n9572;
  assign n9575 = ~n9573 & n9574;
  assign n9576 = x60 & x106;
  assign n9577 = n9575 & n9576;
  assign n9578 = n9575 | n9576;
  assign n9579 = ~n9577 & n9578;
  assign n9580 = n14148 & n9579;
  assign n9581 = n14148 | n9579;
  assign n9582 = ~n9580 & n9581;
  assign n9583 = x59 & x107;
  assign n9584 = n9582 & n9583;
  assign n9585 = n9582 | n9583;
  assign n9586 = ~n9584 & n9585;
  assign n9587 = n14146 & n9586;
  assign n9588 = n14146 | n9586;
  assign n9589 = ~n9587 & n9588;
  assign n9590 = x58 & x108;
  assign n9591 = n9589 & n9590;
  assign n9592 = n9589 | n9590;
  assign n9593 = ~n9591 & n9592;
  assign n9594 = n14144 & n9593;
  assign n9595 = n14144 | n9593;
  assign n9596 = ~n9594 & n9595;
  assign n9597 = x57 & x109;
  assign n9598 = n9596 & n9597;
  assign n9599 = n9596 | n9597;
  assign n9600 = ~n9598 & n9599;
  assign n9601 = n9419 & n9600;
  assign n9602 = n9419 | n9600;
  assign n9603 = ~n9601 & n9602;
  assign n9604 = x56 & x110;
  assign n9605 = n9603 & n9604;
  assign n9606 = n9603 | n9604;
  assign n9607 = ~n9605 & n9606;
  assign n9608 = n9418 & n9607;
  assign n9609 = n9418 | n9607;
  assign n9610 = ~n9608 & n9609;
  assign n9611 = x55 & x111;
  assign n9612 = n9610 & n9611;
  assign n9613 = n9610 | n9611;
  assign n9614 = ~n9612 & n9613;
  assign n9615 = n9417 & n9614;
  assign n9616 = n9417 | n9614;
  assign n9617 = ~n9615 & n9616;
  assign n9618 = n9612 | n9615;
  assign n9619 = n9605 | n9608;
  assign n14233 = n9598 | n9600;
  assign n14234 = (n9419 & n9598) | (n9419 & n14233) | (n9598 & n14233);
  assign n14235 = n9591 | n9593;
  assign n14236 = (n9591 & n14144) | (n9591 & n14235) | (n14144 & n14235);
  assign n14237 = n9584 | n9586;
  assign n14238 = (n9584 & n14146) | (n9584 & n14237) | (n14146 & n14237);
  assign n14239 = n9577 | n9579;
  assign n14240 = (n9577 & n14148) | (n9577 & n14239) | (n14148 & n14239);
  assign n14241 = n9570 | n9572;
  assign n14242 = (n9570 & n14150) | (n9570 & n14241) | (n14150 & n14241);
  assign n14154 = (n9355 & n14057) | (n9355 & n14153) | (n14057 & n14153);
  assign n14156 = (n9348 & n14059) | (n9348 & n14155) | (n14059 & n14155);
  assign n14161 = (n16872 & n16949) | (n16872 & n14160) | (n16949 & n14160);
  assign n14252 = n9486 | n9488;
  assign n17002 = n9285 | n9486;
  assign n17003 = (n9486 & n9488) | (n9486 & n17002) | (n9488 & n17002);
  assign n17004 = (n14108 & n14252) | (n14108 & n17003) | (n14252 & n17003);
  assign n17005 = (n14107 & n14252) | (n14107 & n17003) | (n14252 & n17003);
  assign n17006 = (n13977 & n17004) | (n13977 & n17005) | (n17004 & n17005);
  assign n14257 = n9465 | n9467;
  assign n17007 = n9264 | n9465;
  assign n17008 = (n9465 & n9467) | (n9465 & n17007) | (n9467 & n17007);
  assign n17009 = (n14097 & n14257) | (n14097 & n17008) | (n14257 & n17008);
  assign n17010 = (n14098 & n14257) | (n14098 & n17008) | (n14257 & n17008);
  assign n17011 = (n13982 & n17009) | (n13982 & n17010) | (n17009 & n17010);
  assign n9643 = x79 & x88;
  assign n17013 = n9643 & n16963;
  assign n17825 = n9443 & n9643;
  assign n17826 = n16909 & n17825;
  assign n17015 = (n16901 & n17013) | (n16901 & n17826) | (n17013 & n17826);
  assign n17012 = (n9446 & n9643) | (n9446 & n17015) | (n9643 & n17015);
  assign n14265 = (n14174 & n17012) | (n14174 & n17015) | (n17012 & n17015);
  assign n17017 = n9643 | n16963;
  assign n17827 = n9443 | n9643;
  assign n17828 = (n9643 & n16909) | (n9643 & n17827) | (n16909 & n17827);
  assign n17019 = (n16901 & n17017) | (n16901 & n17828) | (n17017 & n17828);
  assign n17016 = n9446 | n17019;
  assign n14268 = (n14174 & n17016) | (n14174 & n17019) | (n17016 & n17019);
  assign n9646 = ~n14265 & n14268;
  assign n14270 = n9451 & n9646;
  assign n17020 = (n9453 & n9646) | (n9453 & n14270) | (n9646 & n14270);
  assign n14271 = (n16959 & n17020) | (n16959 & n14270) | (n17020 & n14270);
  assign n14273 = n9451 | n9646;
  assign n17021 = n9453 | n14273;
  assign n14274 = (n16959 & n17021) | (n16959 & n14273) | (n17021 & n14273);
  assign n9649 = ~n14271 & n14274;
  assign n9650 = x78 & x89;
  assign n9651 = n9649 & n9650;
  assign n9652 = n9649 | n9650;
  assign n9653 = ~n9651 & n9652;
  assign n14275 = n9458 & n9653;
  assign n17022 = (n9653 & n14184) | (n9653 & n14275) | (n14184 & n14275);
  assign n17023 = (n9653 & n14183) | (n9653 & n14275) | (n14183 & n14275);
  assign n17024 = (n14073 & n17022) | (n14073 & n17023) | (n17022 & n17023);
  assign n14277 = n9458 | n9653;
  assign n17025 = n14184 | n14277;
  assign n17026 = n14183 | n14277;
  assign n17027 = (n14073 & n17025) | (n14073 & n17026) | (n17025 & n17026);
  assign n9656 = ~n17024 & n17027;
  assign n9657 = x77 & x90;
  assign n9658 = n9656 & n9657;
  assign n9659 = n9656 | n9657;
  assign n9660 = ~n9658 & n9659;
  assign n9661 = n17011 & n9660;
  assign n9662 = n17011 | n9660;
  assign n9663 = ~n9661 & n9662;
  assign n9664 = x76 & x91;
  assign n9665 = n9663 & n9664;
  assign n9666 = n9663 | n9664;
  assign n9667 = ~n9665 & n9666;
  assign n14254 = n9472 | n9474;
  assign n14279 = n9667 & n14254;
  assign n14280 = n9472 & n9667;
  assign n14281 = (n16954 & n14279) | (n16954 & n14280) | (n14279 & n14280);
  assign n14282 = n9667 | n14254;
  assign n14283 = n9472 | n9667;
  assign n14284 = (n16954 & n14282) | (n16954 & n14283) | (n14282 & n14283);
  assign n9670 = ~n14281 & n14284;
  assign n9671 = x75 & x92;
  assign n9672 = n9670 & n9671;
  assign n9673 = n9670 | n9671;
  assign n9674 = ~n9672 & n9673;
  assign n14285 = n9479 & n9674;
  assign n17028 = (n9674 & n14194) | (n9674 & n14285) | (n14194 & n14285);
  assign n17029 = (n9674 & n14193) | (n9674 & n14285) | (n14193 & n14285);
  assign n17030 = (n16892 & n17028) | (n16892 & n17029) | (n17028 & n17029);
  assign n14287 = n9479 | n9674;
  assign n17031 = n14194 | n14287;
  assign n17032 = n14193 | n14287;
  assign n17033 = (n16892 & n17031) | (n16892 & n17032) | (n17031 & n17032);
  assign n9677 = ~n17030 & n17033;
  assign n9678 = x74 & x93;
  assign n9679 = n9677 & n9678;
  assign n9680 = n9677 | n9678;
  assign n9681 = ~n9679 & n9680;
  assign n9682 = n17006 & n9681;
  assign n9683 = n17006 | n9681;
  assign n9684 = ~n9682 & n9683;
  assign n9685 = x73 & x94;
  assign n9686 = n9684 & n9685;
  assign n9687 = n9684 | n9685;
  assign n9688 = ~n9686 & n9687;
  assign n14249 = n9493 | n9495;
  assign n14289 = n9688 & n14249;
  assign n14290 = n9493 & n9688;
  assign n14291 = (n14161 & n14289) | (n14161 & n14290) | (n14289 & n14290);
  assign n14292 = n9688 | n14249;
  assign n14293 = n9493 | n9688;
  assign n14294 = (n14161 & n14292) | (n14161 & n14293) | (n14292 & n14293);
  assign n9691 = ~n14291 & n14294;
  assign n9692 = x72 & x95;
  assign n9693 = n9691 & n9692;
  assign n9694 = n9691 | n9692;
  assign n9695 = ~n9693 & n9694;
  assign n14295 = n9500 & n9695;
  assign n14296 = (n9695 & n16986) | (n9695 & n14295) | (n16986 & n14295);
  assign n14297 = n9500 | n9695;
  assign n14298 = n16986 | n14297;
  assign n9698 = ~n14296 & n14298;
  assign n9699 = x71 & x96;
  assign n9700 = n9698 & n9699;
  assign n9701 = n9698 | n9699;
  assign n9702 = ~n9700 & n9701;
  assign n14299 = n9507 & n9702;
  assign n14300 = (n9702 & n14208) | (n9702 & n14299) | (n14208 & n14299);
  assign n14301 = n9507 | n9702;
  assign n14302 = n14208 | n14301;
  assign n9705 = ~n14300 & n14302;
  assign n9706 = x70 & x97;
  assign n9707 = n9705 & n9706;
  assign n9708 = n9705 | n9706;
  assign n9709 = ~n9707 & n9708;
  assign n14303 = n9514 & n9709;
  assign n14304 = (n9709 & n14212) | (n9709 & n14303) | (n14212 & n14303);
  assign n14305 = n9514 | n9709;
  assign n14306 = n14212 | n14305;
  assign n9712 = ~n14304 & n14306;
  assign n9713 = x69 & x98;
  assign n9714 = n9712 & n9713;
  assign n9715 = n9712 | n9713;
  assign n9716 = ~n9714 & n9715;
  assign n14307 = n9521 & n9716;
  assign n14308 = (n9716 & n14216) | (n9716 & n14307) | (n14216 & n14307);
  assign n14309 = n9521 | n9716;
  assign n14310 = n14216 | n14309;
  assign n9719 = ~n14308 & n14310;
  assign n9720 = x68 & x99;
  assign n9721 = n9719 & n9720;
  assign n9722 = n9719 | n9720;
  assign n9723 = ~n9721 & n9722;
  assign n14311 = n9528 & n9723;
  assign n14312 = (n9723 & n14220) | (n9723 & n14311) | (n14220 & n14311);
  assign n14313 = n9528 | n9723;
  assign n14314 = n14220 | n14313;
  assign n9726 = ~n14312 & n14314;
  assign n9727 = x67 & x100;
  assign n9728 = n9726 & n9727;
  assign n9729 = n9726 | n9727;
  assign n9730 = ~n9728 & n9729;
  assign n14315 = n9535 & n9730;
  assign n14316 = (n9730 & n14224) | (n9730 & n14315) | (n14224 & n14315);
  assign n14317 = n9535 | n9730;
  assign n14318 = n14224 | n14317;
  assign n9733 = ~n14316 & n14318;
  assign n9734 = x66 & x101;
  assign n9735 = n9733 & n9734;
  assign n9736 = n9733 | n9734;
  assign n9737 = ~n9735 & n9736;
  assign n14319 = n9542 & n9737;
  assign n14320 = (n9737 & n14229) | (n9737 & n14319) | (n14229 & n14319);
  assign n14321 = n9542 | n9737;
  assign n14322 = n14229 | n14321;
  assign n9740 = ~n14320 & n14322;
  assign n9741 = x65 & x102;
  assign n9742 = n9740 & n9741;
  assign n9743 = n9740 | n9741;
  assign n9744 = ~n9742 & n9743;
  assign n14247 = n9549 | n9551;
  assign n14323 = n9744 & n14247;
  assign n14324 = n9549 & n9744;
  assign n14325 = (n14156 & n14323) | (n14156 & n14324) | (n14323 & n14324);
  assign n14326 = n9744 | n14247;
  assign n14327 = n9549 | n9744;
  assign n14328 = (n14156 & n14326) | (n14156 & n14327) | (n14326 & n14327);
  assign n9747 = ~n14325 & n14328;
  assign n9748 = x64 & x103;
  assign n9749 = n9747 & n9748;
  assign n9750 = n9747 | n9748;
  assign n9751 = ~n9749 & n9750;
  assign n14245 = n9556 | n9558;
  assign n17034 = n9751 & n14245;
  assign n17035 = n9556 & n9751;
  assign n17036 = (n14154 & n17034) | (n14154 & n17035) | (n17034 & n17035);
  assign n17037 = n9751 | n14245;
  assign n17038 = n9556 | n9751;
  assign n17039 = (n14154 & n17037) | (n14154 & n17038) | (n17037 & n17038);
  assign n9754 = ~n17036 & n17039;
  assign n9755 = x63 & x104;
  assign n9756 = n9754 & n9755;
  assign n9757 = n9754 | n9755;
  assign n9758 = ~n9756 & n9757;
  assign n14243 = n9563 | n9565;
  assign n17040 = n9758 & n14243;
  assign n17041 = n9563 & n9758;
  assign n17042 = (n14152 & n17040) | (n14152 & n17041) | (n17040 & n17041);
  assign n17043 = n9758 | n14243;
  assign n17044 = n9563 | n9758;
  assign n17045 = (n14152 & n17043) | (n14152 & n17044) | (n17043 & n17044);
  assign n9761 = ~n17042 & n17045;
  assign n9762 = x62 & x105;
  assign n9763 = n9761 & n9762;
  assign n9764 = n9761 | n9762;
  assign n9765 = ~n9763 & n9764;
  assign n9766 = n14242 & n9765;
  assign n9767 = n14242 | n9765;
  assign n9768 = ~n9766 & n9767;
  assign n9769 = x61 & x106;
  assign n9770 = n9768 & n9769;
  assign n9771 = n9768 | n9769;
  assign n9772 = ~n9770 & n9771;
  assign n9773 = n14240 & n9772;
  assign n9774 = n14240 | n9772;
  assign n9775 = ~n9773 & n9774;
  assign n9776 = x60 & x107;
  assign n9777 = n9775 & n9776;
  assign n9778 = n9775 | n9776;
  assign n9779 = ~n9777 & n9778;
  assign n9780 = n14238 & n9779;
  assign n9781 = n14238 | n9779;
  assign n9782 = ~n9780 & n9781;
  assign n9783 = x59 & x108;
  assign n9784 = n9782 & n9783;
  assign n9785 = n9782 | n9783;
  assign n9786 = ~n9784 & n9785;
  assign n9787 = n14236 & n9786;
  assign n9788 = n14236 | n9786;
  assign n9789 = ~n9787 & n9788;
  assign n9790 = x58 & x109;
  assign n9791 = n9789 & n9790;
  assign n9792 = n9789 | n9790;
  assign n9793 = ~n9791 & n9792;
  assign n9794 = n14234 & n9793;
  assign n9795 = n14234 | n9793;
  assign n9796 = ~n9794 & n9795;
  assign n9797 = x57 & x110;
  assign n9798 = n9796 & n9797;
  assign n9799 = n9796 | n9797;
  assign n9800 = ~n9798 & n9799;
  assign n9801 = n9619 & n9800;
  assign n9802 = n9619 | n9800;
  assign n9803 = ~n9801 & n9802;
  assign n9804 = x56 & x111;
  assign n9805 = n9803 & n9804;
  assign n9806 = n9803 | n9804;
  assign n9807 = ~n9805 & n9806;
  assign n9808 = n9618 & n9807;
  assign n9809 = n9618 | n9807;
  assign n9810 = ~n9808 & n9809;
  assign n9811 = n9805 | n9808;
  assign n14329 = n9798 | n9800;
  assign n14330 = (n9619 & n9798) | (n9619 & n14329) | (n9798 & n14329);
  assign n14331 = n9791 | n9793;
  assign n14332 = (n9791 & n14234) | (n9791 & n14331) | (n14234 & n14331);
  assign n14333 = n9784 | n9786;
  assign n14334 = (n9784 & n14236) | (n9784 & n14333) | (n14236 & n14333);
  assign n14335 = n9777 | n9779;
  assign n14336 = (n9777 & n14238) | (n9777 & n14335) | (n14238 & n14335);
  assign n14337 = n9770 | n9772;
  assign n14338 = (n9770 & n14240) | (n9770 & n14337) | (n14240 & n14337);
  assign n14244 = (n9563 & n14152) | (n9563 & n14243) | (n14152 & n14243);
  assign n14246 = (n9556 & n14154) | (n9556 & n14245) | (n14154 & n14245);
  assign n14351 = n9672 | n9674;
  assign n17048 = n9479 | n9672;
  assign n17049 = (n9672 & n9674) | (n9672 & n17048) | (n9674 & n17048);
  assign n17050 = (n14194 & n14351) | (n14194 & n17049) | (n14351 & n17049);
  assign n17051 = (n14193 & n14351) | (n14193 & n17049) | (n14351 & n17049);
  assign n17052 = (n16892 & n17050) | (n16892 & n17051) | (n17050 & n17051);
  assign n14356 = n9651 | n9653;
  assign n17053 = n9458 | n9651;
  assign n17054 = (n9651 & n9653) | (n9651 & n17053) | (n9653 & n17053);
  assign n17055 = (n14184 & n14356) | (n14184 & n17054) | (n14356 & n17054);
  assign n17056 = (n14183 & n14356) | (n14183 & n17054) | (n14356 & n17054);
  assign n17057 = (n14073 & n17055) | (n14073 & n17056) | (n17055 & n17056);
  assign n9835 = x79 & x89;
  assign n17829 = n9643 & n9835;
  assign n17969 = n16963 & n17829;
  assign n17970 = n9835 & n17825;
  assign n17971 = n16909 & n17970;
  assign n17833 = (n16901 & n17969) | (n16901 & n17971) | (n17969 & n17971);
  assign n17830 = (n9446 & n17833) | (n9446 & n17829) | (n17833 & n17829);
  assign n17060 = (n14174 & n17830) | (n14174 & n17833) | (n17830 & n17833);
  assign n17061 = (n9835 & n17020) | (n9835 & n17060) | (n17020 & n17060);
  assign n17834 = (n9646 & n9835) | (n9646 & n17060) | (n9835 & n17060);
  assign n18077 = n9835 & n17829;
  assign n18166 = n16963 & n18077;
  assign n18168 = n16909 & n17970;
  assign n18081 = (n16901 & n18166) | (n16901 & n18168) | (n18166 & n18168);
  assign n18078 = (n9446 & n18081) | (n9446 & n18077) | (n18081 & n18077);
  assign n17974 = (n14174 & n18078) | (n14174 & n18081) | (n18078 & n18081);
  assign n17836 = (n9451 & n17834) | (n9451 & n17974) | (n17834 & n17974);
  assign n17063 = (n16959 & n17061) | (n16959 & n17836) | (n17061 & n17836);
  assign n17837 = n9643 | n9835;
  assign n17975 = (n9835 & n16963) | (n9835 & n17837) | (n16963 & n17837);
  assign n17976 = n9835 | n17825;
  assign n17977 = (n9835 & n16909) | (n9835 & n17976) | (n16909 & n17976);
  assign n17841 = (n16901 & n17975) | (n16901 & n17977) | (n17975 & n17977);
  assign n17838 = (n9446 & n17841) | (n9446 & n17837) | (n17841 & n17837);
  assign n17066 = (n14174 & n17838) | (n14174 & n17841) | (n17838 & n17841);
  assign n17067 = n17020 | n17066;
  assign n17842 = n9646 | n17066;
  assign n17843 = (n9451 & n17066) | (n9451 & n17842) | (n17066 & n17842);
  assign n17069 = (n16959 & n17067) | (n16959 & n17843) | (n17067 & n17843);
  assign n9838 = ~n17063 & n17069;
  assign n9839 = n17057 & n9838;
  assign n9840 = n17057 | n9838;
  assign n9841 = ~n9839 & n9840;
  assign n9842 = x78 & x90;
  assign n9843 = n9841 & n9842;
  assign n9844 = n9841 | n9842;
  assign n9845 = ~n9843 & n9844;
  assign n14353 = n9658 | n9660;
  assign n14362 = n9845 & n14353;
  assign n14363 = n9658 & n9845;
  assign n14364 = (n17011 & n14362) | (n17011 & n14363) | (n14362 & n14363);
  assign n14365 = n9845 | n14353;
  assign n14366 = n9658 | n9845;
  assign n14367 = (n17011 & n14365) | (n17011 & n14366) | (n14365 & n14366);
  assign n9848 = ~n14364 & n14367;
  assign n9849 = x77 & x91;
  assign n9850 = n9848 & n9849;
  assign n9851 = n9848 | n9849;
  assign n9852 = ~n9850 & n9851;
  assign n14368 = n9665 & n9852;
  assign n17070 = (n9852 & n14280) | (n9852 & n14368) | (n14280 & n14368);
  assign n17071 = (n9852 & n14279) | (n9852 & n14368) | (n14279 & n14368);
  assign n17072 = (n16954 & n17070) | (n16954 & n17071) | (n17070 & n17071);
  assign n14370 = n9665 | n9852;
  assign n17073 = n14280 | n14370;
  assign n17074 = n14279 | n14370;
  assign n17075 = (n16954 & n17073) | (n16954 & n17074) | (n17073 & n17074);
  assign n9855 = ~n17072 & n17075;
  assign n9856 = x76 & x92;
  assign n9857 = n9855 & n9856;
  assign n9858 = n9855 | n9856;
  assign n9859 = ~n9857 & n9858;
  assign n9860 = n17052 & n9859;
  assign n9861 = n17052 | n9859;
  assign n9862 = ~n9860 & n9861;
  assign n9863 = x75 & x93;
  assign n9864 = n9862 & n9863;
  assign n9865 = n9862 | n9863;
  assign n9866 = ~n9864 & n9865;
  assign n14348 = n9679 | n9681;
  assign n14372 = n9866 & n14348;
  assign n14373 = n9679 & n9866;
  assign n14374 = (n17006 & n14372) | (n17006 & n14373) | (n14372 & n14373);
  assign n14375 = n9866 | n14348;
  assign n14376 = n9679 | n9866;
  assign n14377 = (n17006 & n14375) | (n17006 & n14376) | (n14375 & n14376);
  assign n9869 = ~n14374 & n14377;
  assign n9870 = x74 & x94;
  assign n9871 = n9869 & n9870;
  assign n9872 = n9869 | n9870;
  assign n9873 = ~n9871 & n9872;
  assign n14378 = n9686 & n9873;
  assign n17076 = (n9873 & n14290) | (n9873 & n14378) | (n14290 & n14378);
  assign n17077 = (n9873 & n14289) | (n9873 & n14378) | (n14289 & n14378);
  assign n17078 = (n14161 & n17076) | (n14161 & n17077) | (n17076 & n17077);
  assign n14380 = n9686 | n9873;
  assign n17079 = n14290 | n14380;
  assign n17080 = n14289 | n14380;
  assign n17081 = (n14161 & n17079) | (n14161 & n17080) | (n17079 & n17080);
  assign n9876 = ~n17078 & n17081;
  assign n9877 = x73 & x95;
  assign n9878 = n9876 & n9877;
  assign n9879 = n9876 | n9877;
  assign n9880 = ~n9878 & n9879;
  assign n14346 = n9693 | n9695;
  assign n17082 = n9880 & n14346;
  assign n17046 = n9500 | n9693;
  assign n17047 = (n9693 & n9695) | (n9693 & n17046) | (n9695 & n17046);
  assign n17083 = n9880 & n17047;
  assign n17084 = (n16986 & n17082) | (n16986 & n17083) | (n17082 & n17083);
  assign n17085 = n9880 | n14346;
  assign n17086 = n9880 | n17047;
  assign n17087 = (n16986 & n17085) | (n16986 & n17086) | (n17085 & n17086);
  assign n9883 = ~n17084 & n17087;
  assign n9884 = x72 & x96;
  assign n9885 = n9883 & n9884;
  assign n9886 = n9883 | n9884;
  assign n9887 = ~n9885 & n9886;
  assign n14382 = n9700 & n9887;
  assign n17088 = (n9887 & n14299) | (n9887 & n14382) | (n14299 & n14382);
  assign n17089 = (n9702 & n9887) | (n9702 & n14382) | (n9887 & n14382);
  assign n17090 = (n14208 & n17088) | (n14208 & n17089) | (n17088 & n17089);
  assign n14384 = n9700 | n9887;
  assign n17091 = n14299 | n14384;
  assign n17092 = n9702 | n14384;
  assign n17093 = (n14208 & n17091) | (n14208 & n17092) | (n17091 & n17092);
  assign n9890 = ~n17090 & n17093;
  assign n9891 = x71 & x97;
  assign n9892 = n9890 & n9891;
  assign n9893 = n9890 | n9891;
  assign n9894 = ~n9892 & n9893;
  assign n14386 = n9707 & n9894;
  assign n14387 = (n9894 & n14304) | (n9894 & n14386) | (n14304 & n14386);
  assign n14388 = n9707 | n9894;
  assign n14389 = n14304 | n14388;
  assign n9897 = ~n14387 & n14389;
  assign n9898 = x70 & x98;
  assign n9899 = n9897 & n9898;
  assign n9900 = n9897 | n9898;
  assign n9901 = ~n9899 & n9900;
  assign n14390 = n9714 & n9901;
  assign n14391 = (n9901 & n14308) | (n9901 & n14390) | (n14308 & n14390);
  assign n14392 = n9714 | n9901;
  assign n14393 = n14308 | n14392;
  assign n9904 = ~n14391 & n14393;
  assign n9905 = x69 & x99;
  assign n9906 = n9904 & n9905;
  assign n9907 = n9904 | n9905;
  assign n9908 = ~n9906 & n9907;
  assign n14394 = n9721 & n9908;
  assign n14395 = (n9908 & n14312) | (n9908 & n14394) | (n14312 & n14394);
  assign n14396 = n9721 | n9908;
  assign n14397 = n14312 | n14396;
  assign n9911 = ~n14395 & n14397;
  assign n9912 = x68 & x100;
  assign n9913 = n9911 & n9912;
  assign n9914 = n9911 | n9912;
  assign n9915 = ~n9913 & n9914;
  assign n14398 = n9728 & n9915;
  assign n14399 = (n9915 & n14316) | (n9915 & n14398) | (n14316 & n14398);
  assign n14400 = n9728 | n9915;
  assign n14401 = n14316 | n14400;
  assign n9918 = ~n14399 & n14401;
  assign n9919 = x67 & x101;
  assign n9920 = n9918 & n9919;
  assign n9921 = n9918 | n9919;
  assign n9922 = ~n9920 & n9921;
  assign n14402 = n9735 & n9922;
  assign n14403 = (n9922 & n14320) | (n9922 & n14402) | (n14320 & n14402);
  assign n14404 = n9735 | n9922;
  assign n14405 = n14320 | n14404;
  assign n9925 = ~n14403 & n14405;
  assign n9926 = x66 & x102;
  assign n9927 = n9925 & n9926;
  assign n9928 = n9925 | n9926;
  assign n9929 = ~n9927 & n9928;
  assign n14406 = n9742 & n9929;
  assign n14407 = (n9929 & n14325) | (n9929 & n14406) | (n14325 & n14406);
  assign n14408 = n9742 | n9929;
  assign n14409 = n14325 | n14408;
  assign n9932 = ~n14407 & n14409;
  assign n9933 = x65 & x103;
  assign n9934 = n9932 & n9933;
  assign n9935 = n9932 | n9933;
  assign n9936 = ~n9934 & n9935;
  assign n14343 = n9749 | n9751;
  assign n14410 = n9936 & n14343;
  assign n14411 = n9749 & n9936;
  assign n14412 = (n14246 & n14410) | (n14246 & n14411) | (n14410 & n14411);
  assign n14413 = n9936 | n14343;
  assign n14414 = n9749 | n9936;
  assign n14415 = (n14246 & n14413) | (n14246 & n14414) | (n14413 & n14414);
  assign n9939 = ~n14412 & n14415;
  assign n9940 = x64 & x104;
  assign n9941 = n9939 & n9940;
  assign n9942 = n9939 | n9940;
  assign n9943 = ~n9941 & n9942;
  assign n14341 = n9756 | n9758;
  assign n17094 = n9943 & n14341;
  assign n17095 = n9756 & n9943;
  assign n17096 = (n14244 & n17094) | (n14244 & n17095) | (n17094 & n17095);
  assign n17097 = n9943 | n14341;
  assign n17098 = n9756 | n9943;
  assign n17099 = (n14244 & n17097) | (n14244 & n17098) | (n17097 & n17098);
  assign n9946 = ~n17096 & n17099;
  assign n9947 = x63 & x105;
  assign n9948 = n9946 & n9947;
  assign n9949 = n9946 | n9947;
  assign n9950 = ~n9948 & n9949;
  assign n14339 = n9763 | n9765;
  assign n17100 = n9950 & n14339;
  assign n17101 = n9763 & n9950;
  assign n17102 = (n14242 & n17100) | (n14242 & n17101) | (n17100 & n17101);
  assign n17103 = n9950 | n14339;
  assign n17104 = n9763 | n9950;
  assign n17105 = (n14242 & n17103) | (n14242 & n17104) | (n17103 & n17104);
  assign n9953 = ~n17102 & n17105;
  assign n9954 = x62 & x106;
  assign n9955 = n9953 & n9954;
  assign n9956 = n9953 | n9954;
  assign n9957 = ~n9955 & n9956;
  assign n9958 = n14338 & n9957;
  assign n9959 = n14338 | n9957;
  assign n9960 = ~n9958 & n9959;
  assign n9961 = x61 & x107;
  assign n9962 = n9960 & n9961;
  assign n9963 = n9960 | n9961;
  assign n9964 = ~n9962 & n9963;
  assign n9965 = n14336 & n9964;
  assign n9966 = n14336 | n9964;
  assign n9967 = ~n9965 & n9966;
  assign n9968 = x60 & x108;
  assign n9969 = n9967 & n9968;
  assign n9970 = n9967 | n9968;
  assign n9971 = ~n9969 & n9970;
  assign n9972 = n14334 & n9971;
  assign n9973 = n14334 | n9971;
  assign n9974 = ~n9972 & n9973;
  assign n9975 = x59 & x109;
  assign n9976 = n9974 & n9975;
  assign n9977 = n9974 | n9975;
  assign n9978 = ~n9976 & n9977;
  assign n9979 = n14332 & n9978;
  assign n9980 = n14332 | n9978;
  assign n9981 = ~n9979 & n9980;
  assign n9982 = x58 & x110;
  assign n9983 = n9981 & n9982;
  assign n9984 = n9981 | n9982;
  assign n9985 = ~n9983 & n9984;
  assign n9986 = n14330 & n9985;
  assign n9987 = n14330 | n9985;
  assign n9988 = ~n9986 & n9987;
  assign n9989 = x57 & x111;
  assign n9990 = n9988 & n9989;
  assign n9991 = n9988 | n9989;
  assign n9992 = ~n9990 & n9991;
  assign n9993 = n9811 & n9992;
  assign n9994 = n9811 | n9992;
  assign n9995 = ~n9993 & n9994;
  assign n14416 = n9990 | n9992;
  assign n14417 = (n9811 & n9990) | (n9811 & n14416) | (n9990 & n14416);
  assign n14418 = n9983 | n9985;
  assign n14419 = (n9983 & n14330) | (n9983 & n14418) | (n14330 & n14418);
  assign n14420 = n9976 | n9978;
  assign n14421 = (n9976 & n14332) | (n9976 & n14420) | (n14332 & n14420);
  assign n14422 = n9969 | n9971;
  assign n14423 = (n9969 & n14334) | (n9969 & n14422) | (n14334 & n14422);
  assign n14424 = n9962 | n9964;
  assign n14425 = (n9962 & n14336) | (n9962 & n14424) | (n14336 & n14424);
  assign n14340 = (n9763 & n14242) | (n9763 & n14339) | (n14242 & n14339);
  assign n14342 = (n9756 & n14244) | (n9756 & n14341) | (n14244 & n14341);
  assign n14347 = (n16986 & n17047) | (n16986 & n14346) | (n17047 & n14346);
  assign n14435 = n9871 | n9873;
  assign n17106 = n9686 | n9871;
  assign n17107 = (n9871 & n9873) | (n9871 & n17106) | (n9873 & n17106);
  assign n17108 = (n14290 & n14435) | (n14290 & n17107) | (n14435 & n17107);
  assign n17109 = (n14289 & n14435) | (n14289 & n17107) | (n14435 & n17107);
  assign n17110 = (n14161 & n17108) | (n14161 & n17109) | (n17108 & n17109);
  assign n14440 = n9850 | n9852;
  assign n17111 = n9665 | n9850;
  assign n17112 = (n9850 & n9852) | (n9850 & n17111) | (n9852 & n17111);
  assign n17113 = (n14280 & n14440) | (n14280 & n17112) | (n14440 & n17112);
  assign n17114 = (n14279 & n14440) | (n14279 & n17112) | (n14440 & n17112);
  assign n17115 = (n16954 & n17113) | (n16954 & n17114) | (n17113 & n17114);
  assign n10019 = x79 & x90;
  assign n17116 = n10019 & n17063;
  assign n17117 = (n9838 & n10019) | (n9838 & n17116) | (n10019 & n17116);
  assign n14445 = n10019 & n17063;
  assign n14446 = (n17057 & n17117) | (n17057 & n14445) | (n17117 & n14445);
  assign n17118 = n10019 | n17063;
  assign n17119 = n9838 | n17118;
  assign n14448 = n10019 | n17063;
  assign n14449 = (n17057 & n17119) | (n17057 & n14448) | (n17119 & n14448);
  assign n10022 = ~n14446 & n14449;
  assign n14450 = n9843 & n10022;
  assign n17120 = (n10022 & n14363) | (n10022 & n14450) | (n14363 & n14450);
  assign n17121 = (n10022 & n14362) | (n10022 & n14450) | (n14362 & n14450);
  assign n17122 = (n17011 & n17120) | (n17011 & n17121) | (n17120 & n17121);
  assign n14452 = n9843 | n10022;
  assign n17123 = n14363 | n14452;
  assign n17124 = n14362 | n14452;
  assign n17125 = (n17011 & n17123) | (n17011 & n17124) | (n17123 & n17124);
  assign n10025 = ~n17122 & n17125;
  assign n10026 = x78 & x91;
  assign n10027 = n10025 & n10026;
  assign n10028 = n10025 | n10026;
  assign n10029 = ~n10027 & n10028;
  assign n10030 = n17115 & n10029;
  assign n10031 = n17115 | n10029;
  assign n10032 = ~n10030 & n10031;
  assign n10033 = x77 & x92;
  assign n10034 = n10032 & n10033;
  assign n10035 = n10032 | n10033;
  assign n10036 = ~n10034 & n10035;
  assign n14437 = n9857 | n9859;
  assign n14454 = n10036 & n14437;
  assign n14455 = n9857 & n10036;
  assign n14456 = (n17052 & n14454) | (n17052 & n14455) | (n14454 & n14455);
  assign n14457 = n10036 | n14437;
  assign n14458 = n9857 | n10036;
  assign n14459 = (n17052 & n14457) | (n17052 & n14458) | (n14457 & n14458);
  assign n10039 = ~n14456 & n14459;
  assign n10040 = x76 & x93;
  assign n10041 = n10039 & n10040;
  assign n10042 = n10039 | n10040;
  assign n10043 = ~n10041 & n10042;
  assign n14460 = n9864 & n10043;
  assign n17126 = (n10043 & n14373) | (n10043 & n14460) | (n14373 & n14460);
  assign n17127 = (n10043 & n14372) | (n10043 & n14460) | (n14372 & n14460);
  assign n17128 = (n17006 & n17126) | (n17006 & n17127) | (n17126 & n17127);
  assign n14462 = n9864 | n10043;
  assign n17129 = n14373 | n14462;
  assign n17130 = n14372 | n14462;
  assign n17131 = (n17006 & n17129) | (n17006 & n17130) | (n17129 & n17130);
  assign n10046 = ~n17128 & n17131;
  assign n10047 = x75 & x94;
  assign n10048 = n10046 & n10047;
  assign n10049 = n10046 | n10047;
  assign n10050 = ~n10048 & n10049;
  assign n10051 = n17110 & n10050;
  assign n10052 = n17110 | n10050;
  assign n10053 = ~n10051 & n10052;
  assign n10054 = x74 & x95;
  assign n10055 = n10053 & n10054;
  assign n10056 = n10053 | n10054;
  assign n10057 = ~n10055 & n10056;
  assign n14432 = n9878 | n9880;
  assign n14464 = n10057 & n14432;
  assign n14465 = n9878 & n10057;
  assign n14466 = (n14347 & n14464) | (n14347 & n14465) | (n14464 & n14465);
  assign n14467 = n10057 | n14432;
  assign n14468 = n9878 | n10057;
  assign n14469 = (n14347 & n14467) | (n14347 & n14468) | (n14467 & n14468);
  assign n10060 = ~n14466 & n14469;
  assign n10061 = x73 & x96;
  assign n10062 = n10060 & n10061;
  assign n10063 = n10060 | n10061;
  assign n10064 = ~n10062 & n10063;
  assign n14470 = n9885 & n10064;
  assign n14471 = (n10064 & n17090) | (n10064 & n14470) | (n17090 & n14470);
  assign n14472 = n9885 | n10064;
  assign n14473 = n17090 | n14472;
  assign n10067 = ~n14471 & n14473;
  assign n10068 = x72 & x97;
  assign n10069 = n10067 & n10068;
  assign n10070 = n10067 | n10068;
  assign n10071 = ~n10069 & n10070;
  assign n14474 = n9892 & n10071;
  assign n14475 = (n10071 & n14387) | (n10071 & n14474) | (n14387 & n14474);
  assign n14476 = n9892 | n10071;
  assign n14477 = n14387 | n14476;
  assign n10074 = ~n14475 & n14477;
  assign n10075 = x71 & x98;
  assign n10076 = n10074 & n10075;
  assign n10077 = n10074 | n10075;
  assign n10078 = ~n10076 & n10077;
  assign n14478 = n9899 & n10078;
  assign n14479 = (n10078 & n14391) | (n10078 & n14478) | (n14391 & n14478);
  assign n14480 = n9899 | n10078;
  assign n14481 = n14391 | n14480;
  assign n10081 = ~n14479 & n14481;
  assign n10082 = x70 & x99;
  assign n10083 = n10081 & n10082;
  assign n10084 = n10081 | n10082;
  assign n10085 = ~n10083 & n10084;
  assign n14482 = n9906 & n10085;
  assign n14483 = (n10085 & n14395) | (n10085 & n14482) | (n14395 & n14482);
  assign n14484 = n9906 | n10085;
  assign n14485 = n14395 | n14484;
  assign n10088 = ~n14483 & n14485;
  assign n10089 = x69 & x100;
  assign n10090 = n10088 & n10089;
  assign n10091 = n10088 | n10089;
  assign n10092 = ~n10090 & n10091;
  assign n14486 = n9913 & n10092;
  assign n14487 = (n10092 & n14399) | (n10092 & n14486) | (n14399 & n14486);
  assign n14488 = n9913 | n10092;
  assign n14489 = n14399 | n14488;
  assign n10095 = ~n14487 & n14489;
  assign n10096 = x68 & x101;
  assign n10097 = n10095 & n10096;
  assign n10098 = n10095 | n10096;
  assign n10099 = ~n10097 & n10098;
  assign n14490 = n9920 & n10099;
  assign n14491 = (n10099 & n14403) | (n10099 & n14490) | (n14403 & n14490);
  assign n14492 = n9920 | n10099;
  assign n14493 = n14403 | n14492;
  assign n10102 = ~n14491 & n14493;
  assign n10103 = x67 & x102;
  assign n10104 = n10102 & n10103;
  assign n10105 = n10102 | n10103;
  assign n10106 = ~n10104 & n10105;
  assign n14494 = n9927 & n10106;
  assign n14495 = (n10106 & n14407) | (n10106 & n14494) | (n14407 & n14494);
  assign n14496 = n9927 | n10106;
  assign n14497 = n14407 | n14496;
  assign n10109 = ~n14495 & n14497;
  assign n10110 = x66 & x103;
  assign n10111 = n10109 & n10110;
  assign n10112 = n10109 | n10110;
  assign n10113 = ~n10111 & n10112;
  assign n14498 = n9934 & n10113;
  assign n14499 = (n10113 & n14412) | (n10113 & n14498) | (n14412 & n14498);
  assign n14500 = n9934 | n10113;
  assign n14501 = n14412 | n14500;
  assign n10116 = ~n14499 & n14501;
  assign n10117 = x65 & x104;
  assign n10118 = n10116 & n10117;
  assign n10119 = n10116 | n10117;
  assign n10120 = ~n10118 & n10119;
  assign n14430 = n9941 | n9943;
  assign n14502 = n10120 & n14430;
  assign n14503 = n9941 & n10120;
  assign n14504 = (n14342 & n14502) | (n14342 & n14503) | (n14502 & n14503);
  assign n14505 = n10120 | n14430;
  assign n14506 = n9941 | n10120;
  assign n14507 = (n14342 & n14505) | (n14342 & n14506) | (n14505 & n14506);
  assign n10123 = ~n14504 & n14507;
  assign n10124 = x64 & x105;
  assign n10125 = n10123 & n10124;
  assign n10126 = n10123 | n10124;
  assign n10127 = ~n10125 & n10126;
  assign n14428 = n9948 | n9950;
  assign n17132 = n10127 & n14428;
  assign n17133 = n9948 & n10127;
  assign n17134 = (n14340 & n17132) | (n14340 & n17133) | (n17132 & n17133);
  assign n17135 = n10127 | n14428;
  assign n17136 = n9948 | n10127;
  assign n17137 = (n14340 & n17135) | (n14340 & n17136) | (n17135 & n17136);
  assign n10130 = ~n17134 & n17137;
  assign n10131 = x63 & x106;
  assign n10132 = n10130 & n10131;
  assign n10133 = n10130 | n10131;
  assign n10134 = ~n10132 & n10133;
  assign n14426 = n9955 | n9957;
  assign n17138 = n10134 & n14426;
  assign n17139 = n9955 & n10134;
  assign n17140 = (n14338 & n17138) | (n14338 & n17139) | (n17138 & n17139);
  assign n17141 = n10134 | n14426;
  assign n17142 = n9955 | n10134;
  assign n17143 = (n14338 & n17141) | (n14338 & n17142) | (n17141 & n17142);
  assign n10137 = ~n17140 & n17143;
  assign n10138 = x62 & x107;
  assign n10139 = n10137 & n10138;
  assign n10140 = n10137 | n10138;
  assign n10141 = ~n10139 & n10140;
  assign n10142 = n14425 & n10141;
  assign n10143 = n14425 | n10141;
  assign n10144 = ~n10142 & n10143;
  assign n10145 = x61 & x108;
  assign n10146 = n10144 & n10145;
  assign n10147 = n10144 | n10145;
  assign n10148 = ~n10146 & n10147;
  assign n10149 = n14423 & n10148;
  assign n10150 = n14423 | n10148;
  assign n10151 = ~n10149 & n10150;
  assign n10152 = x60 & x109;
  assign n10153 = n10151 & n10152;
  assign n10154 = n10151 | n10152;
  assign n10155 = ~n10153 & n10154;
  assign n10156 = n14421 & n10155;
  assign n10157 = n14421 | n10155;
  assign n10158 = ~n10156 & n10157;
  assign n10159 = x59 & x110;
  assign n10160 = n10158 & n10159;
  assign n10161 = n10158 | n10159;
  assign n10162 = ~n10160 & n10161;
  assign n10163 = n14419 & n10162;
  assign n10164 = n14419 | n10162;
  assign n10165 = ~n10163 & n10164;
  assign n10166 = x58 & x111;
  assign n10167 = n10165 & n10166;
  assign n10168 = n10165 | n10166;
  assign n10169 = ~n10167 & n10168;
  assign n10170 = n14417 & n10169;
  assign n10171 = n14417 | n10169;
  assign n10172 = ~n10170 & n10171;
  assign n14508 = n10167 | n10169;
  assign n14509 = (n10167 & n14417) | (n10167 & n14508) | (n14417 & n14508);
  assign n14510 = n10160 | n10162;
  assign n14511 = (n10160 & n14419) | (n10160 & n14510) | (n14419 & n14510);
  assign n14512 = n10153 | n10155;
  assign n14513 = (n10153 & n14421) | (n10153 & n14512) | (n14421 & n14512);
  assign n14514 = n10146 | n10148;
  assign n14515 = (n10146 & n14423) | (n10146 & n14514) | (n14423 & n14514);
  assign n14427 = (n9955 & n14338) | (n9955 & n14426) | (n14338 & n14426);
  assign n14429 = (n9948 & n14340) | (n9948 & n14428) | (n14340 & n14428);
  assign n14528 = n10041 | n10043;
  assign n17146 = n9864 | n10041;
  assign n17147 = (n10041 & n10043) | (n10041 & n17146) | (n10043 & n17146);
  assign n17148 = (n14373 & n14528) | (n14373 & n17147) | (n14528 & n17147);
  assign n17149 = (n14372 & n14528) | (n14372 & n17147) | (n14528 & n17147);
  assign n17150 = (n17006 & n17148) | (n17006 & n17149) | (n17148 & n17149);
  assign n10195 = x79 & x91;
  assign n14533 = n10022 | n14446;
  assign n17151 = (n9843 & n14446) | (n9843 & n14533) | (n14446 & n14533);
  assign n14535 = n10195 & n17151;
  assign n17844 = n10195 & n17117;
  assign n17978 = n10019 & n10195;
  assign n17979 = n17063 & n17978;
  assign n17846 = (n17057 & n17844) | (n17057 & n17979) | (n17844 & n17979);
  assign n17153 = (n10022 & n10195) | (n10022 & n17846) | (n10195 & n17846);
  assign n17154 = (n14363 & n14535) | (n14363 & n17153) | (n14535 & n17153);
  assign n17155 = (n14362 & n14535) | (n14362 & n17153) | (n14535 & n17153);
  assign n17156 = (n17011 & n17154) | (n17011 & n17155) | (n17154 & n17155);
  assign n14538 = n10195 | n17151;
  assign n17847 = n10195 | n17117;
  assign n17980 = n10019 | n10195;
  assign n17981 = (n10195 & n17063) | (n10195 & n17980) | (n17063 & n17980);
  assign n17849 = (n17057 & n17847) | (n17057 & n17981) | (n17847 & n17981);
  assign n17158 = n10022 | n17849;
  assign n17159 = (n14363 & n14538) | (n14363 & n17158) | (n14538 & n17158);
  assign n17160 = (n14362 & n14538) | (n14362 & n17158) | (n14538 & n17158);
  assign n17161 = (n17011 & n17159) | (n17011 & n17160) | (n17159 & n17160);
  assign n10198 = ~n17156 & n17161;
  assign n14542 = n10027 & n10198;
  assign n17162 = (n10029 & n10198) | (n10029 & n14542) | (n10198 & n14542);
  assign n14543 = (n17115 & n17162) | (n17115 & n14542) | (n17162 & n14542);
  assign n14545 = n10027 | n10198;
  assign n17163 = n10029 | n14545;
  assign n14546 = (n17115 & n17163) | (n17115 & n14545) | (n17163 & n14545);
  assign n10201 = ~n14543 & n14546;
  assign n10202 = x78 & x92;
  assign n10203 = n10201 & n10202;
  assign n10204 = n10201 | n10202;
  assign n10205 = ~n10203 & n10204;
  assign n14547 = n10034 & n10205;
  assign n17164 = (n10205 & n14455) | (n10205 & n14547) | (n14455 & n14547);
  assign n17165 = (n10205 & n14454) | (n10205 & n14547) | (n14454 & n14547);
  assign n17166 = (n17052 & n17164) | (n17052 & n17165) | (n17164 & n17165);
  assign n14549 = n10034 | n10205;
  assign n17167 = n14455 | n14549;
  assign n17168 = n14454 | n14549;
  assign n17169 = (n17052 & n17167) | (n17052 & n17168) | (n17167 & n17168);
  assign n10208 = ~n17166 & n17169;
  assign n10209 = x77 & x93;
  assign n10210 = n10208 & n10209;
  assign n10211 = n10208 | n10209;
  assign n10212 = ~n10210 & n10211;
  assign n10213 = n17150 & n10212;
  assign n10214 = n17150 | n10212;
  assign n10215 = ~n10213 & n10214;
  assign n10216 = x76 & x94;
  assign n10217 = n10215 & n10216;
  assign n10218 = n10215 | n10216;
  assign n10219 = ~n10217 & n10218;
  assign n14525 = n10048 | n10050;
  assign n14551 = n10219 & n14525;
  assign n14552 = n10048 & n10219;
  assign n14553 = (n17110 & n14551) | (n17110 & n14552) | (n14551 & n14552);
  assign n14554 = n10219 | n14525;
  assign n14555 = n10048 | n10219;
  assign n14556 = (n17110 & n14554) | (n17110 & n14555) | (n14554 & n14555);
  assign n10222 = ~n14553 & n14556;
  assign n10223 = x75 & x95;
  assign n10224 = n10222 & n10223;
  assign n10225 = n10222 | n10223;
  assign n10226 = ~n10224 & n10225;
  assign n14557 = n10055 & n10226;
  assign n17170 = (n10226 & n14465) | (n10226 & n14557) | (n14465 & n14557);
  assign n17171 = (n10226 & n14464) | (n10226 & n14557) | (n14464 & n14557);
  assign n17172 = (n14347 & n17170) | (n14347 & n17171) | (n17170 & n17171);
  assign n14559 = n10055 | n10226;
  assign n17173 = n14465 | n14559;
  assign n17174 = n14464 | n14559;
  assign n17175 = (n14347 & n17173) | (n14347 & n17174) | (n17173 & n17174);
  assign n10229 = ~n17172 & n17175;
  assign n10230 = x74 & x96;
  assign n10231 = n10229 & n10230;
  assign n10232 = n10229 | n10230;
  assign n10233 = ~n10231 & n10232;
  assign n14523 = n10062 | n10064;
  assign n17176 = n10233 & n14523;
  assign n17144 = n9885 | n10062;
  assign n17145 = (n10062 & n10064) | (n10062 & n17144) | (n10064 & n17144);
  assign n17177 = n10233 & n17145;
  assign n17178 = (n17090 & n17176) | (n17090 & n17177) | (n17176 & n17177);
  assign n17179 = n10233 | n14523;
  assign n17180 = n10233 | n17145;
  assign n17181 = (n17090 & n17179) | (n17090 & n17180) | (n17179 & n17180);
  assign n10236 = ~n17178 & n17181;
  assign n10237 = x73 & x97;
  assign n10238 = n10236 & n10237;
  assign n10239 = n10236 | n10237;
  assign n10240 = ~n10238 & n10239;
  assign n14561 = n10069 & n10240;
  assign n17182 = (n10240 & n14474) | (n10240 & n14561) | (n14474 & n14561);
  assign n17183 = (n10071 & n10240) | (n10071 & n14561) | (n10240 & n14561);
  assign n17184 = (n14387 & n17182) | (n14387 & n17183) | (n17182 & n17183);
  assign n14563 = n10069 | n10240;
  assign n17185 = n14474 | n14563;
  assign n17186 = n10071 | n14563;
  assign n17187 = (n14387 & n17185) | (n14387 & n17186) | (n17185 & n17186);
  assign n10243 = ~n17184 & n17187;
  assign n10244 = x72 & x98;
  assign n10245 = n10243 & n10244;
  assign n10246 = n10243 | n10244;
  assign n10247 = ~n10245 & n10246;
  assign n14565 = n10076 & n10247;
  assign n14566 = (n10247 & n14479) | (n10247 & n14565) | (n14479 & n14565);
  assign n14567 = n10076 | n10247;
  assign n14568 = n14479 | n14567;
  assign n10250 = ~n14566 & n14568;
  assign n10251 = x71 & x99;
  assign n10252 = n10250 & n10251;
  assign n10253 = n10250 | n10251;
  assign n10254 = ~n10252 & n10253;
  assign n14569 = n10083 & n10254;
  assign n14570 = (n10254 & n14483) | (n10254 & n14569) | (n14483 & n14569);
  assign n14571 = n10083 | n10254;
  assign n14572 = n14483 | n14571;
  assign n10257 = ~n14570 & n14572;
  assign n10258 = x70 & x100;
  assign n10259 = n10257 & n10258;
  assign n10260 = n10257 | n10258;
  assign n10261 = ~n10259 & n10260;
  assign n14573 = n10090 & n10261;
  assign n14574 = (n10261 & n14487) | (n10261 & n14573) | (n14487 & n14573);
  assign n14575 = n10090 | n10261;
  assign n14576 = n14487 | n14575;
  assign n10264 = ~n14574 & n14576;
  assign n10265 = x69 & x101;
  assign n10266 = n10264 & n10265;
  assign n10267 = n10264 | n10265;
  assign n10268 = ~n10266 & n10267;
  assign n14577 = n10097 & n10268;
  assign n14578 = (n10268 & n14491) | (n10268 & n14577) | (n14491 & n14577);
  assign n14579 = n10097 | n10268;
  assign n14580 = n14491 | n14579;
  assign n10271 = ~n14578 & n14580;
  assign n10272 = x68 & x102;
  assign n10273 = n10271 & n10272;
  assign n10274 = n10271 | n10272;
  assign n10275 = ~n10273 & n10274;
  assign n14581 = n10104 & n10275;
  assign n14582 = (n10275 & n14495) | (n10275 & n14581) | (n14495 & n14581);
  assign n14583 = n10104 | n10275;
  assign n14584 = n14495 | n14583;
  assign n10278 = ~n14582 & n14584;
  assign n10279 = x67 & x103;
  assign n10280 = n10278 & n10279;
  assign n10281 = n10278 | n10279;
  assign n10282 = ~n10280 & n10281;
  assign n14585 = n10111 & n10282;
  assign n14586 = (n10282 & n14499) | (n10282 & n14585) | (n14499 & n14585);
  assign n14587 = n10111 | n10282;
  assign n14588 = n14499 | n14587;
  assign n10285 = ~n14586 & n14588;
  assign n10286 = x66 & x104;
  assign n10287 = n10285 & n10286;
  assign n10288 = n10285 | n10286;
  assign n10289 = ~n10287 & n10288;
  assign n14589 = n10118 & n10289;
  assign n14590 = (n10289 & n14504) | (n10289 & n14589) | (n14504 & n14589);
  assign n14591 = n10118 | n10289;
  assign n14592 = n14504 | n14591;
  assign n10292 = ~n14590 & n14592;
  assign n10293 = x65 & x105;
  assign n10294 = n10292 & n10293;
  assign n10295 = n10292 | n10293;
  assign n10296 = ~n10294 & n10295;
  assign n14520 = n10125 | n10127;
  assign n14593 = n10296 & n14520;
  assign n14594 = n10125 & n10296;
  assign n14595 = (n14429 & n14593) | (n14429 & n14594) | (n14593 & n14594);
  assign n14596 = n10296 | n14520;
  assign n14597 = n10125 | n10296;
  assign n14598 = (n14429 & n14596) | (n14429 & n14597) | (n14596 & n14597);
  assign n10299 = ~n14595 & n14598;
  assign n10300 = x64 & x106;
  assign n10301 = n10299 & n10300;
  assign n10302 = n10299 | n10300;
  assign n10303 = ~n10301 & n10302;
  assign n14518 = n10132 | n10134;
  assign n17188 = n10303 & n14518;
  assign n17189 = n10132 & n10303;
  assign n17190 = (n14427 & n17188) | (n14427 & n17189) | (n17188 & n17189);
  assign n17191 = n10303 | n14518;
  assign n17192 = n10132 | n10303;
  assign n17193 = (n14427 & n17191) | (n14427 & n17192) | (n17191 & n17192);
  assign n10306 = ~n17190 & n17193;
  assign n10307 = x63 & x107;
  assign n10308 = n10306 & n10307;
  assign n10309 = n10306 | n10307;
  assign n10310 = ~n10308 & n10309;
  assign n14516 = n10139 | n10141;
  assign n17194 = n10310 & n14516;
  assign n17195 = n10139 & n10310;
  assign n17196 = (n14425 & n17194) | (n14425 & n17195) | (n17194 & n17195);
  assign n17197 = n10310 | n14516;
  assign n17198 = n10139 | n10310;
  assign n17199 = (n14425 & n17197) | (n14425 & n17198) | (n17197 & n17198);
  assign n10313 = ~n17196 & n17199;
  assign n10314 = x62 & x108;
  assign n10315 = n10313 & n10314;
  assign n10316 = n10313 | n10314;
  assign n10317 = ~n10315 & n10316;
  assign n10318 = n14515 & n10317;
  assign n10319 = n14515 | n10317;
  assign n10320 = ~n10318 & n10319;
  assign n10321 = x61 & x109;
  assign n10322 = n10320 & n10321;
  assign n10323 = n10320 | n10321;
  assign n10324 = ~n10322 & n10323;
  assign n10325 = n14513 & n10324;
  assign n10326 = n14513 | n10324;
  assign n10327 = ~n10325 & n10326;
  assign n10328 = x60 & x110;
  assign n10329 = n10327 & n10328;
  assign n10330 = n10327 | n10328;
  assign n10331 = ~n10329 & n10330;
  assign n10332 = n14511 & n10331;
  assign n10333 = n14511 | n10331;
  assign n10334 = ~n10332 & n10333;
  assign n10335 = x59 & x111;
  assign n10336 = n10334 & n10335;
  assign n10337 = n10334 | n10335;
  assign n10338 = ~n10336 & n10337;
  assign n10339 = n14509 & n10338;
  assign n10340 = n14509 | n10338;
  assign n10341 = ~n10339 & n10340;
  assign n14599 = n10336 | n10338;
  assign n14600 = (n10336 & n14509) | (n10336 & n14599) | (n14509 & n14599);
  assign n14601 = n10329 | n10331;
  assign n14602 = (n10329 & n14511) | (n10329 & n14601) | (n14511 & n14601);
  assign n14603 = n10322 | n10324;
  assign n14604 = (n10322 & n14513) | (n10322 & n14603) | (n14513 & n14603);
  assign n14517 = (n10139 & n14425) | (n10139 & n14516) | (n14425 & n14516);
  assign n14519 = (n10132 & n14427) | (n10132 & n14518) | (n14427 & n14518);
  assign n14524 = (n17090 & n17145) | (n17090 & n14523) | (n17145 & n14523);
  assign n14614 = n10224 | n10226;
  assign n17200 = n10055 | n10224;
  assign n17201 = (n10224 & n10226) | (n10224 & n17200) | (n10226 & n17200);
  assign n17202 = (n14465 & n14614) | (n14465 & n17201) | (n14614 & n17201);
  assign n17203 = (n14464 & n14614) | (n14464 & n17201) | (n14614 & n17201);
  assign n17204 = (n14347 & n17202) | (n14347 & n17203) | (n17202 & n17203);
  assign n14619 = n10203 | n10205;
  assign n17205 = n10034 | n10203;
  assign n17206 = (n10203 & n10205) | (n10203 & n17205) | (n10205 & n17205);
  assign n17207 = (n14455 & n14619) | (n14455 & n17206) | (n14619 & n17206);
  assign n17208 = (n14454 & n14619) | (n14454 & n17206) | (n14619 & n17206);
  assign n17209 = (n17052 & n17207) | (n17052 & n17208) | (n17207 & n17208);
  assign n10363 = x79 & x92;
  assign n14621 = n10363 & n17156;
  assign n17210 = (n10363 & n14621) | (n10363 & n17162) | (n14621 & n17162);
  assign n17850 = (n10198 & n10363) | (n10198 & n14621) | (n10363 & n14621);
  assign n17982 = n10363 & n17156;
  assign n17852 = (n10027 & n17850) | (n10027 & n17982) | (n17850 & n17982);
  assign n17212 = (n17115 & n17210) | (n17115 & n17852) | (n17210 & n17852);
  assign n14623 = n10363 | n17156;
  assign n17213 = n14623 | n17162;
  assign n17853 = n10198 | n14623;
  assign n17854 = (n10027 & n14623) | (n10027 & n17853) | (n14623 & n17853);
  assign n17215 = (n17115 & n17213) | (n17115 & n17854) | (n17213 & n17854);
  assign n10366 = ~n17212 & n17215;
  assign n10367 = n17209 & n10366;
  assign n10368 = n17209 | n10366;
  assign n10369 = ~n10367 & n10368;
  assign n10370 = x78 & x93;
  assign n10371 = n10369 & n10370;
  assign n10372 = n10369 | n10370;
  assign n10373 = ~n10371 & n10372;
  assign n14616 = n10210 | n10212;
  assign n14625 = n10373 & n14616;
  assign n14626 = n10210 & n10373;
  assign n14627 = (n17150 & n14625) | (n17150 & n14626) | (n14625 & n14626);
  assign n14628 = n10373 | n14616;
  assign n14629 = n10210 | n10373;
  assign n14630 = (n17150 & n14628) | (n17150 & n14629) | (n14628 & n14629);
  assign n10376 = ~n14627 & n14630;
  assign n10377 = x77 & x94;
  assign n10378 = n10376 & n10377;
  assign n10379 = n10376 | n10377;
  assign n10380 = ~n10378 & n10379;
  assign n14631 = n10217 & n10380;
  assign n17216 = (n10380 & n14552) | (n10380 & n14631) | (n14552 & n14631);
  assign n17217 = (n10380 & n14551) | (n10380 & n14631) | (n14551 & n14631);
  assign n17218 = (n17110 & n17216) | (n17110 & n17217) | (n17216 & n17217);
  assign n14633 = n10217 | n10380;
  assign n17219 = n14552 | n14633;
  assign n17220 = n14551 | n14633;
  assign n17221 = (n17110 & n17219) | (n17110 & n17220) | (n17219 & n17220);
  assign n10383 = ~n17218 & n17221;
  assign n10384 = x76 & x95;
  assign n10385 = n10383 & n10384;
  assign n10386 = n10383 | n10384;
  assign n10387 = ~n10385 & n10386;
  assign n10388 = n17204 & n10387;
  assign n10389 = n17204 | n10387;
  assign n10390 = ~n10388 & n10389;
  assign n10391 = x75 & x96;
  assign n10392 = n10390 & n10391;
  assign n10393 = n10390 | n10391;
  assign n10394 = ~n10392 & n10393;
  assign n14611 = n10231 | n10233;
  assign n14635 = n10394 & n14611;
  assign n14636 = n10231 & n10394;
  assign n14637 = (n14524 & n14635) | (n14524 & n14636) | (n14635 & n14636);
  assign n14638 = n10394 | n14611;
  assign n14639 = n10231 | n10394;
  assign n14640 = (n14524 & n14638) | (n14524 & n14639) | (n14638 & n14639);
  assign n10397 = ~n14637 & n14640;
  assign n10398 = x74 & x97;
  assign n10399 = n10397 & n10398;
  assign n10400 = n10397 | n10398;
  assign n10401 = ~n10399 & n10400;
  assign n14641 = n10238 & n10401;
  assign n14642 = (n10401 & n17184) | (n10401 & n14641) | (n17184 & n14641);
  assign n14643 = n10238 | n10401;
  assign n14644 = n17184 | n14643;
  assign n10404 = ~n14642 & n14644;
  assign n10405 = x73 & x98;
  assign n10406 = n10404 & n10405;
  assign n10407 = n10404 | n10405;
  assign n10408 = ~n10406 & n10407;
  assign n14645 = n10245 & n10408;
  assign n14646 = (n10408 & n14566) | (n10408 & n14645) | (n14566 & n14645);
  assign n14647 = n10245 | n10408;
  assign n14648 = n14566 | n14647;
  assign n10411 = ~n14646 & n14648;
  assign n10412 = x72 & x99;
  assign n10413 = n10411 & n10412;
  assign n10414 = n10411 | n10412;
  assign n10415 = ~n10413 & n10414;
  assign n14649 = n10252 & n10415;
  assign n14650 = (n10415 & n14570) | (n10415 & n14649) | (n14570 & n14649);
  assign n14651 = n10252 | n10415;
  assign n14652 = n14570 | n14651;
  assign n10418 = ~n14650 & n14652;
  assign n10419 = x71 & x100;
  assign n10420 = n10418 & n10419;
  assign n10421 = n10418 | n10419;
  assign n10422 = ~n10420 & n10421;
  assign n14653 = n10259 & n10422;
  assign n14654 = (n10422 & n14574) | (n10422 & n14653) | (n14574 & n14653);
  assign n14655 = n10259 | n10422;
  assign n14656 = n14574 | n14655;
  assign n10425 = ~n14654 & n14656;
  assign n10426 = x70 & x101;
  assign n10427 = n10425 & n10426;
  assign n10428 = n10425 | n10426;
  assign n10429 = ~n10427 & n10428;
  assign n14657 = n10266 & n10429;
  assign n14658 = (n10429 & n14578) | (n10429 & n14657) | (n14578 & n14657);
  assign n14659 = n10266 | n10429;
  assign n14660 = n14578 | n14659;
  assign n10432 = ~n14658 & n14660;
  assign n10433 = x69 & x102;
  assign n10434 = n10432 & n10433;
  assign n10435 = n10432 | n10433;
  assign n10436 = ~n10434 & n10435;
  assign n14661 = n10273 & n10436;
  assign n14662 = (n10436 & n14582) | (n10436 & n14661) | (n14582 & n14661);
  assign n14663 = n10273 | n10436;
  assign n14664 = n14582 | n14663;
  assign n10439 = ~n14662 & n14664;
  assign n10440 = x68 & x103;
  assign n10441 = n10439 & n10440;
  assign n10442 = n10439 | n10440;
  assign n10443 = ~n10441 & n10442;
  assign n14665 = n10280 & n10443;
  assign n14666 = (n10443 & n14586) | (n10443 & n14665) | (n14586 & n14665);
  assign n14667 = n10280 | n10443;
  assign n14668 = n14586 | n14667;
  assign n10446 = ~n14666 & n14668;
  assign n10447 = x67 & x104;
  assign n10448 = n10446 & n10447;
  assign n10449 = n10446 | n10447;
  assign n10450 = ~n10448 & n10449;
  assign n14669 = n10287 & n10450;
  assign n14670 = (n10450 & n14590) | (n10450 & n14669) | (n14590 & n14669);
  assign n14671 = n10287 | n10450;
  assign n14672 = n14590 | n14671;
  assign n10453 = ~n14670 & n14672;
  assign n10454 = x66 & x105;
  assign n10455 = n10453 & n10454;
  assign n10456 = n10453 | n10454;
  assign n10457 = ~n10455 & n10456;
  assign n14673 = n10294 & n10457;
  assign n14674 = (n10457 & n14595) | (n10457 & n14673) | (n14595 & n14673);
  assign n14675 = n10294 | n10457;
  assign n14676 = n14595 | n14675;
  assign n10460 = ~n14674 & n14676;
  assign n10461 = x65 & x106;
  assign n10462 = n10460 & n10461;
  assign n10463 = n10460 | n10461;
  assign n10464 = ~n10462 & n10463;
  assign n14609 = n10301 | n10303;
  assign n14677 = n10464 & n14609;
  assign n14678 = n10301 & n10464;
  assign n14679 = (n14519 & n14677) | (n14519 & n14678) | (n14677 & n14678);
  assign n14680 = n10464 | n14609;
  assign n14681 = n10301 | n10464;
  assign n14682 = (n14519 & n14680) | (n14519 & n14681) | (n14680 & n14681);
  assign n10467 = ~n14679 & n14682;
  assign n10468 = x64 & x107;
  assign n10469 = n10467 & n10468;
  assign n10470 = n10467 | n10468;
  assign n10471 = ~n10469 & n10470;
  assign n14607 = n10308 | n10310;
  assign n17222 = n10471 & n14607;
  assign n17223 = n10308 & n10471;
  assign n17224 = (n14517 & n17222) | (n14517 & n17223) | (n17222 & n17223);
  assign n17225 = n10471 | n14607;
  assign n17226 = n10308 | n10471;
  assign n17227 = (n14517 & n17225) | (n14517 & n17226) | (n17225 & n17226);
  assign n10474 = ~n17224 & n17227;
  assign n10475 = x63 & x108;
  assign n10476 = n10474 & n10475;
  assign n10477 = n10474 | n10475;
  assign n10478 = ~n10476 & n10477;
  assign n14605 = n10315 | n10317;
  assign n17228 = n10478 & n14605;
  assign n17229 = n10315 & n10478;
  assign n17230 = (n14515 & n17228) | (n14515 & n17229) | (n17228 & n17229);
  assign n17231 = n10478 | n14605;
  assign n17232 = n10315 | n10478;
  assign n17233 = (n14515 & n17231) | (n14515 & n17232) | (n17231 & n17232);
  assign n10481 = ~n17230 & n17233;
  assign n10482 = x62 & x109;
  assign n10483 = n10481 & n10482;
  assign n10484 = n10481 | n10482;
  assign n10485 = ~n10483 & n10484;
  assign n10486 = n14604 & n10485;
  assign n10487 = n14604 | n10485;
  assign n10488 = ~n10486 & n10487;
  assign n10489 = x61 & x110;
  assign n10490 = n10488 & n10489;
  assign n10491 = n10488 | n10489;
  assign n10492 = ~n10490 & n10491;
  assign n10493 = n14602 & n10492;
  assign n10494 = n14602 | n10492;
  assign n10495 = ~n10493 & n10494;
  assign n10496 = x60 & x111;
  assign n10497 = n10495 & n10496;
  assign n10498 = n10495 | n10496;
  assign n10499 = ~n10497 & n10498;
  assign n10500 = n14600 & n10499;
  assign n10501 = n14600 | n10499;
  assign n10502 = ~n10500 & n10501;
  assign n14683 = n10497 | n10499;
  assign n14684 = (n10497 & n14600) | (n10497 & n14683) | (n14600 & n14683);
  assign n14685 = n10490 | n10492;
  assign n14686 = (n10490 & n14602) | (n10490 & n14685) | (n14602 & n14685);
  assign n14606 = (n10315 & n14515) | (n10315 & n14605) | (n14515 & n14605);
  assign n14608 = (n10308 & n14517) | (n10308 & n14607) | (n14517 & n14607);
  assign n14699 = n10378 | n10380;
  assign n17236 = n10217 | n10378;
  assign n17237 = (n10378 & n10380) | (n10378 & n17236) | (n10380 & n17236);
  assign n17238 = (n14552 & n14699) | (n14552 & n17237) | (n14699 & n17237);
  assign n17239 = (n14551 & n14699) | (n14551 & n17237) | (n14699 & n17237);
  assign n17240 = (n17110 & n17238) | (n17110 & n17239) | (n17238 & n17239);
  assign n10523 = x79 & x93;
  assign n17858 = n10363 & n10523;
  assign n17983 = n17156 & n17858;
  assign n17859 = (n17162 & n17983) | (n17162 & n17858) | (n17983 & n17858);
  assign n17855 = n10523 & n17852;
  assign n17856 = (n17115 & n17859) | (n17115 & n17855) | (n17859 & n17855);
  assign n17242 = (n10366 & n10523) | (n10366 & n17856) | (n10523 & n17856);
  assign n17244 = n10523 & n17852;
  assign n17245 = (n17115 & n17859) | (n17115 & n17244) | (n17859 & n17244);
  assign n14705 = (n17209 & n17242) | (n17209 & n17245) | (n17242 & n17245);
  assign n17863 = n10363 | n10523;
  assign n17984 = (n10523 & n17156) | (n10523 & n17863) | (n17156 & n17863);
  assign n17864 = (n17162 & n17984) | (n17162 & n17863) | (n17984 & n17863);
  assign n17860 = n10523 | n17852;
  assign n17861 = (n17115 & n17864) | (n17115 & n17860) | (n17864 & n17860);
  assign n17247 = n10366 | n17861;
  assign n17249 = n10523 | n17852;
  assign n17250 = (n17115 & n17864) | (n17115 & n17249) | (n17864 & n17249);
  assign n14708 = (n17209 & n17247) | (n17209 & n17250) | (n17247 & n17250);
  assign n10526 = ~n14705 & n14708;
  assign n14709 = n10371 & n10526;
  assign n17251 = (n10526 & n14626) | (n10526 & n14709) | (n14626 & n14709);
  assign n17252 = (n10526 & n14625) | (n10526 & n14709) | (n14625 & n14709);
  assign n17253 = (n17150 & n17251) | (n17150 & n17252) | (n17251 & n17252);
  assign n14711 = n10371 | n10526;
  assign n17254 = n14626 | n14711;
  assign n17255 = n14625 | n14711;
  assign n17256 = (n17150 & n17254) | (n17150 & n17255) | (n17254 & n17255);
  assign n10529 = ~n17253 & n17256;
  assign n10530 = x78 & x94;
  assign n10531 = n10529 & n10530;
  assign n10532 = n10529 | n10530;
  assign n10533 = ~n10531 & n10532;
  assign n10534 = n17240 & n10533;
  assign n10535 = n17240 | n10533;
  assign n10536 = ~n10534 & n10535;
  assign n10537 = x77 & x95;
  assign n10538 = n10536 & n10537;
  assign n10539 = n10536 | n10537;
  assign n10540 = ~n10538 & n10539;
  assign n14696 = n10385 | n10387;
  assign n14713 = n10540 & n14696;
  assign n14714 = n10385 & n10540;
  assign n14715 = (n17204 & n14713) | (n17204 & n14714) | (n14713 & n14714);
  assign n14716 = n10540 | n14696;
  assign n14717 = n10385 | n10540;
  assign n14718 = (n17204 & n14716) | (n17204 & n14717) | (n14716 & n14717);
  assign n10543 = ~n14715 & n14718;
  assign n10544 = x76 & x96;
  assign n10545 = n10543 & n10544;
  assign n10546 = n10543 | n10544;
  assign n10547 = ~n10545 & n10546;
  assign n14719 = n10392 & n10547;
  assign n17257 = (n10547 & n14636) | (n10547 & n14719) | (n14636 & n14719);
  assign n17258 = (n10547 & n14635) | (n10547 & n14719) | (n14635 & n14719);
  assign n17259 = (n14524 & n17257) | (n14524 & n17258) | (n17257 & n17258);
  assign n14721 = n10392 | n10547;
  assign n17260 = n14636 | n14721;
  assign n17261 = n14635 | n14721;
  assign n17262 = (n14524 & n17260) | (n14524 & n17261) | (n17260 & n17261);
  assign n10550 = ~n17259 & n17262;
  assign n10551 = x75 & x97;
  assign n10552 = n10550 & n10551;
  assign n10553 = n10550 | n10551;
  assign n10554 = ~n10552 & n10553;
  assign n14694 = n10399 | n10401;
  assign n17263 = n10554 & n14694;
  assign n17234 = n10238 | n10399;
  assign n17235 = (n10399 & n10401) | (n10399 & n17234) | (n10401 & n17234);
  assign n17264 = n10554 & n17235;
  assign n17265 = (n17184 & n17263) | (n17184 & n17264) | (n17263 & n17264);
  assign n17266 = n10554 | n14694;
  assign n17267 = n10554 | n17235;
  assign n17268 = (n17184 & n17266) | (n17184 & n17267) | (n17266 & n17267);
  assign n10557 = ~n17265 & n17268;
  assign n10558 = x74 & x98;
  assign n10559 = n10557 & n10558;
  assign n10560 = n10557 | n10558;
  assign n10561 = ~n10559 & n10560;
  assign n14723 = n10406 & n10561;
  assign n17269 = (n10561 & n14645) | (n10561 & n14723) | (n14645 & n14723);
  assign n17270 = (n10408 & n10561) | (n10408 & n14723) | (n10561 & n14723);
  assign n17271 = (n14566 & n17269) | (n14566 & n17270) | (n17269 & n17270);
  assign n14725 = n10406 | n10561;
  assign n17272 = n14645 | n14725;
  assign n17273 = n10408 | n14725;
  assign n17274 = (n14566 & n17272) | (n14566 & n17273) | (n17272 & n17273);
  assign n10564 = ~n17271 & n17274;
  assign n10565 = x73 & x99;
  assign n10566 = n10564 & n10565;
  assign n10567 = n10564 | n10565;
  assign n10568 = ~n10566 & n10567;
  assign n14727 = n10413 & n10568;
  assign n14728 = (n10568 & n14650) | (n10568 & n14727) | (n14650 & n14727);
  assign n14729 = n10413 | n10568;
  assign n14730 = n14650 | n14729;
  assign n10571 = ~n14728 & n14730;
  assign n10572 = x72 & x100;
  assign n10573 = n10571 & n10572;
  assign n10574 = n10571 | n10572;
  assign n10575 = ~n10573 & n10574;
  assign n14731 = n10420 & n10575;
  assign n14732 = (n10575 & n14654) | (n10575 & n14731) | (n14654 & n14731);
  assign n14733 = n10420 | n10575;
  assign n14734 = n14654 | n14733;
  assign n10578 = ~n14732 & n14734;
  assign n10579 = x71 & x101;
  assign n10580 = n10578 & n10579;
  assign n10581 = n10578 | n10579;
  assign n10582 = ~n10580 & n10581;
  assign n14735 = n10427 & n10582;
  assign n14736 = (n10582 & n14658) | (n10582 & n14735) | (n14658 & n14735);
  assign n14737 = n10427 | n10582;
  assign n14738 = n14658 | n14737;
  assign n10585 = ~n14736 & n14738;
  assign n10586 = x70 & x102;
  assign n10587 = n10585 & n10586;
  assign n10588 = n10585 | n10586;
  assign n10589 = ~n10587 & n10588;
  assign n14739 = n10434 & n10589;
  assign n14740 = (n10589 & n14662) | (n10589 & n14739) | (n14662 & n14739);
  assign n14741 = n10434 | n10589;
  assign n14742 = n14662 | n14741;
  assign n10592 = ~n14740 & n14742;
  assign n10593 = x69 & x103;
  assign n10594 = n10592 & n10593;
  assign n10595 = n10592 | n10593;
  assign n10596 = ~n10594 & n10595;
  assign n14743 = n10441 & n10596;
  assign n14744 = (n10596 & n14666) | (n10596 & n14743) | (n14666 & n14743);
  assign n14745 = n10441 | n10596;
  assign n14746 = n14666 | n14745;
  assign n10599 = ~n14744 & n14746;
  assign n10600 = x68 & x104;
  assign n10601 = n10599 & n10600;
  assign n10602 = n10599 | n10600;
  assign n10603 = ~n10601 & n10602;
  assign n14747 = n10448 & n10603;
  assign n14748 = (n10603 & n14670) | (n10603 & n14747) | (n14670 & n14747);
  assign n14749 = n10448 | n10603;
  assign n14750 = n14670 | n14749;
  assign n10606 = ~n14748 & n14750;
  assign n10607 = x67 & x105;
  assign n10608 = n10606 & n10607;
  assign n10609 = n10606 | n10607;
  assign n10610 = ~n10608 & n10609;
  assign n14751 = n10455 & n10610;
  assign n14752 = (n10610 & n14674) | (n10610 & n14751) | (n14674 & n14751);
  assign n14753 = n10455 | n10610;
  assign n14754 = n14674 | n14753;
  assign n10613 = ~n14752 & n14754;
  assign n10614 = x66 & x106;
  assign n10615 = n10613 & n10614;
  assign n10616 = n10613 | n10614;
  assign n10617 = ~n10615 & n10616;
  assign n14755 = n10462 & n10617;
  assign n14756 = (n10617 & n14679) | (n10617 & n14755) | (n14679 & n14755);
  assign n14757 = n10462 | n10617;
  assign n14758 = n14679 | n14757;
  assign n10620 = ~n14756 & n14758;
  assign n10621 = x65 & x107;
  assign n10622 = n10620 & n10621;
  assign n10623 = n10620 | n10621;
  assign n10624 = ~n10622 & n10623;
  assign n14691 = n10469 | n10471;
  assign n14759 = n10624 & n14691;
  assign n14760 = n10469 & n10624;
  assign n14761 = (n14608 & n14759) | (n14608 & n14760) | (n14759 & n14760);
  assign n14762 = n10624 | n14691;
  assign n14763 = n10469 | n10624;
  assign n14764 = (n14608 & n14762) | (n14608 & n14763) | (n14762 & n14763);
  assign n10627 = ~n14761 & n14764;
  assign n10628 = x64 & x108;
  assign n10629 = n10627 & n10628;
  assign n10630 = n10627 | n10628;
  assign n10631 = ~n10629 & n10630;
  assign n14689 = n10476 | n10478;
  assign n17275 = n10631 & n14689;
  assign n17276 = n10476 & n10631;
  assign n17277 = (n14606 & n17275) | (n14606 & n17276) | (n17275 & n17276);
  assign n17278 = n10631 | n14689;
  assign n17279 = n10476 | n10631;
  assign n17280 = (n14606 & n17278) | (n14606 & n17279) | (n17278 & n17279);
  assign n10634 = ~n17277 & n17280;
  assign n10635 = x63 & x109;
  assign n10636 = n10634 & n10635;
  assign n10637 = n10634 | n10635;
  assign n10638 = ~n10636 & n10637;
  assign n14687 = n10483 | n10485;
  assign n17281 = n10638 & n14687;
  assign n17282 = n10483 & n10638;
  assign n17283 = (n14604 & n17281) | (n14604 & n17282) | (n17281 & n17282);
  assign n17284 = n10638 | n14687;
  assign n17285 = n10483 | n10638;
  assign n17286 = (n14604 & n17284) | (n14604 & n17285) | (n17284 & n17285);
  assign n10641 = ~n17283 & n17286;
  assign n10642 = x62 & x110;
  assign n10643 = n10641 & n10642;
  assign n10644 = n10641 | n10642;
  assign n10645 = ~n10643 & n10644;
  assign n10646 = n14686 & n10645;
  assign n10647 = n14686 | n10645;
  assign n10648 = ~n10646 & n10647;
  assign n10649 = x61 & x111;
  assign n10650 = n10648 & n10649;
  assign n10651 = n10648 | n10649;
  assign n10652 = ~n10650 & n10651;
  assign n10653 = n14684 & n10652;
  assign n10654 = n14684 | n10652;
  assign n10655 = ~n10653 & n10654;
  assign n14765 = n10650 | n10652;
  assign n14766 = (n10650 & n14684) | (n10650 & n14765) | (n14684 & n14765);
  assign n14688 = (n10483 & n14604) | (n10483 & n14687) | (n14604 & n14687);
  assign n14690 = (n10476 & n14606) | (n10476 & n14689) | (n14606 & n14689);
  assign n14695 = (n17184 & n17235) | (n17184 & n14694) | (n17235 & n14694);
  assign n14776 = n10545 | n10547;
  assign n17287 = n10392 | n10545;
  assign n17288 = (n10545 & n10547) | (n10545 & n17287) | (n10547 & n17287);
  assign n17289 = (n14636 & n14776) | (n14636 & n17288) | (n14776 & n17288);
  assign n17290 = (n14635 & n14776) | (n14635 & n17288) | (n14776 & n17288);
  assign n17291 = (n14524 & n17289) | (n14524 & n17290) | (n17289 & n17290);
  assign n10675 = x79 & x94;
  assign n14781 = n10526 | n14705;
  assign n17292 = (n10371 & n14705) | (n10371 & n14781) | (n14705 & n14781);
  assign n14783 = n10675 & n17292;
  assign n18085 = n10675 & n17858;
  assign n18169 = n17156 & n18085;
  assign n18086 = (n17162 & n18169) | (n17162 & n18085) | (n18169 & n18085);
  assign n17986 = n10523 & n10675;
  assign n18087 = n17852 & n17986;
  assign n18083 = (n17115 & n18086) | (n17115 & n18087) | (n18086 & n18087);
  assign n17987 = (n10366 & n18083) | (n10366 & n17986) | (n18083 & n17986);
  assign n17990 = (n17115 & n18086) | (n17115 & n18087) | (n18086 & n18087);
  assign n17867 = (n17209 & n17987) | (n17209 & n17990) | (n17987 & n17990);
  assign n17294 = (n10526 & n10675) | (n10526 & n17867) | (n10675 & n17867);
  assign n17295 = (n14626 & n14783) | (n14626 & n17294) | (n14783 & n17294);
  assign n17296 = (n14625 & n14783) | (n14625 & n17294) | (n14783 & n17294);
  assign n17297 = (n17150 & n17295) | (n17150 & n17296) | (n17295 & n17296);
  assign n14786 = n10675 | n17292;
  assign n18091 = n10675 | n17858;
  assign n18170 = (n10675 & n17156) | (n10675 & n18091) | (n17156 & n18091);
  assign n18092 = (n17162 & n18170) | (n17162 & n18091) | (n18170 & n18091);
  assign n17992 = n10523 | n10675;
  assign n18093 = (n10675 & n17852) | (n10675 & n17992) | (n17852 & n17992);
  assign n18089 = (n17115 & n18092) | (n17115 & n18093) | (n18092 & n18093);
  assign n17993 = (n10366 & n18089) | (n10366 & n17992) | (n18089 & n17992);
  assign n17996 = (n17115 & n18092) | (n17115 & n18093) | (n18092 & n18093);
  assign n17870 = (n17209 & n17993) | (n17209 & n17996) | (n17993 & n17996);
  assign n17299 = n10526 | n17870;
  assign n17300 = (n14626 & n14786) | (n14626 & n17299) | (n14786 & n17299);
  assign n17301 = (n14625 & n14786) | (n14625 & n17299) | (n14786 & n17299);
  assign n17302 = (n17150 & n17300) | (n17150 & n17301) | (n17300 & n17301);
  assign n10678 = ~n17297 & n17302;
  assign n14790 = n10531 & n10678;
  assign n17303 = (n10533 & n10678) | (n10533 & n14790) | (n10678 & n14790);
  assign n14791 = (n17240 & n17303) | (n17240 & n14790) | (n17303 & n14790);
  assign n14793 = n10531 | n10678;
  assign n17304 = n10533 | n14793;
  assign n14794 = (n17240 & n17304) | (n17240 & n14793) | (n17304 & n14793);
  assign n10681 = ~n14791 & n14794;
  assign n10682 = x78 & x95;
  assign n10683 = n10681 & n10682;
  assign n10684 = n10681 | n10682;
  assign n10685 = ~n10683 & n10684;
  assign n14795 = n10538 & n10685;
  assign n17305 = (n10685 & n14714) | (n10685 & n14795) | (n14714 & n14795);
  assign n17306 = (n10685 & n14713) | (n10685 & n14795) | (n14713 & n14795);
  assign n17307 = (n17204 & n17305) | (n17204 & n17306) | (n17305 & n17306);
  assign n14797 = n10538 | n10685;
  assign n17308 = n14714 | n14797;
  assign n17309 = n14713 | n14797;
  assign n17310 = (n17204 & n17308) | (n17204 & n17309) | (n17308 & n17309);
  assign n10688 = ~n17307 & n17310;
  assign n10689 = x77 & x96;
  assign n10690 = n10688 & n10689;
  assign n10691 = n10688 | n10689;
  assign n10692 = ~n10690 & n10691;
  assign n10693 = n17291 & n10692;
  assign n10694 = n17291 | n10692;
  assign n10695 = ~n10693 & n10694;
  assign n10696 = x76 & x97;
  assign n10697 = n10695 & n10696;
  assign n10698 = n10695 | n10696;
  assign n10699 = ~n10697 & n10698;
  assign n14773 = n10552 | n10554;
  assign n14799 = n10699 & n14773;
  assign n14800 = n10552 & n10699;
  assign n14801 = (n14695 & n14799) | (n14695 & n14800) | (n14799 & n14800);
  assign n14802 = n10699 | n14773;
  assign n14803 = n10552 | n10699;
  assign n14804 = (n14695 & n14802) | (n14695 & n14803) | (n14802 & n14803);
  assign n10702 = ~n14801 & n14804;
  assign n10703 = x75 & x98;
  assign n10704 = n10702 & n10703;
  assign n10705 = n10702 | n10703;
  assign n10706 = ~n10704 & n10705;
  assign n14805 = n10559 & n10706;
  assign n14806 = (n10706 & n17271) | (n10706 & n14805) | (n17271 & n14805);
  assign n14807 = n10559 | n10706;
  assign n14808 = n17271 | n14807;
  assign n10709 = ~n14806 & n14808;
  assign n10710 = x74 & x99;
  assign n10711 = n10709 & n10710;
  assign n10712 = n10709 | n10710;
  assign n10713 = ~n10711 & n10712;
  assign n14809 = n10566 & n10713;
  assign n14810 = (n10713 & n14728) | (n10713 & n14809) | (n14728 & n14809);
  assign n14811 = n10566 | n10713;
  assign n14812 = n14728 | n14811;
  assign n10716 = ~n14810 & n14812;
  assign n10717 = x73 & x100;
  assign n10718 = n10716 & n10717;
  assign n10719 = n10716 | n10717;
  assign n10720 = ~n10718 & n10719;
  assign n14813 = n10573 & n10720;
  assign n14814 = (n10720 & n14732) | (n10720 & n14813) | (n14732 & n14813);
  assign n14815 = n10573 | n10720;
  assign n14816 = n14732 | n14815;
  assign n10723 = ~n14814 & n14816;
  assign n10724 = x72 & x101;
  assign n10725 = n10723 & n10724;
  assign n10726 = n10723 | n10724;
  assign n10727 = ~n10725 & n10726;
  assign n14817 = n10580 & n10727;
  assign n14818 = (n10727 & n14736) | (n10727 & n14817) | (n14736 & n14817);
  assign n14819 = n10580 | n10727;
  assign n14820 = n14736 | n14819;
  assign n10730 = ~n14818 & n14820;
  assign n10731 = x71 & x102;
  assign n10732 = n10730 & n10731;
  assign n10733 = n10730 | n10731;
  assign n10734 = ~n10732 & n10733;
  assign n14821 = n10587 & n10734;
  assign n14822 = (n10734 & n14740) | (n10734 & n14821) | (n14740 & n14821);
  assign n14823 = n10587 | n10734;
  assign n14824 = n14740 | n14823;
  assign n10737 = ~n14822 & n14824;
  assign n10738 = x70 & x103;
  assign n10739 = n10737 & n10738;
  assign n10740 = n10737 | n10738;
  assign n10741 = ~n10739 & n10740;
  assign n14825 = n10594 & n10741;
  assign n14826 = (n10741 & n14744) | (n10741 & n14825) | (n14744 & n14825);
  assign n14827 = n10594 | n10741;
  assign n14828 = n14744 | n14827;
  assign n10744 = ~n14826 & n14828;
  assign n10745 = x69 & x104;
  assign n10746 = n10744 & n10745;
  assign n10747 = n10744 | n10745;
  assign n10748 = ~n10746 & n10747;
  assign n14829 = n10601 & n10748;
  assign n14830 = (n10748 & n14748) | (n10748 & n14829) | (n14748 & n14829);
  assign n14831 = n10601 | n10748;
  assign n14832 = n14748 | n14831;
  assign n10751 = ~n14830 & n14832;
  assign n10752 = x68 & x105;
  assign n10753 = n10751 & n10752;
  assign n10754 = n10751 | n10752;
  assign n10755 = ~n10753 & n10754;
  assign n14833 = n10608 & n10755;
  assign n14834 = (n10755 & n14752) | (n10755 & n14833) | (n14752 & n14833);
  assign n14835 = n10608 | n10755;
  assign n14836 = n14752 | n14835;
  assign n10758 = ~n14834 & n14836;
  assign n10759 = x67 & x106;
  assign n10760 = n10758 & n10759;
  assign n10761 = n10758 | n10759;
  assign n10762 = ~n10760 & n10761;
  assign n14837 = n10615 & n10762;
  assign n14838 = (n10762 & n14756) | (n10762 & n14837) | (n14756 & n14837);
  assign n14839 = n10615 | n10762;
  assign n14840 = n14756 | n14839;
  assign n10765 = ~n14838 & n14840;
  assign n10766 = x66 & x107;
  assign n10767 = n10765 & n10766;
  assign n10768 = n10765 | n10766;
  assign n10769 = ~n10767 & n10768;
  assign n14841 = n10622 & n10769;
  assign n14842 = (n10769 & n14761) | (n10769 & n14841) | (n14761 & n14841);
  assign n14843 = n10622 | n10769;
  assign n14844 = n14761 | n14843;
  assign n10772 = ~n14842 & n14844;
  assign n10773 = x65 & x108;
  assign n10774 = n10772 & n10773;
  assign n10775 = n10772 | n10773;
  assign n10776 = ~n10774 & n10775;
  assign n14771 = n10629 | n10631;
  assign n14845 = n10776 & n14771;
  assign n14846 = n10629 & n10776;
  assign n14847 = (n14690 & n14845) | (n14690 & n14846) | (n14845 & n14846);
  assign n14848 = n10776 | n14771;
  assign n14849 = n10629 | n10776;
  assign n14850 = (n14690 & n14848) | (n14690 & n14849) | (n14848 & n14849);
  assign n10779 = ~n14847 & n14850;
  assign n10780 = x64 & x109;
  assign n10781 = n10779 & n10780;
  assign n10782 = n10779 | n10780;
  assign n10783 = ~n10781 & n10782;
  assign n14769 = n10636 | n10638;
  assign n17311 = n10783 & n14769;
  assign n17312 = n10636 & n10783;
  assign n17313 = (n14688 & n17311) | (n14688 & n17312) | (n17311 & n17312);
  assign n17314 = n10783 | n14769;
  assign n17315 = n10636 | n10783;
  assign n17316 = (n14688 & n17314) | (n14688 & n17315) | (n17314 & n17315);
  assign n10786 = ~n17313 & n17316;
  assign n10787 = x63 & x110;
  assign n10788 = n10786 & n10787;
  assign n10789 = n10786 | n10787;
  assign n10790 = ~n10788 & n10789;
  assign n14767 = n10643 | n10645;
  assign n17317 = n10790 & n14767;
  assign n17318 = n10643 & n10790;
  assign n17319 = (n14686 & n17317) | (n14686 & n17318) | (n17317 & n17318);
  assign n17320 = n10790 | n14767;
  assign n17321 = n10643 | n10790;
  assign n17322 = (n14686 & n17320) | (n14686 & n17321) | (n17320 & n17321);
  assign n10793 = ~n17319 & n17322;
  assign n10794 = x62 & x111;
  assign n10795 = n10793 & n10794;
  assign n10796 = n10793 | n10794;
  assign n10797 = ~n10795 & n10796;
  assign n10798 = n14766 & n10797;
  assign n10799 = n14766 | n10797;
  assign n10800 = ~n10798 & n10799;
  assign n14768 = (n10643 & n14686) | (n10643 & n14767) | (n14686 & n14767);
  assign n14770 = (n10636 & n14688) | (n10636 & n14769) | (n14688 & n14769);
  assign n14863 = n10683 | n10685;
  assign n17325 = n10538 | n10683;
  assign n17326 = (n10683 & n10685) | (n10683 & n17325) | (n10685 & n17325);
  assign n17327 = (n14714 & n14863) | (n14714 & n17326) | (n14863 & n17326);
  assign n17328 = (n14713 & n14863) | (n14713 & n17326) | (n14863 & n17326);
  assign n17329 = (n17204 & n17327) | (n17204 & n17328) | (n17327 & n17328);
  assign n10819 = x79 & x95;
  assign n14865 = n10819 & n17297;
  assign n17330 = (n10819 & n14865) | (n10819 & n17303) | (n14865 & n17303);
  assign n17871 = (n10678 & n10819) | (n10678 & n14865) | (n10819 & n14865);
  assign n17997 = n10819 & n17297;
  assign n17873 = (n10531 & n17871) | (n10531 & n17997) | (n17871 & n17997);
  assign n17332 = (n17240 & n17330) | (n17240 & n17873) | (n17330 & n17873);
  assign n14867 = n10819 | n17297;
  assign n17333 = n14867 | n17303;
  assign n17874 = n10678 | n14867;
  assign n17875 = (n10531 & n14867) | (n10531 & n17874) | (n14867 & n17874);
  assign n17335 = (n17240 & n17333) | (n17240 & n17875) | (n17333 & n17875);
  assign n10822 = ~n17332 & n17335;
  assign n10823 = n17329 & n10822;
  assign n10824 = n17329 | n10822;
  assign n10825 = ~n10823 & n10824;
  assign n10826 = x78 & x96;
  assign n10827 = n10825 & n10826;
  assign n10828 = n10825 | n10826;
  assign n10829 = ~n10827 & n10828;
  assign n14860 = n10690 | n10692;
  assign n14869 = n10829 & n14860;
  assign n14870 = n10690 & n10829;
  assign n14871 = (n17291 & n14869) | (n17291 & n14870) | (n14869 & n14870);
  assign n14872 = n10829 | n14860;
  assign n14873 = n10690 | n10829;
  assign n14874 = (n17291 & n14872) | (n17291 & n14873) | (n14872 & n14873);
  assign n10832 = ~n14871 & n14874;
  assign n10833 = x77 & x97;
  assign n10834 = n10832 & n10833;
  assign n10835 = n10832 | n10833;
  assign n10836 = ~n10834 & n10835;
  assign n14875 = n10697 & n10836;
  assign n17336 = (n10836 & n14800) | (n10836 & n14875) | (n14800 & n14875);
  assign n17337 = (n10836 & n14799) | (n10836 & n14875) | (n14799 & n14875);
  assign n17338 = (n14695 & n17336) | (n14695 & n17337) | (n17336 & n17337);
  assign n14877 = n10697 | n10836;
  assign n17339 = n14800 | n14877;
  assign n17340 = n14799 | n14877;
  assign n17341 = (n14695 & n17339) | (n14695 & n17340) | (n17339 & n17340);
  assign n10839 = ~n17338 & n17341;
  assign n10840 = x76 & x98;
  assign n10841 = n10839 & n10840;
  assign n10842 = n10839 | n10840;
  assign n10843 = ~n10841 & n10842;
  assign n14858 = n10704 | n10706;
  assign n17342 = n10843 & n14858;
  assign n17323 = n10559 | n10704;
  assign n17324 = (n10704 & n10706) | (n10704 & n17323) | (n10706 & n17323);
  assign n17343 = n10843 & n17324;
  assign n17344 = (n17271 & n17342) | (n17271 & n17343) | (n17342 & n17343);
  assign n17345 = n10843 | n14858;
  assign n17346 = n10843 | n17324;
  assign n17347 = (n17271 & n17345) | (n17271 & n17346) | (n17345 & n17346);
  assign n10846 = ~n17344 & n17347;
  assign n10847 = x75 & x99;
  assign n10848 = n10846 & n10847;
  assign n10849 = n10846 | n10847;
  assign n10850 = ~n10848 & n10849;
  assign n14879 = n10711 & n10850;
  assign n17348 = (n10850 & n14809) | (n10850 & n14879) | (n14809 & n14879);
  assign n17349 = (n10713 & n10850) | (n10713 & n14879) | (n10850 & n14879);
  assign n17350 = (n14728 & n17348) | (n14728 & n17349) | (n17348 & n17349);
  assign n14881 = n10711 | n10850;
  assign n17351 = n14809 | n14881;
  assign n17352 = n10713 | n14881;
  assign n17353 = (n14728 & n17351) | (n14728 & n17352) | (n17351 & n17352);
  assign n10853 = ~n17350 & n17353;
  assign n10854 = x74 & x100;
  assign n10855 = n10853 & n10854;
  assign n10856 = n10853 | n10854;
  assign n10857 = ~n10855 & n10856;
  assign n14883 = n10718 & n10857;
  assign n14884 = (n10857 & n14814) | (n10857 & n14883) | (n14814 & n14883);
  assign n14885 = n10718 | n10857;
  assign n14886 = n14814 | n14885;
  assign n10860 = ~n14884 & n14886;
  assign n10861 = x73 & x101;
  assign n10862 = n10860 & n10861;
  assign n10863 = n10860 | n10861;
  assign n10864 = ~n10862 & n10863;
  assign n14887 = n10725 & n10864;
  assign n14888 = (n10864 & n14818) | (n10864 & n14887) | (n14818 & n14887);
  assign n14889 = n10725 | n10864;
  assign n14890 = n14818 | n14889;
  assign n10867 = ~n14888 & n14890;
  assign n10868 = x72 & x102;
  assign n10869 = n10867 & n10868;
  assign n10870 = n10867 | n10868;
  assign n10871 = ~n10869 & n10870;
  assign n14891 = n10732 & n10871;
  assign n14892 = (n10871 & n14822) | (n10871 & n14891) | (n14822 & n14891);
  assign n14893 = n10732 | n10871;
  assign n14894 = n14822 | n14893;
  assign n10874 = ~n14892 & n14894;
  assign n10875 = x71 & x103;
  assign n10876 = n10874 & n10875;
  assign n10877 = n10874 | n10875;
  assign n10878 = ~n10876 & n10877;
  assign n14895 = n10739 & n10878;
  assign n14896 = (n10878 & n14826) | (n10878 & n14895) | (n14826 & n14895);
  assign n14897 = n10739 | n10878;
  assign n14898 = n14826 | n14897;
  assign n10881 = ~n14896 & n14898;
  assign n10882 = x70 & x104;
  assign n10883 = n10881 & n10882;
  assign n10884 = n10881 | n10882;
  assign n10885 = ~n10883 & n10884;
  assign n14899 = n10746 & n10885;
  assign n14900 = (n10885 & n14830) | (n10885 & n14899) | (n14830 & n14899);
  assign n14901 = n10746 | n10885;
  assign n14902 = n14830 | n14901;
  assign n10888 = ~n14900 & n14902;
  assign n10889 = x69 & x105;
  assign n10890 = n10888 & n10889;
  assign n10891 = n10888 | n10889;
  assign n10892 = ~n10890 & n10891;
  assign n14903 = n10753 & n10892;
  assign n14904 = (n10892 & n14834) | (n10892 & n14903) | (n14834 & n14903);
  assign n14905 = n10753 | n10892;
  assign n14906 = n14834 | n14905;
  assign n10895 = ~n14904 & n14906;
  assign n10896 = x68 & x106;
  assign n10897 = n10895 & n10896;
  assign n10898 = n10895 | n10896;
  assign n10899 = ~n10897 & n10898;
  assign n14907 = n10760 & n10899;
  assign n14908 = (n10899 & n14838) | (n10899 & n14907) | (n14838 & n14907);
  assign n14909 = n10760 | n10899;
  assign n14910 = n14838 | n14909;
  assign n10902 = ~n14908 & n14910;
  assign n10903 = x67 & x107;
  assign n10904 = n10902 & n10903;
  assign n10905 = n10902 | n10903;
  assign n10906 = ~n10904 & n10905;
  assign n14911 = n10767 & n10906;
  assign n14912 = (n10906 & n14842) | (n10906 & n14911) | (n14842 & n14911);
  assign n14913 = n10767 | n10906;
  assign n14914 = n14842 | n14913;
  assign n10909 = ~n14912 & n14914;
  assign n10910 = x66 & x108;
  assign n10911 = n10909 & n10910;
  assign n10912 = n10909 | n10910;
  assign n10913 = ~n10911 & n10912;
  assign n14915 = n10774 & n10913;
  assign n14916 = (n10913 & n14847) | (n10913 & n14915) | (n14847 & n14915);
  assign n14917 = n10774 | n10913;
  assign n14918 = n14847 | n14917;
  assign n10916 = ~n14916 & n14918;
  assign n10917 = x65 & x109;
  assign n10918 = n10916 & n10917;
  assign n10919 = n10916 | n10917;
  assign n10920 = ~n10918 & n10919;
  assign n14855 = n10781 | n10783;
  assign n14919 = n10920 & n14855;
  assign n14920 = n10781 & n10920;
  assign n14921 = (n14770 & n14919) | (n14770 & n14920) | (n14919 & n14920);
  assign n14922 = n10920 | n14855;
  assign n14923 = n10781 | n10920;
  assign n14924 = (n14770 & n14922) | (n14770 & n14923) | (n14922 & n14923);
  assign n10923 = ~n14921 & n14924;
  assign n10924 = x64 & x110;
  assign n10925 = n10923 & n10924;
  assign n10926 = n10923 | n10924;
  assign n10927 = ~n10925 & n10926;
  assign n14853 = n10788 | n10790;
  assign n17354 = n10927 & n14853;
  assign n17355 = n10788 & n10927;
  assign n17356 = (n14768 & n17354) | (n14768 & n17355) | (n17354 & n17355);
  assign n17357 = n10927 | n14853;
  assign n17358 = n10788 | n10927;
  assign n17359 = (n14768 & n17357) | (n14768 & n17358) | (n17357 & n17358);
  assign n10930 = ~n17356 & n17359;
  assign n10931 = x63 & x111;
  assign n10932 = n10930 & n10931;
  assign n10933 = n10930 | n10931;
  assign n10934 = ~n10932 & n10933;
  assign n14851 = n10795 | n10797;
  assign n17360 = n10934 & n14851;
  assign n17361 = n10795 & n10934;
  assign n17362 = (n14766 & n17360) | (n14766 & n17361) | (n17360 & n17361);
  assign n17363 = n10934 | n14851;
  assign n17364 = n10795 | n10934;
  assign n17365 = (n14766 & n17363) | (n14766 & n17364) | (n17363 & n17364);
  assign n10937 = ~n17362 & n17365;
  assign n14852 = (n10795 & n14766) | (n10795 & n14851) | (n14766 & n14851);
  assign n14854 = (n10788 & n14768) | (n10788 & n14853) | (n14768 & n14853);
  assign n14859 = (n17271 & n17324) | (n17271 & n14858) | (n17324 & n14858);
  assign n14932 = n10834 | n10836;
  assign n17366 = n10697 | n10834;
  assign n17367 = (n10834 & n10836) | (n10834 & n17366) | (n10836 & n17366);
  assign n17368 = (n14800 & n14932) | (n14800 & n17367) | (n14932 & n17367);
  assign n17369 = (n14799 & n14932) | (n14799 & n17367) | (n14932 & n17367);
  assign n17370 = (n14695 & n17368) | (n14695 & n17369) | (n17368 & n17369);
  assign n10955 = x79 & x96;
  assign n17879 = n10819 & n10955;
  assign n17998 = n17297 & n17879;
  assign n17880 = (n17303 & n17998) | (n17303 & n17879) | (n17998 & n17879);
  assign n17876 = n10955 & n17873;
  assign n17877 = (n17240 & n17880) | (n17240 & n17876) | (n17880 & n17876);
  assign n17372 = (n10822 & n10955) | (n10822 & n17877) | (n10955 & n17877);
  assign n17374 = n10955 & n17873;
  assign n17375 = (n17240 & n17880) | (n17240 & n17374) | (n17880 & n17374);
  assign n14938 = (n17329 & n17372) | (n17329 & n17375) | (n17372 & n17375);
  assign n17884 = n10819 | n10955;
  assign n17999 = (n10955 & n17297) | (n10955 & n17884) | (n17297 & n17884);
  assign n17885 = (n17303 & n17999) | (n17303 & n17884) | (n17999 & n17884);
  assign n17881 = n10955 | n17873;
  assign n17882 = (n17240 & n17885) | (n17240 & n17881) | (n17885 & n17881);
  assign n17377 = n10822 | n17882;
  assign n17379 = n10955 | n17873;
  assign n17380 = (n17240 & n17885) | (n17240 & n17379) | (n17885 & n17379);
  assign n14941 = (n17329 & n17377) | (n17329 & n17380) | (n17377 & n17380);
  assign n10958 = ~n14938 & n14941;
  assign n14942 = n10827 & n10958;
  assign n17381 = (n10958 & n14870) | (n10958 & n14942) | (n14870 & n14942);
  assign n17382 = (n10958 & n14869) | (n10958 & n14942) | (n14869 & n14942);
  assign n17383 = (n17291 & n17381) | (n17291 & n17382) | (n17381 & n17382);
  assign n14944 = n10827 | n10958;
  assign n17384 = n14870 | n14944;
  assign n17385 = n14869 | n14944;
  assign n17386 = (n17291 & n17384) | (n17291 & n17385) | (n17384 & n17385);
  assign n10961 = ~n17383 & n17386;
  assign n10962 = x78 & x97;
  assign n10963 = n10961 & n10962;
  assign n10964 = n10961 | n10962;
  assign n10965 = ~n10963 & n10964;
  assign n10966 = n17370 & n10965;
  assign n10967 = n17370 | n10965;
  assign n10968 = ~n10966 & n10967;
  assign n10969 = x77 & x98;
  assign n10970 = n10968 & n10969;
  assign n10971 = n10968 | n10969;
  assign n10972 = ~n10970 & n10971;
  assign n14929 = n10841 | n10843;
  assign n14946 = n10972 & n14929;
  assign n14947 = n10841 & n10972;
  assign n14948 = (n14859 & n14946) | (n14859 & n14947) | (n14946 & n14947);
  assign n14949 = n10972 | n14929;
  assign n14950 = n10841 | n10972;
  assign n14951 = (n14859 & n14949) | (n14859 & n14950) | (n14949 & n14950);
  assign n10975 = ~n14948 & n14951;
  assign n10976 = x76 & x99;
  assign n10977 = n10975 & n10976;
  assign n10978 = n10975 | n10976;
  assign n10979 = ~n10977 & n10978;
  assign n14952 = n10848 & n10979;
  assign n14953 = (n10979 & n17350) | (n10979 & n14952) | (n17350 & n14952);
  assign n14954 = n10848 | n10979;
  assign n14955 = n17350 | n14954;
  assign n10982 = ~n14953 & n14955;
  assign n10983 = x75 & x100;
  assign n10984 = n10982 & n10983;
  assign n10985 = n10982 | n10983;
  assign n10986 = ~n10984 & n10985;
  assign n14956 = n10855 & n10986;
  assign n14957 = (n10986 & n14884) | (n10986 & n14956) | (n14884 & n14956);
  assign n14958 = n10855 | n10986;
  assign n14959 = n14884 | n14958;
  assign n10989 = ~n14957 & n14959;
  assign n10990 = x74 & x101;
  assign n10991 = n10989 & n10990;
  assign n10992 = n10989 | n10990;
  assign n10993 = ~n10991 & n10992;
  assign n14960 = n10862 & n10993;
  assign n14961 = (n10993 & n14888) | (n10993 & n14960) | (n14888 & n14960);
  assign n14962 = n10862 | n10993;
  assign n14963 = n14888 | n14962;
  assign n10996 = ~n14961 & n14963;
  assign n10997 = x73 & x102;
  assign n10998 = n10996 & n10997;
  assign n10999 = n10996 | n10997;
  assign n11000 = ~n10998 & n10999;
  assign n14964 = n10869 & n11000;
  assign n14965 = (n11000 & n14892) | (n11000 & n14964) | (n14892 & n14964);
  assign n14966 = n10869 | n11000;
  assign n14967 = n14892 | n14966;
  assign n11003 = ~n14965 & n14967;
  assign n11004 = x72 & x103;
  assign n11005 = n11003 & n11004;
  assign n11006 = n11003 | n11004;
  assign n11007 = ~n11005 & n11006;
  assign n14968 = n10876 & n11007;
  assign n14969 = (n11007 & n14896) | (n11007 & n14968) | (n14896 & n14968);
  assign n14970 = n10876 | n11007;
  assign n14971 = n14896 | n14970;
  assign n11010 = ~n14969 & n14971;
  assign n11011 = x71 & x104;
  assign n11012 = n11010 & n11011;
  assign n11013 = n11010 | n11011;
  assign n11014 = ~n11012 & n11013;
  assign n14972 = n10883 & n11014;
  assign n14973 = (n11014 & n14900) | (n11014 & n14972) | (n14900 & n14972);
  assign n14974 = n10883 | n11014;
  assign n14975 = n14900 | n14974;
  assign n11017 = ~n14973 & n14975;
  assign n11018 = x70 & x105;
  assign n11019 = n11017 & n11018;
  assign n11020 = n11017 | n11018;
  assign n11021 = ~n11019 & n11020;
  assign n14976 = n10890 & n11021;
  assign n14977 = (n11021 & n14904) | (n11021 & n14976) | (n14904 & n14976);
  assign n14978 = n10890 | n11021;
  assign n14979 = n14904 | n14978;
  assign n11024 = ~n14977 & n14979;
  assign n11025 = x69 & x106;
  assign n11026 = n11024 & n11025;
  assign n11027 = n11024 | n11025;
  assign n11028 = ~n11026 & n11027;
  assign n14980 = n10897 & n11028;
  assign n14981 = (n11028 & n14908) | (n11028 & n14980) | (n14908 & n14980);
  assign n14982 = n10897 | n11028;
  assign n14983 = n14908 | n14982;
  assign n11031 = ~n14981 & n14983;
  assign n11032 = x68 & x107;
  assign n11033 = n11031 & n11032;
  assign n11034 = n11031 | n11032;
  assign n11035 = ~n11033 & n11034;
  assign n14984 = n10904 & n11035;
  assign n14985 = (n11035 & n14912) | (n11035 & n14984) | (n14912 & n14984);
  assign n14986 = n10904 | n11035;
  assign n14987 = n14912 | n14986;
  assign n11038 = ~n14985 & n14987;
  assign n11039 = x67 & x108;
  assign n11040 = n11038 & n11039;
  assign n11041 = n11038 | n11039;
  assign n11042 = ~n11040 & n11041;
  assign n14988 = n10911 & n11042;
  assign n14989 = (n11042 & n14916) | (n11042 & n14988) | (n14916 & n14988);
  assign n14990 = n10911 | n11042;
  assign n14991 = n14916 | n14990;
  assign n11045 = ~n14989 & n14991;
  assign n11046 = x66 & x109;
  assign n11047 = n11045 & n11046;
  assign n11048 = n11045 | n11046;
  assign n11049 = ~n11047 & n11048;
  assign n14992 = n10918 & n11049;
  assign n14993 = (n11049 & n14921) | (n11049 & n14992) | (n14921 & n14992);
  assign n14994 = n10918 | n11049;
  assign n14995 = n14921 | n14994;
  assign n11052 = ~n14993 & n14995;
  assign n11053 = x65 & x110;
  assign n11054 = n11052 & n11053;
  assign n11055 = n11052 | n11053;
  assign n11056 = ~n11054 & n11055;
  assign n14927 = n10925 | n10927;
  assign n14996 = n11056 & n14927;
  assign n14997 = n10925 & n11056;
  assign n14998 = (n14854 & n14996) | (n14854 & n14997) | (n14996 & n14997);
  assign n14999 = n11056 | n14927;
  assign n15000 = n10925 | n11056;
  assign n15001 = (n14854 & n14999) | (n14854 & n15000) | (n14999 & n15000);
  assign n11059 = ~n14998 & n15001;
  assign n11060 = x64 & x111;
  assign n11061 = n11059 & n11060;
  assign n11062 = n11059 | n11060;
  assign n11063 = ~n11061 & n11062;
  assign n14925 = n10932 | n10934;
  assign n17387 = n11063 & n14925;
  assign n17388 = n10932 & n11063;
  assign n17389 = (n14852 & n17387) | (n14852 & n17388) | (n17387 & n17388);
  assign n17390 = n11063 | n14925;
  assign n17391 = n10932 | n11063;
  assign n17392 = (n14852 & n17390) | (n14852 & n17391) | (n17390 & n17391);
  assign n11066 = ~n17389 & n17392;
  assign n14926 = (n10932 & n14852) | (n10932 & n14925) | (n14852 & n14925);
  assign n11083 = x79 & x97;
  assign n15010 = n10958 | n14938;
  assign n17395 = (n10827 & n14938) | (n10827 & n15010) | (n14938 & n15010);
  assign n15012 = n11083 & n17395;
  assign n18097 = n11083 & n17879;
  assign n18171 = n17297 & n18097;
  assign n18098 = (n17303 & n18171) | (n17303 & n18097) | (n18171 & n18097);
  assign n18001 = n10955 & n11083;
  assign n18099 = n17873 & n18001;
  assign n18095 = (n17240 & n18098) | (n17240 & n18099) | (n18098 & n18099);
  assign n18002 = (n10822 & n18095) | (n10822 & n18001) | (n18095 & n18001);
  assign n18005 = (n17240 & n18098) | (n17240 & n18099) | (n18098 & n18099);
  assign n17888 = (n17329 & n18002) | (n17329 & n18005) | (n18002 & n18005);
  assign n17397 = (n10958 & n11083) | (n10958 & n17888) | (n11083 & n17888);
  assign n17398 = (n14870 & n15012) | (n14870 & n17397) | (n15012 & n17397);
  assign n17399 = (n14869 & n15012) | (n14869 & n17397) | (n15012 & n17397);
  assign n17400 = (n17291 & n17398) | (n17291 & n17399) | (n17398 & n17399);
  assign n15015 = n11083 | n17395;
  assign n18103 = n11083 | n17879;
  assign n18172 = (n11083 & n17297) | (n11083 & n18103) | (n17297 & n18103);
  assign n18104 = (n17303 & n18172) | (n17303 & n18103) | (n18172 & n18103);
  assign n18007 = n10955 | n11083;
  assign n18105 = (n11083 & n17873) | (n11083 & n18007) | (n17873 & n18007);
  assign n18101 = (n17240 & n18104) | (n17240 & n18105) | (n18104 & n18105);
  assign n18008 = (n10822 & n18101) | (n10822 & n18007) | (n18101 & n18007);
  assign n18011 = (n17240 & n18104) | (n17240 & n18105) | (n18104 & n18105);
  assign n17891 = (n17329 & n18008) | (n17329 & n18011) | (n18008 & n18011);
  assign n17402 = n10958 | n17891;
  assign n17403 = (n14870 & n15015) | (n14870 & n17402) | (n15015 & n17402);
  assign n17404 = (n14869 & n15015) | (n14869 & n17402) | (n15015 & n17402);
  assign n17405 = (n17291 & n17403) | (n17291 & n17404) | (n17403 & n17404);
  assign n11086 = ~n17400 & n17405;
  assign n15019 = n10963 & n11086;
  assign n17406 = (n10965 & n11086) | (n10965 & n15019) | (n11086 & n15019);
  assign n15020 = (n17370 & n17406) | (n17370 & n15019) | (n17406 & n15019);
  assign n15022 = n10963 | n11086;
  assign n17407 = n10965 | n15022;
  assign n15023 = (n17370 & n17407) | (n17370 & n15022) | (n17407 & n15022);
  assign n11089 = ~n15020 & n15023;
  assign n11090 = x78 & x98;
  assign n11091 = n11089 & n11090;
  assign n11092 = n11089 | n11090;
  assign n11093 = ~n11091 & n11092;
  assign n15024 = n10970 & n11093;
  assign n17408 = (n11093 & n14947) | (n11093 & n15024) | (n14947 & n15024);
  assign n17409 = (n11093 & n14946) | (n11093 & n15024) | (n14946 & n15024);
  assign n17410 = (n14859 & n17408) | (n14859 & n17409) | (n17408 & n17409);
  assign n15026 = n10970 | n11093;
  assign n17411 = n14947 | n15026;
  assign n17412 = n14946 | n15026;
  assign n17413 = (n14859 & n17411) | (n14859 & n17412) | (n17411 & n17412);
  assign n11096 = ~n17410 & n17413;
  assign n11097 = x77 & x99;
  assign n11098 = n11096 & n11097;
  assign n11099 = n11096 | n11097;
  assign n11100 = ~n11098 & n11099;
  assign n15005 = n10977 | n10979;
  assign n17414 = n11100 & n15005;
  assign n17393 = n10848 | n10977;
  assign n17394 = (n10977 & n10979) | (n10977 & n17393) | (n10979 & n17393);
  assign n17415 = n11100 & n17394;
  assign n17416 = (n17350 & n17414) | (n17350 & n17415) | (n17414 & n17415);
  assign n17417 = n11100 | n15005;
  assign n17418 = n11100 | n17394;
  assign n17419 = (n17350 & n17417) | (n17350 & n17418) | (n17417 & n17418);
  assign n11103 = ~n17416 & n17419;
  assign n11104 = x76 & x100;
  assign n11105 = n11103 & n11104;
  assign n11106 = n11103 | n11104;
  assign n11107 = ~n11105 & n11106;
  assign n15028 = n10984 & n11107;
  assign n17420 = (n11107 & n14956) | (n11107 & n15028) | (n14956 & n15028);
  assign n17421 = (n10986 & n11107) | (n10986 & n15028) | (n11107 & n15028);
  assign n17422 = (n14884 & n17420) | (n14884 & n17421) | (n17420 & n17421);
  assign n15030 = n10984 | n11107;
  assign n17423 = n14956 | n15030;
  assign n17424 = n10986 | n15030;
  assign n17425 = (n14884 & n17423) | (n14884 & n17424) | (n17423 & n17424);
  assign n11110 = ~n17422 & n17425;
  assign n11111 = x75 & x101;
  assign n11112 = n11110 & n11111;
  assign n11113 = n11110 | n11111;
  assign n11114 = ~n11112 & n11113;
  assign n15032 = n10991 & n11114;
  assign n15033 = (n11114 & n14961) | (n11114 & n15032) | (n14961 & n15032);
  assign n15034 = n10991 | n11114;
  assign n15035 = n14961 | n15034;
  assign n11117 = ~n15033 & n15035;
  assign n11118 = x74 & x102;
  assign n11119 = n11117 & n11118;
  assign n11120 = n11117 | n11118;
  assign n11121 = ~n11119 & n11120;
  assign n15036 = n10998 & n11121;
  assign n15037 = (n11121 & n14965) | (n11121 & n15036) | (n14965 & n15036);
  assign n15038 = n10998 | n11121;
  assign n15039 = n14965 | n15038;
  assign n11124 = ~n15037 & n15039;
  assign n11125 = x73 & x103;
  assign n11126 = n11124 & n11125;
  assign n11127 = n11124 | n11125;
  assign n11128 = ~n11126 & n11127;
  assign n15040 = n11005 & n11128;
  assign n15041 = (n11128 & n14969) | (n11128 & n15040) | (n14969 & n15040);
  assign n15042 = n11005 | n11128;
  assign n15043 = n14969 | n15042;
  assign n11131 = ~n15041 & n15043;
  assign n11132 = x72 & x104;
  assign n11133 = n11131 & n11132;
  assign n11134 = n11131 | n11132;
  assign n11135 = ~n11133 & n11134;
  assign n15044 = n11012 & n11135;
  assign n15045 = (n11135 & n14973) | (n11135 & n15044) | (n14973 & n15044);
  assign n15046 = n11012 | n11135;
  assign n15047 = n14973 | n15046;
  assign n11138 = ~n15045 & n15047;
  assign n11139 = x71 & x105;
  assign n11140 = n11138 & n11139;
  assign n11141 = n11138 | n11139;
  assign n11142 = ~n11140 & n11141;
  assign n15048 = n11019 & n11142;
  assign n15049 = (n11142 & n14977) | (n11142 & n15048) | (n14977 & n15048);
  assign n15050 = n11019 | n11142;
  assign n15051 = n14977 | n15050;
  assign n11145 = ~n15049 & n15051;
  assign n11146 = x70 & x106;
  assign n11147 = n11145 & n11146;
  assign n11148 = n11145 | n11146;
  assign n11149 = ~n11147 & n11148;
  assign n15052 = n11026 & n11149;
  assign n15053 = (n11149 & n14981) | (n11149 & n15052) | (n14981 & n15052);
  assign n15054 = n11026 | n11149;
  assign n15055 = n14981 | n15054;
  assign n11152 = ~n15053 & n15055;
  assign n11153 = x69 & x107;
  assign n11154 = n11152 & n11153;
  assign n11155 = n11152 | n11153;
  assign n11156 = ~n11154 & n11155;
  assign n15056 = n11033 & n11156;
  assign n15057 = (n11156 & n14985) | (n11156 & n15056) | (n14985 & n15056);
  assign n15058 = n11033 | n11156;
  assign n15059 = n14985 | n15058;
  assign n11159 = ~n15057 & n15059;
  assign n11160 = x68 & x108;
  assign n11161 = n11159 & n11160;
  assign n11162 = n11159 | n11160;
  assign n11163 = ~n11161 & n11162;
  assign n15060 = n11040 & n11163;
  assign n15061 = (n11163 & n14989) | (n11163 & n15060) | (n14989 & n15060);
  assign n15062 = n11040 | n11163;
  assign n15063 = n14989 | n15062;
  assign n11166 = ~n15061 & n15063;
  assign n11167 = x67 & x109;
  assign n11168 = n11166 & n11167;
  assign n11169 = n11166 | n11167;
  assign n11170 = ~n11168 & n11169;
  assign n15064 = n11047 & n11170;
  assign n15065 = (n11170 & n14993) | (n11170 & n15064) | (n14993 & n15064);
  assign n15066 = n11047 | n11170;
  assign n15067 = n14993 | n15066;
  assign n11173 = ~n15065 & n15067;
  assign n11174 = x66 & x110;
  assign n11175 = n11173 & n11174;
  assign n11176 = n11173 | n11174;
  assign n11177 = ~n11175 & n11176;
  assign n15068 = n11054 & n11177;
  assign n15069 = (n11177 & n14998) | (n11177 & n15068) | (n14998 & n15068);
  assign n15070 = n11054 | n11177;
  assign n15071 = n14998 | n15070;
  assign n11180 = ~n15069 & n15071;
  assign n11181 = x65 & x111;
  assign n11182 = n11180 & n11181;
  assign n11183 = n11180 | n11181;
  assign n11184 = ~n11182 & n11183;
  assign n15002 = n11061 | n11063;
  assign n15072 = n11184 & n15002;
  assign n15073 = n11061 & n11184;
  assign n15074 = (n14926 & n15072) | (n14926 & n15073) | (n15072 & n15073);
  assign n15075 = n11184 | n15002;
  assign n15076 = n11061 | n11184;
  assign n15077 = (n14926 & n15075) | (n14926 & n15076) | (n15075 & n15076);
  assign n11187 = ~n15074 & n15077;
  assign n15006 = (n17350 & n17394) | (n17350 & n15005) | (n17394 & n15005);
  assign n15081 = n11091 | n11093;
  assign n17426 = n10970 | n11091;
  assign n17427 = (n11091 & n11093) | (n11091 & n17426) | (n11093 & n17426);
  assign n17428 = (n14947 & n15081) | (n14947 & n17427) | (n15081 & n17427);
  assign n17429 = (n14946 & n15081) | (n14946 & n17427) | (n15081 & n17427);
  assign n17430 = (n14859 & n17428) | (n14859 & n17429) | (n17428 & n17429);
  assign n11203 = x79 & x98;
  assign n15083 = n11203 & n17400;
  assign n17431 = (n11203 & n15083) | (n11203 & n17406) | (n15083 & n17406);
  assign n17892 = (n11086 & n11203) | (n11086 & n15083) | (n11203 & n15083);
  assign n18012 = n11203 & n17400;
  assign n17894 = (n10963 & n17892) | (n10963 & n18012) | (n17892 & n18012);
  assign n17433 = (n17370 & n17431) | (n17370 & n17894) | (n17431 & n17894);
  assign n15085 = n11203 | n17400;
  assign n17434 = n15085 | n17406;
  assign n17895 = n11086 | n15085;
  assign n17896 = (n10963 & n15085) | (n10963 & n17895) | (n15085 & n17895);
  assign n17436 = (n17370 & n17434) | (n17370 & n17896) | (n17434 & n17896);
  assign n11206 = ~n17433 & n17436;
  assign n11207 = n17430 & n11206;
  assign n11208 = n17430 | n11206;
  assign n11209 = ~n11207 & n11208;
  assign n11210 = x78 & x99;
  assign n11211 = n11209 & n11210;
  assign n11212 = n11209 | n11210;
  assign n11213 = ~n11211 & n11212;
  assign n15078 = n11098 | n11100;
  assign n15087 = n11213 & n15078;
  assign n15088 = n11098 & n11213;
  assign n15089 = (n15006 & n15087) | (n15006 & n15088) | (n15087 & n15088);
  assign n15090 = n11213 | n15078;
  assign n15091 = n11098 | n11213;
  assign n15092 = (n15006 & n15090) | (n15006 & n15091) | (n15090 & n15091);
  assign n11216 = ~n15089 & n15092;
  assign n11217 = x77 & x100;
  assign n11218 = n11216 & n11217;
  assign n11219 = n11216 | n11217;
  assign n11220 = ~n11218 & n11219;
  assign n15093 = n11105 & n11220;
  assign n15094 = (n11220 & n17422) | (n11220 & n15093) | (n17422 & n15093);
  assign n15095 = n11105 | n11220;
  assign n15096 = n17422 | n15095;
  assign n11223 = ~n15094 & n15096;
  assign n11224 = x76 & x101;
  assign n11225 = n11223 & n11224;
  assign n11226 = n11223 | n11224;
  assign n11227 = ~n11225 & n11226;
  assign n15097 = n11112 & n11227;
  assign n15098 = (n11227 & n15033) | (n11227 & n15097) | (n15033 & n15097);
  assign n15099 = n11112 | n11227;
  assign n15100 = n15033 | n15099;
  assign n11230 = ~n15098 & n15100;
  assign n11231 = x75 & x102;
  assign n11232 = n11230 & n11231;
  assign n11233 = n11230 | n11231;
  assign n11234 = ~n11232 & n11233;
  assign n15101 = n11119 & n11234;
  assign n15102 = (n11234 & n15037) | (n11234 & n15101) | (n15037 & n15101);
  assign n15103 = n11119 | n11234;
  assign n15104 = n15037 | n15103;
  assign n11237 = ~n15102 & n15104;
  assign n11238 = x74 & x103;
  assign n11239 = n11237 & n11238;
  assign n11240 = n11237 | n11238;
  assign n11241 = ~n11239 & n11240;
  assign n15105 = n11126 & n11241;
  assign n15106 = (n11241 & n15041) | (n11241 & n15105) | (n15041 & n15105);
  assign n15107 = n11126 | n11241;
  assign n15108 = n15041 | n15107;
  assign n11244 = ~n15106 & n15108;
  assign n11245 = x73 & x104;
  assign n11246 = n11244 & n11245;
  assign n11247 = n11244 | n11245;
  assign n11248 = ~n11246 & n11247;
  assign n15109 = n11133 & n11248;
  assign n15110 = (n11248 & n15045) | (n11248 & n15109) | (n15045 & n15109);
  assign n15111 = n11133 | n11248;
  assign n15112 = n15045 | n15111;
  assign n11251 = ~n15110 & n15112;
  assign n11252 = x72 & x105;
  assign n11253 = n11251 & n11252;
  assign n11254 = n11251 | n11252;
  assign n11255 = ~n11253 & n11254;
  assign n15113 = n11140 & n11255;
  assign n15114 = (n11255 & n15049) | (n11255 & n15113) | (n15049 & n15113);
  assign n15115 = n11140 | n11255;
  assign n15116 = n15049 | n15115;
  assign n11258 = ~n15114 & n15116;
  assign n11259 = x71 & x106;
  assign n11260 = n11258 & n11259;
  assign n11261 = n11258 | n11259;
  assign n11262 = ~n11260 & n11261;
  assign n15117 = n11147 & n11262;
  assign n15118 = (n11262 & n15053) | (n11262 & n15117) | (n15053 & n15117);
  assign n15119 = n11147 | n11262;
  assign n15120 = n15053 | n15119;
  assign n11265 = ~n15118 & n15120;
  assign n11266 = x70 & x107;
  assign n11267 = n11265 & n11266;
  assign n11268 = n11265 | n11266;
  assign n11269 = ~n11267 & n11268;
  assign n15121 = n11154 & n11269;
  assign n15122 = (n11269 & n15057) | (n11269 & n15121) | (n15057 & n15121);
  assign n15123 = n11154 | n11269;
  assign n15124 = n15057 | n15123;
  assign n11272 = ~n15122 & n15124;
  assign n11273 = x69 & x108;
  assign n11274 = n11272 & n11273;
  assign n11275 = n11272 | n11273;
  assign n11276 = ~n11274 & n11275;
  assign n15125 = n11161 & n11276;
  assign n15126 = (n11276 & n15061) | (n11276 & n15125) | (n15061 & n15125);
  assign n15127 = n11161 | n11276;
  assign n15128 = n15061 | n15127;
  assign n11279 = ~n15126 & n15128;
  assign n11280 = x68 & x109;
  assign n11281 = n11279 & n11280;
  assign n11282 = n11279 | n11280;
  assign n11283 = ~n11281 & n11282;
  assign n15129 = n11168 & n11283;
  assign n15130 = (n11283 & n15065) | (n11283 & n15129) | (n15065 & n15129);
  assign n15131 = n11168 | n11283;
  assign n15132 = n15065 | n15131;
  assign n11286 = ~n15130 & n15132;
  assign n11287 = x67 & x110;
  assign n11288 = n11286 & n11287;
  assign n11289 = n11286 | n11287;
  assign n11290 = ~n11288 & n11289;
  assign n15133 = n11175 & n11290;
  assign n15134 = (n11290 & n15069) | (n11290 & n15133) | (n15069 & n15133);
  assign n15135 = n11175 | n11290;
  assign n15136 = n15069 | n15135;
  assign n11293 = ~n15134 & n15136;
  assign n11294 = x66 & x111;
  assign n11295 = n11293 & n11294;
  assign n11296 = n11293 | n11294;
  assign n11297 = ~n11295 & n11296;
  assign n15137 = n11182 & n11297;
  assign n15138 = (n11297 & n15074) | (n11297 & n15137) | (n15074 & n15137);
  assign n15139 = n11182 | n11297;
  assign n15140 = n15074 | n15139;
  assign n11300 = ~n15138 & n15140;
  assign n11315 = x79 & x99;
  assign n17900 = n11203 & n11315;
  assign n18013 = n17400 & n17900;
  assign n17901 = (n17406 & n18013) | (n17406 & n17900) | (n18013 & n17900);
  assign n17897 = n11315 & n17894;
  assign n17898 = (n17370 & n17901) | (n17370 & n17897) | (n17901 & n17897);
  assign n17440 = (n11206 & n11315) | (n11206 & n17898) | (n11315 & n17898);
  assign n17442 = n11315 & n17894;
  assign n17443 = (n17370 & n17901) | (n17370 & n17442) | (n17901 & n17442);
  assign n15148 = (n17430 & n17440) | (n17430 & n17443) | (n17440 & n17443);
  assign n17905 = n11203 | n11315;
  assign n18014 = (n11315 & n17400) | (n11315 & n17905) | (n17400 & n17905);
  assign n17906 = (n17406 & n18014) | (n17406 & n17905) | (n18014 & n17905);
  assign n17902 = n11315 | n17894;
  assign n17903 = (n17370 & n17906) | (n17370 & n17902) | (n17906 & n17902);
  assign n17445 = n11206 | n17903;
  assign n17447 = n11315 | n17894;
  assign n17448 = (n17370 & n17906) | (n17370 & n17447) | (n17906 & n17447);
  assign n15151 = (n17430 & n17445) | (n17430 & n17448) | (n17445 & n17448);
  assign n11318 = ~n15148 & n15151;
  assign n15152 = n11211 & n11318;
  assign n17449 = (n11318 & n15088) | (n11318 & n15152) | (n15088 & n15152);
  assign n17450 = (n11318 & n15087) | (n11318 & n15152) | (n15087 & n15152);
  assign n17451 = (n15006 & n17449) | (n15006 & n17450) | (n17449 & n17450);
  assign n15154 = n11211 | n11318;
  assign n17452 = n15088 | n15154;
  assign n17453 = n15087 | n15154;
  assign n17454 = (n15006 & n17452) | (n15006 & n17453) | (n17452 & n17453);
  assign n11321 = ~n17451 & n17454;
  assign n11322 = x78 & x100;
  assign n11323 = n11321 & n11322;
  assign n11324 = n11321 | n11322;
  assign n11325 = ~n11323 & n11324;
  assign n15142 = n11218 | n11220;
  assign n17455 = n11325 & n15142;
  assign n17437 = n11105 | n11218;
  assign n17438 = (n11218 & n11220) | (n11218 & n17437) | (n11220 & n17437);
  assign n17456 = n11325 & n17438;
  assign n17457 = (n17422 & n17455) | (n17422 & n17456) | (n17455 & n17456);
  assign n17458 = n11325 | n15142;
  assign n17459 = n11325 | n17438;
  assign n17460 = (n17422 & n17458) | (n17422 & n17459) | (n17458 & n17459);
  assign n11328 = ~n17457 & n17460;
  assign n11329 = x77 & x101;
  assign n11330 = n11328 & n11329;
  assign n11331 = n11328 | n11329;
  assign n11332 = ~n11330 & n11331;
  assign n15156 = n11225 & n11332;
  assign n17461 = (n11332 & n15097) | (n11332 & n15156) | (n15097 & n15156);
  assign n17462 = (n11227 & n11332) | (n11227 & n15156) | (n11332 & n15156);
  assign n17463 = (n15033 & n17461) | (n15033 & n17462) | (n17461 & n17462);
  assign n15158 = n11225 | n11332;
  assign n17464 = n15097 | n15158;
  assign n17465 = n11227 | n15158;
  assign n17466 = (n15033 & n17464) | (n15033 & n17465) | (n17464 & n17465);
  assign n11335 = ~n17463 & n17466;
  assign n11336 = x76 & x102;
  assign n11337 = n11335 & n11336;
  assign n11338 = n11335 | n11336;
  assign n11339 = ~n11337 & n11338;
  assign n15160 = n11232 & n11339;
  assign n15161 = (n11339 & n15102) | (n11339 & n15160) | (n15102 & n15160);
  assign n15162 = n11232 | n11339;
  assign n15163 = n15102 | n15162;
  assign n11342 = ~n15161 & n15163;
  assign n11343 = x75 & x103;
  assign n11344 = n11342 & n11343;
  assign n11345 = n11342 | n11343;
  assign n11346 = ~n11344 & n11345;
  assign n15164 = n11239 & n11346;
  assign n15165 = (n11346 & n15106) | (n11346 & n15164) | (n15106 & n15164);
  assign n15166 = n11239 | n11346;
  assign n15167 = n15106 | n15166;
  assign n11349 = ~n15165 & n15167;
  assign n11350 = x74 & x104;
  assign n11351 = n11349 & n11350;
  assign n11352 = n11349 | n11350;
  assign n11353 = ~n11351 & n11352;
  assign n15168 = n11246 & n11353;
  assign n15169 = (n11353 & n15110) | (n11353 & n15168) | (n15110 & n15168);
  assign n15170 = n11246 | n11353;
  assign n15171 = n15110 | n15170;
  assign n11356 = ~n15169 & n15171;
  assign n11357 = x73 & x105;
  assign n11358 = n11356 & n11357;
  assign n11359 = n11356 | n11357;
  assign n11360 = ~n11358 & n11359;
  assign n15172 = n11253 & n11360;
  assign n15173 = (n11360 & n15114) | (n11360 & n15172) | (n15114 & n15172);
  assign n15174 = n11253 | n11360;
  assign n15175 = n15114 | n15174;
  assign n11363 = ~n15173 & n15175;
  assign n11364 = x72 & x106;
  assign n11365 = n11363 & n11364;
  assign n11366 = n11363 | n11364;
  assign n11367 = ~n11365 & n11366;
  assign n15176 = n11260 & n11367;
  assign n15177 = (n11367 & n15118) | (n11367 & n15176) | (n15118 & n15176);
  assign n15178 = n11260 | n11367;
  assign n15179 = n15118 | n15178;
  assign n11370 = ~n15177 & n15179;
  assign n11371 = x71 & x107;
  assign n11372 = n11370 & n11371;
  assign n11373 = n11370 | n11371;
  assign n11374 = ~n11372 & n11373;
  assign n15180 = n11267 & n11374;
  assign n15181 = (n11374 & n15122) | (n11374 & n15180) | (n15122 & n15180);
  assign n15182 = n11267 | n11374;
  assign n15183 = n15122 | n15182;
  assign n11377 = ~n15181 & n15183;
  assign n11378 = x70 & x108;
  assign n11379 = n11377 & n11378;
  assign n11380 = n11377 | n11378;
  assign n11381 = ~n11379 & n11380;
  assign n15184 = n11274 & n11381;
  assign n15185 = (n11381 & n15126) | (n11381 & n15184) | (n15126 & n15184);
  assign n15186 = n11274 | n11381;
  assign n15187 = n15126 | n15186;
  assign n11384 = ~n15185 & n15187;
  assign n11385 = x69 & x109;
  assign n11386 = n11384 & n11385;
  assign n11387 = n11384 | n11385;
  assign n11388 = ~n11386 & n11387;
  assign n15188 = n11281 & n11388;
  assign n15189 = (n11388 & n15130) | (n11388 & n15188) | (n15130 & n15188);
  assign n15190 = n11281 | n11388;
  assign n15191 = n15130 | n15190;
  assign n11391 = ~n15189 & n15191;
  assign n11392 = x68 & x110;
  assign n11393 = n11391 & n11392;
  assign n11394 = n11391 | n11392;
  assign n11395 = ~n11393 & n11394;
  assign n15192 = n11288 & n11395;
  assign n15193 = (n11395 & n15134) | (n11395 & n15192) | (n15134 & n15192);
  assign n15194 = n11288 | n11395;
  assign n15195 = n15134 | n15194;
  assign n11398 = ~n15193 & n15195;
  assign n11399 = x67 & x111;
  assign n11400 = n11398 & n11399;
  assign n11401 = n11398 | n11399;
  assign n11402 = ~n11400 & n11401;
  assign n15196 = n11295 & n11402;
  assign n15197 = (n11402 & n15138) | (n11402 & n15196) | (n15138 & n15196);
  assign n15198 = n11295 | n11402;
  assign n15199 = n15138 | n15198;
  assign n11405 = ~n15197 & n15199;
  assign n11419 = x79 & x100;
  assign n15203 = n11318 | n15148;
  assign n17467 = (n11211 & n15148) | (n11211 & n15203) | (n15148 & n15203);
  assign n15205 = n11419 & n17467;
  assign n18109 = n11419 & n17900;
  assign n18173 = n17400 & n18109;
  assign n18110 = (n17406 & n18173) | (n17406 & n18109) | (n18173 & n18109);
  assign n18016 = n11315 & n11419;
  assign n18111 = n17894 & n18016;
  assign n18107 = (n17370 & n18110) | (n17370 & n18111) | (n18110 & n18111);
  assign n18017 = (n11206 & n18107) | (n11206 & n18016) | (n18107 & n18016);
  assign n18020 = (n17370 & n18110) | (n17370 & n18111) | (n18110 & n18111);
  assign n17909 = (n17430 & n18017) | (n17430 & n18020) | (n18017 & n18020);
  assign n17469 = (n11318 & n11419) | (n11318 & n17909) | (n11419 & n17909);
  assign n17470 = (n15088 & n15205) | (n15088 & n17469) | (n15205 & n17469);
  assign n17471 = (n15087 & n15205) | (n15087 & n17469) | (n15205 & n17469);
  assign n17472 = (n15006 & n17470) | (n15006 & n17471) | (n17470 & n17471);
  assign n15208 = n11419 | n17467;
  assign n18115 = n11419 | n17900;
  assign n18174 = (n11419 & n17400) | (n11419 & n18115) | (n17400 & n18115);
  assign n18116 = (n17406 & n18174) | (n17406 & n18115) | (n18174 & n18115);
  assign n18022 = n11315 | n11419;
  assign n18117 = (n11419 & n17894) | (n11419 & n18022) | (n17894 & n18022);
  assign n18113 = (n17370 & n18116) | (n17370 & n18117) | (n18116 & n18117);
  assign n18023 = (n11206 & n18113) | (n11206 & n18022) | (n18113 & n18022);
  assign n18026 = (n17370 & n18116) | (n17370 & n18117) | (n18116 & n18117);
  assign n17912 = (n17430 & n18023) | (n17430 & n18026) | (n18023 & n18026);
  assign n17474 = n11318 | n17912;
  assign n17475 = (n15088 & n15208) | (n15088 & n17474) | (n15208 & n17474);
  assign n17476 = (n15087 & n15208) | (n15087 & n17474) | (n15208 & n17474);
  assign n17477 = (n15006 & n17475) | (n15006 & n17476) | (n17475 & n17476);
  assign n11422 = ~n17472 & n17477;
  assign n15212 = n11323 & n11422;
  assign n17478 = (n11325 & n11422) | (n11325 & n15212) | (n11422 & n15212);
  assign n17479 = (n15142 & n15212) | (n15142 & n17478) | (n15212 & n17478);
  assign n17480 = (n15212 & n17438) | (n15212 & n17478) | (n17438 & n17478);
  assign n17481 = (n17422 & n17479) | (n17422 & n17480) | (n17479 & n17480);
  assign n15215 = n11323 | n11422;
  assign n17482 = n11325 | n15215;
  assign n17483 = (n15142 & n15215) | (n15142 & n17482) | (n15215 & n17482);
  assign n17484 = (n15215 & n17438) | (n15215 & n17482) | (n17438 & n17482);
  assign n17485 = (n17422 & n17483) | (n17422 & n17484) | (n17483 & n17484);
  assign n11425 = ~n17481 & n17485;
  assign n11426 = x78 & x101;
  assign n11427 = n11425 & n11426;
  assign n11428 = n11425 | n11426;
  assign n11429 = ~n11427 & n11428;
  assign n15217 = n11330 & n11429;
  assign n15218 = (n11429 & n17463) | (n11429 & n15217) | (n17463 & n15217);
  assign n15219 = n11330 | n11429;
  assign n15220 = n17463 | n15219;
  assign n11432 = ~n15218 & n15220;
  assign n11433 = x77 & x102;
  assign n11434 = n11432 & n11433;
  assign n11435 = n11432 | n11433;
  assign n11436 = ~n11434 & n11435;
  assign n15221 = n11337 & n11436;
  assign n15222 = (n11436 & n15161) | (n11436 & n15221) | (n15161 & n15221);
  assign n15223 = n11337 | n11436;
  assign n15224 = n15161 | n15223;
  assign n11439 = ~n15222 & n15224;
  assign n11440 = x76 & x103;
  assign n11441 = n11439 & n11440;
  assign n11442 = n11439 | n11440;
  assign n11443 = ~n11441 & n11442;
  assign n15225 = n11344 & n11443;
  assign n15226 = (n11443 & n15165) | (n11443 & n15225) | (n15165 & n15225);
  assign n15227 = n11344 | n11443;
  assign n15228 = n15165 | n15227;
  assign n11446 = ~n15226 & n15228;
  assign n11447 = x75 & x104;
  assign n11448 = n11446 & n11447;
  assign n11449 = n11446 | n11447;
  assign n11450 = ~n11448 & n11449;
  assign n15229 = n11351 & n11450;
  assign n15230 = (n11450 & n15169) | (n11450 & n15229) | (n15169 & n15229);
  assign n15231 = n11351 | n11450;
  assign n15232 = n15169 | n15231;
  assign n11453 = ~n15230 & n15232;
  assign n11454 = x74 & x105;
  assign n11455 = n11453 & n11454;
  assign n11456 = n11453 | n11454;
  assign n11457 = ~n11455 & n11456;
  assign n15233 = n11358 & n11457;
  assign n15234 = (n11457 & n15173) | (n11457 & n15233) | (n15173 & n15233);
  assign n15235 = n11358 | n11457;
  assign n15236 = n15173 | n15235;
  assign n11460 = ~n15234 & n15236;
  assign n11461 = x73 & x106;
  assign n11462 = n11460 & n11461;
  assign n11463 = n11460 | n11461;
  assign n11464 = ~n11462 & n11463;
  assign n15237 = n11365 & n11464;
  assign n15238 = (n11464 & n15177) | (n11464 & n15237) | (n15177 & n15237);
  assign n15239 = n11365 | n11464;
  assign n15240 = n15177 | n15239;
  assign n11467 = ~n15238 & n15240;
  assign n11468 = x72 & x107;
  assign n11469 = n11467 & n11468;
  assign n11470 = n11467 | n11468;
  assign n11471 = ~n11469 & n11470;
  assign n15241 = n11372 & n11471;
  assign n15242 = (n11471 & n15181) | (n11471 & n15241) | (n15181 & n15241);
  assign n15243 = n11372 | n11471;
  assign n15244 = n15181 | n15243;
  assign n11474 = ~n15242 & n15244;
  assign n11475 = x71 & x108;
  assign n11476 = n11474 & n11475;
  assign n11477 = n11474 | n11475;
  assign n11478 = ~n11476 & n11477;
  assign n15245 = n11379 & n11478;
  assign n15246 = (n11478 & n15185) | (n11478 & n15245) | (n15185 & n15245);
  assign n15247 = n11379 | n11478;
  assign n15248 = n15185 | n15247;
  assign n11481 = ~n15246 & n15248;
  assign n11482 = x70 & x109;
  assign n11483 = n11481 & n11482;
  assign n11484 = n11481 | n11482;
  assign n11485 = ~n11483 & n11484;
  assign n15249 = n11386 & n11485;
  assign n15250 = (n11485 & n15189) | (n11485 & n15249) | (n15189 & n15249);
  assign n15251 = n11386 | n11485;
  assign n15252 = n15189 | n15251;
  assign n11488 = ~n15250 & n15252;
  assign n11489 = x69 & x110;
  assign n11490 = n11488 & n11489;
  assign n11491 = n11488 | n11489;
  assign n11492 = ~n11490 & n11491;
  assign n15253 = n11393 & n11492;
  assign n15254 = (n11492 & n15193) | (n11492 & n15253) | (n15193 & n15253);
  assign n15255 = n11393 | n11492;
  assign n15256 = n15193 | n15255;
  assign n11495 = ~n15254 & n15256;
  assign n11496 = x68 & x111;
  assign n11497 = n11495 & n11496;
  assign n11498 = n11495 | n11496;
  assign n11499 = ~n11497 & n11498;
  assign n15257 = n11400 & n11499;
  assign n15258 = (n11499 & n15197) | (n11499 & n15257) | (n15197 & n15257);
  assign n15259 = n11400 | n11499;
  assign n15260 = n15197 | n15259;
  assign n11502 = ~n15258 & n15260;
  assign n11515 = x79 & x101;
  assign n15264 = n11515 & n17472;
  assign n15265 = (n11515 & n17481) | (n11515 & n15264) | (n17481 & n15264);
  assign n15266 = n11515 | n17472;
  assign n15267 = n17481 | n15266;
  assign n11518 = ~n15265 & n15267;
  assign n17913 = n11427 & n11518;
  assign n17914 = (n11429 & n11518) | (n11429 & n17913) | (n11518 & n17913);
  assign n17486 = n11330 | n11427;
  assign n17487 = (n11427 & n11429) | (n11427 & n17486) | (n11429 & n17486);
  assign n17489 = n11518 & n17487;
  assign n17490 = (n17463 & n17914) | (n17463 & n17489) | (n17914 & n17489);
  assign n17915 = n11427 | n11518;
  assign n17916 = n11429 | n17915;
  assign n17492 = n11518 | n17487;
  assign n17493 = (n17463 & n17916) | (n17463 & n17492) | (n17916 & n17492);
  assign n11521 = ~n17490 & n17493;
  assign n11522 = x78 & x102;
  assign n11523 = n11521 & n11522;
  assign n11524 = n11521 | n11522;
  assign n11525 = ~n11523 & n11524;
  assign n15268 = n11434 & n11525;
  assign n17494 = (n11525 & n15221) | (n11525 & n15268) | (n15221 & n15268);
  assign n17495 = (n11436 & n11525) | (n11436 & n15268) | (n11525 & n15268);
  assign n17496 = (n15161 & n17494) | (n15161 & n17495) | (n17494 & n17495);
  assign n15270 = n11434 | n11525;
  assign n17497 = n15221 | n15270;
  assign n17498 = n11436 | n15270;
  assign n17499 = (n15161 & n17497) | (n15161 & n17498) | (n17497 & n17498);
  assign n11528 = ~n17496 & n17499;
  assign n11529 = x77 & x103;
  assign n11530 = n11528 & n11529;
  assign n11531 = n11528 | n11529;
  assign n11532 = ~n11530 & n11531;
  assign n15272 = n11441 & n11532;
  assign n15273 = (n11532 & n15226) | (n11532 & n15272) | (n15226 & n15272);
  assign n15274 = n11441 | n11532;
  assign n15275 = n15226 | n15274;
  assign n11535 = ~n15273 & n15275;
  assign n11536 = x76 & x104;
  assign n11537 = n11535 & n11536;
  assign n11538 = n11535 | n11536;
  assign n11539 = ~n11537 & n11538;
  assign n15276 = n11448 & n11539;
  assign n15277 = (n11539 & n15230) | (n11539 & n15276) | (n15230 & n15276);
  assign n15278 = n11448 | n11539;
  assign n15279 = n15230 | n15278;
  assign n11542 = ~n15277 & n15279;
  assign n11543 = x75 & x105;
  assign n11544 = n11542 & n11543;
  assign n11545 = n11542 | n11543;
  assign n11546 = ~n11544 & n11545;
  assign n15280 = n11455 & n11546;
  assign n15281 = (n11546 & n15234) | (n11546 & n15280) | (n15234 & n15280);
  assign n15282 = n11455 | n11546;
  assign n15283 = n15234 | n15282;
  assign n11549 = ~n15281 & n15283;
  assign n11550 = x74 & x106;
  assign n11551 = n11549 & n11550;
  assign n11552 = n11549 | n11550;
  assign n11553 = ~n11551 & n11552;
  assign n15284 = n11462 & n11553;
  assign n15285 = (n11553 & n15238) | (n11553 & n15284) | (n15238 & n15284);
  assign n15286 = n11462 | n11553;
  assign n15287 = n15238 | n15286;
  assign n11556 = ~n15285 & n15287;
  assign n11557 = x73 & x107;
  assign n11558 = n11556 & n11557;
  assign n11559 = n11556 | n11557;
  assign n11560 = ~n11558 & n11559;
  assign n15288 = n11469 & n11560;
  assign n15289 = (n11560 & n15242) | (n11560 & n15288) | (n15242 & n15288);
  assign n15290 = n11469 | n11560;
  assign n15291 = n15242 | n15290;
  assign n11563 = ~n15289 & n15291;
  assign n11564 = x72 & x108;
  assign n11565 = n11563 & n11564;
  assign n11566 = n11563 | n11564;
  assign n11567 = ~n11565 & n11566;
  assign n15292 = n11476 & n11567;
  assign n15293 = (n11567 & n15246) | (n11567 & n15292) | (n15246 & n15292);
  assign n15294 = n11476 | n11567;
  assign n15295 = n15246 | n15294;
  assign n11570 = ~n15293 & n15295;
  assign n11571 = x71 & x109;
  assign n11572 = n11570 & n11571;
  assign n11573 = n11570 | n11571;
  assign n11574 = ~n11572 & n11573;
  assign n15296 = n11483 & n11574;
  assign n15297 = (n11574 & n15250) | (n11574 & n15296) | (n15250 & n15296);
  assign n15298 = n11483 | n11574;
  assign n15299 = n15250 | n15298;
  assign n11577 = ~n15297 & n15299;
  assign n11578 = x70 & x110;
  assign n11579 = n11577 & n11578;
  assign n11580 = n11577 | n11578;
  assign n11581 = ~n11579 & n11580;
  assign n15300 = n11490 & n11581;
  assign n15301 = (n11581 & n15254) | (n11581 & n15300) | (n15254 & n15300);
  assign n15302 = n11490 | n11581;
  assign n15303 = n15254 | n15302;
  assign n11584 = ~n15301 & n15303;
  assign n11585 = x69 & x111;
  assign n11586 = n11584 & n11585;
  assign n11587 = n11584 | n11585;
  assign n11588 = ~n11586 & n11587;
  assign n15304 = n11497 & n11588;
  assign n15305 = (n11588 & n15258) | (n11588 & n15304) | (n15258 & n15304);
  assign n15306 = n11497 | n11588;
  assign n15307 = n15258 | n15306;
  assign n11591 = ~n15305 & n15307;
  assign n15262 = n11427 | n11429;
  assign n11603 = x79 & x102;
  assign n17502 = n11515 & n11603;
  assign n17917 = n17472 & n17502;
  assign n17503 = (n17481 & n17917) | (n17481 & n17502) | (n17917 & n17502);
  assign n17500 = (n11518 & n11603) | (n11518 & n17503) | (n11603 & n17503);
  assign n17504 = (n15262 & n17500) | (n15262 & n17503) | (n17500 & n17503);
  assign n17505 = (n17487 & n17500) | (n17487 & n17503) | (n17500 & n17503);
  assign n17506 = (n17463 & n17504) | (n17463 & n17505) | (n17504 & n17505);
  assign n17509 = n11515 | n11603;
  assign n17918 = (n11603 & n17472) | (n11603 & n17509) | (n17472 & n17509);
  assign n17510 = (n17481 & n17918) | (n17481 & n17509) | (n17918 & n17509);
  assign n17507 = n11518 | n17510;
  assign n17511 = (n15262 & n17507) | (n15262 & n17510) | (n17507 & n17510);
  assign n17512 = (n17487 & n17507) | (n17487 & n17510) | (n17507 & n17510);
  assign n17513 = (n17463 & n17511) | (n17463 & n17512) | (n17511 & n17512);
  assign n11606 = ~n17506 & n17513;
  assign n15316 = n11523 & n11606;
  assign n15317 = (n11606 & n17496) | (n11606 & n15316) | (n17496 & n15316);
  assign n15318 = n11523 | n11606;
  assign n15319 = n17496 | n15318;
  assign n11609 = ~n15317 & n15319;
  assign n11610 = x78 & x103;
  assign n11611 = n11609 & n11610;
  assign n11612 = n11609 | n11610;
  assign n11613 = ~n11611 & n11612;
  assign n15320 = n11530 & n11613;
  assign n15321 = (n11613 & n15273) | (n11613 & n15320) | (n15273 & n15320);
  assign n15322 = n11530 | n11613;
  assign n15323 = n15273 | n15322;
  assign n11616 = ~n15321 & n15323;
  assign n11617 = x77 & x104;
  assign n11618 = n11616 & n11617;
  assign n11619 = n11616 | n11617;
  assign n11620 = ~n11618 & n11619;
  assign n15324 = n11537 & n11620;
  assign n15325 = (n11620 & n15277) | (n11620 & n15324) | (n15277 & n15324);
  assign n15326 = n11537 | n11620;
  assign n15327 = n15277 | n15326;
  assign n11623 = ~n15325 & n15327;
  assign n11624 = x76 & x105;
  assign n11625 = n11623 & n11624;
  assign n11626 = n11623 | n11624;
  assign n11627 = ~n11625 & n11626;
  assign n15328 = n11544 & n11627;
  assign n15329 = (n11627 & n15281) | (n11627 & n15328) | (n15281 & n15328);
  assign n15330 = n11544 | n11627;
  assign n15331 = n15281 | n15330;
  assign n11630 = ~n15329 & n15331;
  assign n11631 = x75 & x106;
  assign n11632 = n11630 & n11631;
  assign n11633 = n11630 | n11631;
  assign n11634 = ~n11632 & n11633;
  assign n15332 = n11551 & n11634;
  assign n15333 = (n11634 & n15285) | (n11634 & n15332) | (n15285 & n15332);
  assign n15334 = n11551 | n11634;
  assign n15335 = n15285 | n15334;
  assign n11637 = ~n15333 & n15335;
  assign n11638 = x74 & x107;
  assign n11639 = n11637 & n11638;
  assign n11640 = n11637 | n11638;
  assign n11641 = ~n11639 & n11640;
  assign n15336 = n11558 & n11641;
  assign n15337 = (n11641 & n15289) | (n11641 & n15336) | (n15289 & n15336);
  assign n15338 = n11558 | n11641;
  assign n15339 = n15289 | n15338;
  assign n11644 = ~n15337 & n15339;
  assign n11645 = x73 & x108;
  assign n11646 = n11644 & n11645;
  assign n11647 = n11644 | n11645;
  assign n11648 = ~n11646 & n11647;
  assign n15340 = n11565 & n11648;
  assign n15341 = (n11648 & n15293) | (n11648 & n15340) | (n15293 & n15340);
  assign n15342 = n11565 | n11648;
  assign n15343 = n15293 | n15342;
  assign n11651 = ~n15341 & n15343;
  assign n11652 = x72 & x109;
  assign n11653 = n11651 & n11652;
  assign n11654 = n11651 | n11652;
  assign n11655 = ~n11653 & n11654;
  assign n15344 = n11572 & n11655;
  assign n15345 = (n11655 & n15297) | (n11655 & n15344) | (n15297 & n15344);
  assign n15346 = n11572 | n11655;
  assign n15347 = n15297 | n15346;
  assign n11658 = ~n15345 & n15347;
  assign n11659 = x71 & x110;
  assign n11660 = n11658 & n11659;
  assign n11661 = n11658 | n11659;
  assign n11662 = ~n11660 & n11661;
  assign n15348 = n11579 & n11662;
  assign n15349 = (n11662 & n15301) | (n11662 & n15348) | (n15301 & n15348);
  assign n15350 = n11579 | n11662;
  assign n15351 = n15301 | n15350;
  assign n11665 = ~n15349 & n15351;
  assign n11666 = x70 & x111;
  assign n11667 = n11665 & n11666;
  assign n11668 = n11665 | n11666;
  assign n11669 = ~n11667 & n11668;
  assign n15352 = n11586 & n11669;
  assign n15353 = (n11669 & n15305) | (n11669 & n15352) | (n15305 & n15352);
  assign n15354 = n11586 | n11669;
  assign n15355 = n15305 | n15354;
  assign n11672 = ~n15353 & n15355;
  assign n11683 = x79 & x103;
  assign n17514 = n11606 | n17506;
  assign n17515 = (n11523 & n17506) | (n11523 & n17514) | (n17506 & n17514);
  assign n15359 = n11683 & n17515;
  assign n18121 = n11683 & n17502;
  assign n18175 = n17472 & n18121;
  assign n18122 = (n17481 & n18175) | (n17481 & n18121) | (n18175 & n18121);
  assign n18118 = n11603 & n11683;
  assign n18119 = (n11518 & n18122) | (n11518 & n18118) | (n18122 & n18118);
  assign n18029 = (n17487 & n18119) | (n17487 & n18122) | (n18119 & n18122);
  assign n18030 = (n15262 & n18119) | (n15262 & n18122) | (n18119 & n18122);
  assign n17921 = (n17463 & n18029) | (n17463 & n18030) | (n18029 & n18030);
  assign n17517 = (n11606 & n11683) | (n11606 & n17921) | (n11683 & n17921);
  assign n15361 = (n17496 & n15359) | (n17496 & n17517) | (n15359 & n17517);
  assign n15362 = n11683 | n17515;
  assign n18126 = n11683 | n17502;
  assign n18176 = (n11683 & n17472) | (n11683 & n18126) | (n17472 & n18126);
  assign n18127 = (n17481 & n18176) | (n17481 & n18126) | (n18176 & n18126);
  assign n18123 = n11603 | n11683;
  assign n18124 = (n11518 & n18127) | (n11518 & n18123) | (n18127 & n18123);
  assign n18033 = (n17487 & n18124) | (n17487 & n18127) | (n18124 & n18127);
  assign n18034 = (n15262 & n18124) | (n15262 & n18127) | (n18124 & n18127);
  assign n17924 = (n17463 & n18033) | (n17463 & n18034) | (n18033 & n18034);
  assign n17519 = n11606 | n17924;
  assign n15364 = (n17496 & n15362) | (n17496 & n17519) | (n15362 & n17519);
  assign n11686 = ~n15361 & n15364;
  assign n15365 = n11611 & n11686;
  assign n17520 = (n11686 & n15320) | (n11686 & n15365) | (n15320 & n15365);
  assign n17521 = (n11613 & n11686) | (n11613 & n15365) | (n11686 & n15365);
  assign n17522 = (n15273 & n17520) | (n15273 & n17521) | (n17520 & n17521);
  assign n15367 = n11611 | n11686;
  assign n17523 = n15320 | n15367;
  assign n17524 = n11613 | n15367;
  assign n17525 = (n15273 & n17523) | (n15273 & n17524) | (n17523 & n17524);
  assign n11689 = ~n17522 & n17525;
  assign n11690 = x78 & x104;
  assign n11691 = n11689 & n11690;
  assign n11692 = n11689 | n11690;
  assign n11693 = ~n11691 & n11692;
  assign n15369 = n11618 & n11693;
  assign n15370 = (n11693 & n15325) | (n11693 & n15369) | (n15325 & n15369);
  assign n15371 = n11618 | n11693;
  assign n15372 = n15325 | n15371;
  assign n11696 = ~n15370 & n15372;
  assign n11697 = x77 & x105;
  assign n11698 = n11696 & n11697;
  assign n11699 = n11696 | n11697;
  assign n11700 = ~n11698 & n11699;
  assign n15373 = n11625 & n11700;
  assign n15374 = (n11700 & n15329) | (n11700 & n15373) | (n15329 & n15373);
  assign n15375 = n11625 | n11700;
  assign n15376 = n15329 | n15375;
  assign n11703 = ~n15374 & n15376;
  assign n11704 = x76 & x106;
  assign n11705 = n11703 & n11704;
  assign n11706 = n11703 | n11704;
  assign n11707 = ~n11705 & n11706;
  assign n15377 = n11632 & n11707;
  assign n15378 = (n11707 & n15333) | (n11707 & n15377) | (n15333 & n15377);
  assign n15379 = n11632 | n11707;
  assign n15380 = n15333 | n15379;
  assign n11710 = ~n15378 & n15380;
  assign n11711 = x75 & x107;
  assign n11712 = n11710 & n11711;
  assign n11713 = n11710 | n11711;
  assign n11714 = ~n11712 & n11713;
  assign n15381 = n11639 & n11714;
  assign n15382 = (n11714 & n15337) | (n11714 & n15381) | (n15337 & n15381);
  assign n15383 = n11639 | n11714;
  assign n15384 = n15337 | n15383;
  assign n11717 = ~n15382 & n15384;
  assign n11718 = x74 & x108;
  assign n11719 = n11717 & n11718;
  assign n11720 = n11717 | n11718;
  assign n11721 = ~n11719 & n11720;
  assign n15385 = n11646 & n11721;
  assign n15386 = (n11721 & n15341) | (n11721 & n15385) | (n15341 & n15385);
  assign n15387 = n11646 | n11721;
  assign n15388 = n15341 | n15387;
  assign n11724 = ~n15386 & n15388;
  assign n11725 = x73 & x109;
  assign n11726 = n11724 & n11725;
  assign n11727 = n11724 | n11725;
  assign n11728 = ~n11726 & n11727;
  assign n15389 = n11653 & n11728;
  assign n15390 = (n11728 & n15345) | (n11728 & n15389) | (n15345 & n15389);
  assign n15391 = n11653 | n11728;
  assign n15392 = n15345 | n15391;
  assign n11731 = ~n15390 & n15392;
  assign n11732 = x72 & x110;
  assign n11733 = n11731 & n11732;
  assign n11734 = n11731 | n11732;
  assign n11735 = ~n11733 & n11734;
  assign n15393 = n11660 & n11735;
  assign n15394 = (n11735 & n15349) | (n11735 & n15393) | (n15349 & n15393);
  assign n15395 = n11660 | n11735;
  assign n15396 = n15349 | n15395;
  assign n11738 = ~n15394 & n15396;
  assign n11739 = x71 & x111;
  assign n11740 = n11738 & n11739;
  assign n11741 = n11738 | n11739;
  assign n11742 = ~n11740 & n11741;
  assign n15397 = n11667 & n11742;
  assign n15398 = (n11742 & n15353) | (n11742 & n15397) | (n15353 & n15397);
  assign n15399 = n11667 | n11742;
  assign n15400 = n15353 | n15399;
  assign n11745 = ~n15398 & n15400;
  assign n11755 = x79 & x104;
  assign n15402 = n11686 | n15361;
  assign n17526 = (n11611 & n15361) | (n11611 & n15402) | (n15361 & n15402);
  assign n15404 = n11755 & n17526;
  assign n18035 = n11683 & n11755;
  assign n18036 = n17515 & n18035;
  assign n18240 = n17502 & n18035;
  assign n18239 = n17472 & n18240;
  assign n18215 = (n17481 & n18239) | (n17481 & n18240) | (n18239 & n18240);
  assign n18211 = n11755 & n18118;
  assign n18212 = (n11518 & n18215) | (n11518 & n18211) | (n18215 & n18211);
  assign n18179 = (n15262 & n18212) | (n15262 & n18215) | (n18212 & n18215);
  assign n18180 = (n17487 & n18212) | (n17487 & n18215) | (n18212 & n18215);
  assign n18130 = (n17463 & n18179) | (n17463 & n18180) | (n18179 & n18180);
  assign n18038 = (n11606 & n18035) | (n11606 & n18130) | (n18035 & n18130);
  assign n17927 = (n17496 & n18036) | (n17496 & n18038) | (n18036 & n18038);
  assign n17528 = (n11686 & n11755) | (n11686 & n17927) | (n11755 & n17927);
  assign n17529 = (n15320 & n15404) | (n15320 & n17528) | (n15404 & n17528);
  assign n17530 = (n11613 & n15404) | (n11613 & n17528) | (n15404 & n17528);
  assign n17531 = (n15273 & n17529) | (n15273 & n17530) | (n17529 & n17530);
  assign n15407 = n11755 | n17526;
  assign n18039 = n11683 | n11755;
  assign n18040 = (n11755 & n17515) | (n11755 & n18039) | (n17515 & n18039);
  assign n18242 = (n11755 & n17502) | (n11755 & n18039) | (n17502 & n18039);
  assign n18241 = (n11755 & n17472) | (n11755 & n18242) | (n17472 & n18242);
  assign n18220 = (n17481 & n18241) | (n17481 & n18242) | (n18241 & n18242);
  assign n18216 = n11755 | n18118;
  assign n18217 = (n11518 & n18220) | (n11518 & n18216) | (n18220 & n18216);
  assign n18183 = (n15262 & n18217) | (n15262 & n18220) | (n18217 & n18220);
  assign n18184 = (n17487 & n18217) | (n17487 & n18220) | (n18217 & n18220);
  assign n18133 = (n17463 & n18183) | (n17463 & n18184) | (n18183 & n18184);
  assign n18042 = (n11606 & n18039) | (n11606 & n18133) | (n18039 & n18133);
  assign n17930 = (n17496 & n18040) | (n17496 & n18042) | (n18040 & n18042);
  assign n17533 = n11686 | n17930;
  assign n17534 = (n15320 & n15407) | (n15320 & n17533) | (n15407 & n17533);
  assign n17535 = (n11613 & n15407) | (n11613 & n17533) | (n15407 & n17533);
  assign n17536 = (n15273 & n17534) | (n15273 & n17535) | (n17534 & n17535);
  assign n11758 = ~n17531 & n17536;
  assign n15410 = n11691 & n11758;
  assign n17537 = (n11758 & n15369) | (n11758 & n15410) | (n15369 & n15410);
  assign n17538 = (n11693 & n11758) | (n11693 & n15410) | (n11758 & n15410);
  assign n17539 = (n15325 & n17537) | (n15325 & n17538) | (n17537 & n17538);
  assign n15412 = n11691 | n11758;
  assign n17540 = n15369 | n15412;
  assign n17541 = n11693 | n15412;
  assign n17542 = (n15325 & n17540) | (n15325 & n17541) | (n17540 & n17541);
  assign n11761 = ~n17539 & n17542;
  assign n11762 = x78 & x105;
  assign n11763 = n11761 & n11762;
  assign n11764 = n11761 | n11762;
  assign n11765 = ~n11763 & n11764;
  assign n15414 = n11698 & n11765;
  assign n15415 = (n11765 & n15374) | (n11765 & n15414) | (n15374 & n15414);
  assign n15416 = n11698 | n11765;
  assign n15417 = n15374 | n15416;
  assign n11768 = ~n15415 & n15417;
  assign n11769 = x77 & x106;
  assign n11770 = n11768 & n11769;
  assign n11771 = n11768 | n11769;
  assign n11772 = ~n11770 & n11771;
  assign n15418 = n11705 & n11772;
  assign n15419 = (n11772 & n15378) | (n11772 & n15418) | (n15378 & n15418);
  assign n15420 = n11705 | n11772;
  assign n15421 = n15378 | n15420;
  assign n11775 = ~n15419 & n15421;
  assign n11776 = x76 & x107;
  assign n11777 = n11775 & n11776;
  assign n11778 = n11775 | n11776;
  assign n11779 = ~n11777 & n11778;
  assign n15422 = n11712 & n11779;
  assign n15423 = (n11779 & n15382) | (n11779 & n15422) | (n15382 & n15422);
  assign n15424 = n11712 | n11779;
  assign n15425 = n15382 | n15424;
  assign n11782 = ~n15423 & n15425;
  assign n11783 = x75 & x108;
  assign n11784 = n11782 & n11783;
  assign n11785 = n11782 | n11783;
  assign n11786 = ~n11784 & n11785;
  assign n15426 = n11719 & n11786;
  assign n15427 = (n11786 & n15386) | (n11786 & n15426) | (n15386 & n15426);
  assign n15428 = n11719 | n11786;
  assign n15429 = n15386 | n15428;
  assign n11789 = ~n15427 & n15429;
  assign n11790 = x74 & x109;
  assign n11791 = n11789 & n11790;
  assign n11792 = n11789 | n11790;
  assign n11793 = ~n11791 & n11792;
  assign n15430 = n11726 & n11793;
  assign n15431 = (n11793 & n15390) | (n11793 & n15430) | (n15390 & n15430);
  assign n15432 = n11726 | n11793;
  assign n15433 = n15390 | n15432;
  assign n11796 = ~n15431 & n15433;
  assign n11797 = x73 & x110;
  assign n11798 = n11796 & n11797;
  assign n11799 = n11796 | n11797;
  assign n11800 = ~n11798 & n11799;
  assign n15434 = n11733 & n11800;
  assign n15435 = (n11800 & n15394) | (n11800 & n15434) | (n15394 & n15434);
  assign n15436 = n11733 | n11800;
  assign n15437 = n15394 | n15436;
  assign n11803 = ~n15435 & n15437;
  assign n11804 = x72 & x111;
  assign n11805 = n11803 & n11804;
  assign n11806 = n11803 | n11804;
  assign n11807 = ~n11805 & n11806;
  assign n15438 = n11740 & n11807;
  assign n15439 = (n11807 & n15398) | (n11807 & n15438) | (n15398 & n15438);
  assign n15440 = n11740 | n11807;
  assign n15441 = n15398 | n15440;
  assign n11810 = ~n15439 & n15441;
  assign n11819 = x79 & x105;
  assign n17543 = n11758 | n17531;
  assign n17544 = (n11691 & n17531) | (n11691 & n17543) | (n17531 & n17543);
  assign n15445 = n11819 & n17544;
  assign n17545 = n11819 & n17531;
  assign n17546 = (n11758 & n11819) | (n11758 & n17545) | (n11819 & n17545);
  assign n17547 = (n15369 & n15445) | (n15369 & n17546) | (n15445 & n17546);
  assign n17548 = (n11693 & n15445) | (n11693 & n17546) | (n15445 & n17546);
  assign n17549 = (n15325 & n17547) | (n15325 & n17548) | (n17547 & n17548);
  assign n15448 = n11819 | n17544;
  assign n17550 = n11819 | n17531;
  assign n17551 = n11758 | n17550;
  assign n17552 = (n15369 & n15448) | (n15369 & n17551) | (n15448 & n17551);
  assign n17553 = (n11693 & n15448) | (n11693 & n17551) | (n15448 & n17551);
  assign n17554 = (n15325 & n17552) | (n15325 & n17553) | (n17552 & n17553);
  assign n11822 = ~n17549 & n17554;
  assign n15451 = n11763 & n11822;
  assign n17555 = (n11822 & n15414) | (n11822 & n15451) | (n15414 & n15451);
  assign n17556 = (n11765 & n11822) | (n11765 & n15451) | (n11822 & n15451);
  assign n17557 = (n15374 & n17555) | (n15374 & n17556) | (n17555 & n17556);
  assign n15453 = n11763 | n11822;
  assign n17558 = n15414 | n15453;
  assign n17559 = n11765 | n15453;
  assign n17560 = (n15374 & n17558) | (n15374 & n17559) | (n17558 & n17559);
  assign n11825 = ~n17557 & n17560;
  assign n11826 = x78 & x106;
  assign n11827 = n11825 & n11826;
  assign n11828 = n11825 | n11826;
  assign n11829 = ~n11827 & n11828;
  assign n15455 = n11770 & n11829;
  assign n15456 = (n11829 & n15419) | (n11829 & n15455) | (n15419 & n15455);
  assign n15457 = n11770 | n11829;
  assign n15458 = n15419 | n15457;
  assign n11832 = ~n15456 & n15458;
  assign n11833 = x77 & x107;
  assign n11834 = n11832 & n11833;
  assign n11835 = n11832 | n11833;
  assign n11836 = ~n11834 & n11835;
  assign n15459 = n11777 & n11836;
  assign n15460 = (n11836 & n15423) | (n11836 & n15459) | (n15423 & n15459);
  assign n15461 = n11777 | n11836;
  assign n15462 = n15423 | n15461;
  assign n11839 = ~n15460 & n15462;
  assign n11840 = x76 & x108;
  assign n11841 = n11839 & n11840;
  assign n11842 = n11839 | n11840;
  assign n11843 = ~n11841 & n11842;
  assign n15463 = n11784 & n11843;
  assign n15464 = (n11843 & n15427) | (n11843 & n15463) | (n15427 & n15463);
  assign n15465 = n11784 | n11843;
  assign n15466 = n15427 | n15465;
  assign n11846 = ~n15464 & n15466;
  assign n11847 = x75 & x109;
  assign n11848 = n11846 & n11847;
  assign n11849 = n11846 | n11847;
  assign n11850 = ~n11848 & n11849;
  assign n15467 = n11791 & n11850;
  assign n15468 = (n11850 & n15431) | (n11850 & n15467) | (n15431 & n15467);
  assign n15469 = n11791 | n11850;
  assign n15470 = n15431 | n15469;
  assign n11853 = ~n15468 & n15470;
  assign n11854 = x74 & x110;
  assign n11855 = n11853 & n11854;
  assign n11856 = n11853 | n11854;
  assign n11857 = ~n11855 & n11856;
  assign n15471 = n11798 & n11857;
  assign n15472 = (n11857 & n15435) | (n11857 & n15471) | (n15435 & n15471);
  assign n15473 = n11798 | n11857;
  assign n15474 = n15435 | n15473;
  assign n11860 = ~n15472 & n15474;
  assign n11861 = x73 & x111;
  assign n11862 = n11860 & n11861;
  assign n11863 = n11860 | n11861;
  assign n11864 = ~n11862 & n11863;
  assign n15475 = n11805 & n11864;
  assign n15476 = (n11864 & n15439) | (n11864 & n15475) | (n15439 & n15475);
  assign n15477 = n11805 | n11864;
  assign n15478 = n15439 | n15477;
  assign n11867 = ~n15476 & n15478;
  assign n11875 = x79 & x106;
  assign n17561 = n11822 | n17549;
  assign n17562 = (n11763 & n17549) | (n11763 & n17561) | (n17549 & n17561);
  assign n15482 = n11875 & n17562;
  assign n17563 = n11875 & n17549;
  assign n17564 = (n11822 & n11875) | (n11822 & n17563) | (n11875 & n17563);
  assign n17565 = (n15414 & n15482) | (n15414 & n17564) | (n15482 & n17564);
  assign n17566 = (n11765 & n15482) | (n11765 & n17564) | (n15482 & n17564);
  assign n17567 = (n15374 & n17565) | (n15374 & n17566) | (n17565 & n17566);
  assign n15485 = n11875 | n17562;
  assign n17568 = n11875 | n17549;
  assign n17569 = n11822 | n17568;
  assign n17570 = (n15414 & n15485) | (n15414 & n17569) | (n15485 & n17569);
  assign n17571 = (n11765 & n15485) | (n11765 & n17569) | (n15485 & n17569);
  assign n17572 = (n15374 & n17570) | (n15374 & n17571) | (n17570 & n17571);
  assign n11878 = ~n17567 & n17572;
  assign n15488 = n11827 & n11878;
  assign n17573 = (n11878 & n15455) | (n11878 & n15488) | (n15455 & n15488);
  assign n17574 = (n11829 & n11878) | (n11829 & n15488) | (n11878 & n15488);
  assign n17575 = (n15419 & n17573) | (n15419 & n17574) | (n17573 & n17574);
  assign n15490 = n11827 | n11878;
  assign n17576 = n15455 | n15490;
  assign n17577 = n11829 | n15490;
  assign n17578 = (n15419 & n17576) | (n15419 & n17577) | (n17576 & n17577);
  assign n11881 = ~n17575 & n17578;
  assign n11882 = x78 & x107;
  assign n11883 = n11881 & n11882;
  assign n11884 = n11881 | n11882;
  assign n11885 = ~n11883 & n11884;
  assign n15492 = n11834 & n11885;
  assign n15493 = (n11885 & n15460) | (n11885 & n15492) | (n15460 & n15492);
  assign n15494 = n11834 | n11885;
  assign n15495 = n15460 | n15494;
  assign n11888 = ~n15493 & n15495;
  assign n11889 = x77 & x108;
  assign n11890 = n11888 & n11889;
  assign n11891 = n11888 | n11889;
  assign n11892 = ~n11890 & n11891;
  assign n15496 = n11841 & n11892;
  assign n15497 = (n11892 & n15464) | (n11892 & n15496) | (n15464 & n15496);
  assign n15498 = n11841 | n11892;
  assign n15499 = n15464 | n15498;
  assign n11895 = ~n15497 & n15499;
  assign n11896 = x76 & x109;
  assign n11897 = n11895 & n11896;
  assign n11898 = n11895 | n11896;
  assign n11899 = ~n11897 & n11898;
  assign n15500 = n11848 & n11899;
  assign n15501 = (n11899 & n15468) | (n11899 & n15500) | (n15468 & n15500);
  assign n15502 = n11848 | n11899;
  assign n15503 = n15468 | n15502;
  assign n11902 = ~n15501 & n15503;
  assign n11903 = x75 & x110;
  assign n11904 = n11902 & n11903;
  assign n11905 = n11902 | n11903;
  assign n11906 = ~n11904 & n11905;
  assign n15504 = n11855 & n11906;
  assign n15505 = (n11906 & n15472) | (n11906 & n15504) | (n15472 & n15504);
  assign n15506 = n11855 | n11906;
  assign n15507 = n15472 | n15506;
  assign n11909 = ~n15505 & n15507;
  assign n11910 = x74 & x111;
  assign n11911 = n11909 & n11910;
  assign n11912 = n11909 | n11910;
  assign n11913 = ~n11911 & n11912;
  assign n15508 = n11862 & n11913;
  assign n15509 = (n11913 & n15476) | (n11913 & n15508) | (n15476 & n15508);
  assign n15510 = n11862 | n11913;
  assign n15511 = n15476 | n15510;
  assign n11916 = ~n15509 & n15511;
  assign n11923 = x79 & x107;
  assign n17579 = n11878 | n17567;
  assign n17580 = (n11827 & n17567) | (n11827 & n17579) | (n17567 & n17579);
  assign n15515 = n11923 & n17580;
  assign n17581 = n11923 & n17567;
  assign n17582 = (n11878 & n11923) | (n11878 & n17581) | (n11923 & n17581);
  assign n17583 = (n15455 & n15515) | (n15455 & n17582) | (n15515 & n17582);
  assign n17584 = (n11829 & n15515) | (n11829 & n17582) | (n15515 & n17582);
  assign n17585 = (n15419 & n17583) | (n15419 & n17584) | (n17583 & n17584);
  assign n15518 = n11923 | n17580;
  assign n17586 = n11923 | n17567;
  assign n17587 = n11878 | n17586;
  assign n17588 = (n15455 & n15518) | (n15455 & n17587) | (n15518 & n17587);
  assign n17589 = (n11829 & n15518) | (n11829 & n17587) | (n15518 & n17587);
  assign n17590 = (n15419 & n17588) | (n15419 & n17589) | (n17588 & n17589);
  assign n11926 = ~n17585 & n17590;
  assign n15521 = n11883 & n11926;
  assign n17591 = (n11926 & n15492) | (n11926 & n15521) | (n15492 & n15521);
  assign n17592 = (n11885 & n11926) | (n11885 & n15521) | (n11926 & n15521);
  assign n17593 = (n15460 & n17591) | (n15460 & n17592) | (n17591 & n17592);
  assign n15523 = n11883 | n11926;
  assign n17594 = n15492 | n15523;
  assign n17595 = n11885 | n15523;
  assign n17596 = (n15460 & n17594) | (n15460 & n17595) | (n17594 & n17595);
  assign n11929 = ~n17593 & n17596;
  assign n11930 = x78 & x108;
  assign n11931 = n11929 & n11930;
  assign n11932 = n11929 | n11930;
  assign n11933 = ~n11931 & n11932;
  assign n15525 = n11890 & n11933;
  assign n15526 = (n11933 & n15497) | (n11933 & n15525) | (n15497 & n15525);
  assign n15527 = n11890 | n11933;
  assign n15528 = n15497 | n15527;
  assign n11936 = ~n15526 & n15528;
  assign n11937 = x77 & x109;
  assign n11938 = n11936 & n11937;
  assign n11939 = n11936 | n11937;
  assign n11940 = ~n11938 & n11939;
  assign n15529 = n11897 & n11940;
  assign n15530 = (n11940 & n15501) | (n11940 & n15529) | (n15501 & n15529);
  assign n15531 = n11897 | n11940;
  assign n15532 = n15501 | n15531;
  assign n11943 = ~n15530 & n15532;
  assign n11944 = x76 & x110;
  assign n11945 = n11943 & n11944;
  assign n11946 = n11943 | n11944;
  assign n11947 = ~n11945 & n11946;
  assign n15533 = n11904 & n11947;
  assign n15534 = (n11947 & n15505) | (n11947 & n15533) | (n15505 & n15533);
  assign n15535 = n11904 | n11947;
  assign n15536 = n15505 | n15535;
  assign n11950 = ~n15534 & n15536;
  assign n11951 = x75 & x111;
  assign n11952 = n11950 & n11951;
  assign n11953 = n11950 | n11951;
  assign n11954 = ~n11952 & n11953;
  assign n15537 = n11911 & n11954;
  assign n15538 = (n11954 & n15509) | (n11954 & n15537) | (n15509 & n15537);
  assign n15539 = n11911 | n11954;
  assign n15540 = n15509 | n15539;
  assign n11957 = ~n15538 & n15540;
  assign n11963 = x79 & x108;
  assign n17597 = n11926 | n17585;
  assign n17598 = (n11883 & n17585) | (n11883 & n17597) | (n17585 & n17597);
  assign n15544 = n11963 & n17598;
  assign n17599 = n11963 & n17585;
  assign n17600 = (n11926 & n11963) | (n11926 & n17599) | (n11963 & n17599);
  assign n17601 = (n15492 & n15544) | (n15492 & n17600) | (n15544 & n17600);
  assign n17602 = (n11885 & n15544) | (n11885 & n17600) | (n15544 & n17600);
  assign n17603 = (n15460 & n17601) | (n15460 & n17602) | (n17601 & n17602);
  assign n15547 = n11963 | n17598;
  assign n17604 = n11963 | n17585;
  assign n17605 = n11926 | n17604;
  assign n17606 = (n15492 & n15547) | (n15492 & n17605) | (n15547 & n17605);
  assign n17607 = (n11885 & n15547) | (n11885 & n17605) | (n15547 & n17605);
  assign n17608 = (n15460 & n17606) | (n15460 & n17607) | (n17606 & n17607);
  assign n11966 = ~n17603 & n17608;
  assign n15550 = n11931 & n11966;
  assign n17609 = (n11966 & n15525) | (n11966 & n15550) | (n15525 & n15550);
  assign n17610 = (n11933 & n11966) | (n11933 & n15550) | (n11966 & n15550);
  assign n17611 = (n15497 & n17609) | (n15497 & n17610) | (n17609 & n17610);
  assign n15552 = n11931 | n11966;
  assign n17612 = n15525 | n15552;
  assign n17613 = n11933 | n15552;
  assign n17614 = (n15497 & n17612) | (n15497 & n17613) | (n17612 & n17613);
  assign n11969 = ~n17611 & n17614;
  assign n11970 = x78 & x109;
  assign n11971 = n11969 & n11970;
  assign n11972 = n11969 | n11970;
  assign n11973 = ~n11971 & n11972;
  assign n15554 = n11938 & n11973;
  assign n15555 = (n11973 & n15530) | (n11973 & n15554) | (n15530 & n15554);
  assign n15556 = n11938 | n11973;
  assign n15557 = n15530 | n15556;
  assign n11976 = ~n15555 & n15557;
  assign n11977 = x77 & x110;
  assign n11978 = n11976 & n11977;
  assign n11979 = n11976 | n11977;
  assign n11980 = ~n11978 & n11979;
  assign n15558 = n11945 & n11980;
  assign n15559 = (n11980 & n15534) | (n11980 & n15558) | (n15534 & n15558);
  assign n15560 = n11945 | n11980;
  assign n15561 = n15534 | n15560;
  assign n11983 = ~n15559 & n15561;
  assign n11984 = x76 & x111;
  assign n11985 = n11983 & n11984;
  assign n11986 = n11983 | n11984;
  assign n11987 = ~n11985 & n11986;
  assign n15562 = n11952 & n11987;
  assign n15563 = (n11987 & n15538) | (n11987 & n15562) | (n15538 & n15562);
  assign n15564 = n11952 | n11987;
  assign n15565 = n15538 | n15564;
  assign n11990 = ~n15563 & n15565;
  assign n11995 = x79 & x109;
  assign n17615 = n11966 | n17603;
  assign n17616 = (n11931 & n17603) | (n11931 & n17615) | (n17603 & n17615);
  assign n15569 = n11995 & n17616;
  assign n17617 = n11995 & n17603;
  assign n17618 = (n11966 & n11995) | (n11966 & n17617) | (n11995 & n17617);
  assign n17619 = (n15525 & n15569) | (n15525 & n17618) | (n15569 & n17618);
  assign n17620 = (n11933 & n15569) | (n11933 & n17618) | (n15569 & n17618);
  assign n17621 = (n15497 & n17619) | (n15497 & n17620) | (n17619 & n17620);
  assign n15572 = n11995 | n17616;
  assign n17622 = n11995 | n17603;
  assign n17623 = n11966 | n17622;
  assign n17624 = (n15525 & n15572) | (n15525 & n17623) | (n15572 & n17623);
  assign n17625 = (n11933 & n15572) | (n11933 & n17623) | (n15572 & n17623);
  assign n17626 = (n15497 & n17624) | (n15497 & n17625) | (n17624 & n17625);
  assign n11998 = ~n17621 & n17626;
  assign n15575 = n11971 & n11998;
  assign n17627 = (n11998 & n15554) | (n11998 & n15575) | (n15554 & n15575);
  assign n17628 = (n11973 & n11998) | (n11973 & n15575) | (n11998 & n15575);
  assign n17629 = (n15530 & n17627) | (n15530 & n17628) | (n17627 & n17628);
  assign n15577 = n11971 | n11998;
  assign n17630 = n15554 | n15577;
  assign n17631 = n11973 | n15577;
  assign n17632 = (n15530 & n17630) | (n15530 & n17631) | (n17630 & n17631);
  assign n12001 = ~n17629 & n17632;
  assign n12002 = x78 & x110;
  assign n12003 = n12001 & n12002;
  assign n12004 = n12001 | n12002;
  assign n12005 = ~n12003 & n12004;
  assign n15579 = n11978 & n12005;
  assign n15580 = (n12005 & n15559) | (n12005 & n15579) | (n15559 & n15579);
  assign n15581 = n11978 | n12005;
  assign n15582 = n15559 | n15581;
  assign n12008 = ~n15580 & n15582;
  assign n12009 = x77 & x111;
  assign n12010 = n12008 & n12009;
  assign n12011 = n12008 | n12009;
  assign n12012 = ~n12010 & n12011;
  assign n15583 = n11985 & n12012;
  assign n15584 = (n12012 & n15563) | (n12012 & n15583) | (n15563 & n15583);
  assign n15585 = n11985 | n12012;
  assign n15586 = n15563 | n15585;
  assign n12015 = ~n15584 & n15586;
  assign n12019 = x79 & x110;
  assign n17633 = n11998 | n17621;
  assign n17634 = (n11971 & n17621) | (n11971 & n17633) | (n17621 & n17633);
  assign n15590 = n12019 & n17634;
  assign n17635 = n12019 & n17621;
  assign n17636 = (n11998 & n12019) | (n11998 & n17635) | (n12019 & n17635);
  assign n17637 = (n15554 & n15590) | (n15554 & n17636) | (n15590 & n17636);
  assign n17638 = (n11973 & n15590) | (n11973 & n17636) | (n15590 & n17636);
  assign n17639 = (n15530 & n17637) | (n15530 & n17638) | (n17637 & n17638);
  assign n15593 = n12019 | n17634;
  assign n17640 = n12019 | n17621;
  assign n17641 = n11998 | n17640;
  assign n17642 = (n15554 & n15593) | (n15554 & n17641) | (n15593 & n17641);
  assign n17643 = (n11973 & n15593) | (n11973 & n17641) | (n15593 & n17641);
  assign n17644 = (n15530 & n17642) | (n15530 & n17643) | (n17642 & n17643);
  assign n12022 = ~n17639 & n17644;
  assign n15596 = n12003 & n12022;
  assign n17645 = (n12022 & n15579) | (n12022 & n15596) | (n15579 & n15596);
  assign n17646 = (n12005 & n12022) | (n12005 & n15596) | (n12022 & n15596);
  assign n17647 = (n15559 & n17645) | (n15559 & n17646) | (n17645 & n17646);
  assign n15598 = n12003 | n12022;
  assign n17648 = n15579 | n15598;
  assign n17649 = n12005 | n15598;
  assign n17650 = (n15559 & n17648) | (n15559 & n17649) | (n17648 & n17649);
  assign n12025 = ~n17647 & n17650;
  assign n12026 = x78 & x111;
  assign n12027 = n12025 & n12026;
  assign n12028 = n12025 | n12026;
  assign n12029 = ~n12027 & n12028;
  assign n15600 = n12010 & n12029;
  assign n15601 = (n12029 & n15584) | (n12029 & n15600) | (n15584 & n15600);
  assign n15602 = n12010 | n12029;
  assign n15603 = n15584 | n15602;
  assign n12032 = ~n15601 & n15603;
  assign n12035 = x79 & x111;
  assign n17651 = n12022 | n17639;
  assign n17652 = (n12003 & n17639) | (n12003 & n17651) | (n17639 & n17651);
  assign n15607 = n12035 & n17652;
  assign n17653 = n12035 & n17639;
  assign n17654 = (n12022 & n12035) | (n12022 & n17653) | (n12035 & n17653);
  assign n17655 = (n15579 & n15607) | (n15579 & n17654) | (n15607 & n17654);
  assign n17656 = (n12005 & n15607) | (n12005 & n17654) | (n15607 & n17654);
  assign n17657 = (n15559 & n17655) | (n15559 & n17656) | (n17655 & n17656);
  assign n15610 = n12035 | n17652;
  assign n17658 = n12035 | n17639;
  assign n17659 = n12022 | n17658;
  assign n17660 = (n15579 & n15610) | (n15579 & n17659) | (n15610 & n17659);
  assign n17661 = (n12005 & n15610) | (n12005 & n17659) | (n15610 & n17659);
  assign n17662 = (n15559 & n17660) | (n15559 & n17661) | (n17660 & n17661);
  assign n12038 = ~n17657 & n17662;
  assign n15613 = n12027 & n12038;
  assign n17663 = (n12038 & n15600) | (n12038 & n15613) | (n15600 & n15613);
  assign n17664 = (n12029 & n12038) | (n12029 & n15613) | (n12038 & n15613);
  assign n17665 = (n15584 & n17663) | (n15584 & n17664) | (n17663 & n17664);
  assign n15615 = n12027 | n12038;
  assign n17666 = n15600 | n15615;
  assign n17667 = n12029 | n15615;
  assign n17668 = (n15584 & n17666) | (n15584 & n17667) | (n17666 & n17667);
  assign n12041 = ~n17665 & n17668;
  assign n15618 = n12038 | n17657;
  assign n17669 = n12038 | n17657;
  assign n17670 = (n12027 & n17657) | (n12027 & n17669) | (n17657 & n17669);
  assign n17671 = (n15600 & n15618) | (n15600 & n17670) | (n15618 & n17670);
  assign n17672 = (n12029 & n15618) | (n12029 & n17670) | (n15618 & n17670);
  assign n17673 = (n15584 & n17671) | (n15584 & n17672) | (n17671 & n17672);
  assign n18337 = x112 & x144;
  assign n18338 = x113 & x144;
  assign n18339 = x112 & x145;
  assign n18340 = n18338 & n18339;
  assign n18341 = n18338 | n18339;
  assign n18342 = ~n18340 & n18341;
  assign n18343 = x114 & x144;
  assign n18344 = x113 & x145;
  assign n18345 = n18343 & ~n18344;
  assign n18346 = ~n18343 & n18344;
  assign n18347 = n18345 | n18346;
  assign n18348 = ~n18340 & n18347;
  assign n18349 = n18340 & ~n18347;
  assign n18350 = n18348 | n18349;
  assign n18351 = x112 & x146;
  assign n18352 = n18350 & n18351;
  assign n18353 = n18350 | n18351;
  assign n18354 = ~n18352 & n18353;
  assign n18355 = n18337 | n18343;
  assign n18356 = n18344 & n18355;
  assign n18357 = x115 & x144;
  assign n18358 = x114 & x145;
  assign n18359 = n18357 & n18358;
  assign n18360 = n18357 | n18358;
  assign n18361 = ~n18359 & n18360;
  assign n18362 = n18356 & n18361;
  assign n18363 = n18356 | n18361;
  assign n18364 = ~n18362 & n18363;
  assign n18365 = x113 & x146;
  assign n18366 = n18364 & n18365;
  assign n18367 = n18364 | n18365;
  assign n18368 = ~n18366 & n18367;
  assign n18369 = ~n18352 & n18368;
  assign n18370 = n18352 & ~n18368;
  assign n18371 = n18369 | n18370;
  assign n18372 = x112 & x147;
  assign n18373 = n18371 & n18372;
  assign n18374 = n18371 | n18372;
  assign n18375 = ~n18373 & n18374;
  assign n18376 = n18352 | n18366;
  assign n18377 = n18367 & n18376;
  assign n18378 = n18356 | n18359;
  assign n18379 = x116 & x144;
  assign n18380 = x115 & x145;
  assign n18381 = n18379 | n18380;
  assign n18382 = n18379 & n18380;
  assign n18383 = n18381 & ~n18382;
  assign n18384 = n18360 & n18383;
  assign n18385 = n18378 & n18384;
  assign n18386 = n18359 | n18383;
  assign n18387 = n18362 | n18386;
  assign n18388 = ~n18385 & n18387;
  assign n18389 = x114 & x146;
  assign n18390 = n18388 & n18389;
  assign n18391 = n18388 | n18389;
  assign n18392 = ~n18390 & n18391;
  assign n18393 = n18377 & n18392;
  assign n18394 = n18377 | n18392;
  assign n18395 = ~n18393 & n18394;
  assign n18396 = x113 & x147;
  assign n18397 = n18395 | n18396;
  assign n18398 = n18395 & n18396;
  assign n18399 = n18397 & ~n18398;
  assign n18400 = ~n18373 & n18399;
  assign n18401 = n18373 & ~n18399;
  assign n18402 = n18400 | n18401;
  assign n18403 = x112 & x148;
  assign n18404 = n18402 & n18403;
  assign n18405 = n18402 | n18403;
  assign n18406 = ~n18404 & n18405;
  assign n18407 = n18373 | n18398;
  assign n18408 = n18397 & n18407;
  assign n18409 = n18390 | n18393;
  assign n18410 = n18382 | n18385;
  assign n18411 = x117 & x144;
  assign n18412 = x116 & x145;
  assign n18413 = n18411 & n18412;
  assign n18414 = n18411 | n18412;
  assign n18415 = ~n18413 & n18414;
  assign n18416 = x115 & x146;
  assign n18417 = n18415 & n18416;
  assign n18418 = n18415 | n18416;
  assign n18419 = ~n18417 & n18418;
  assign n18420 = ~n18410 & n18419;
  assign n18421 = n18410 & ~n18419;
  assign n18422 = n18420 | n18421;
  assign n18423 = x114 & x147;
  assign n18424 = n18422 & n18423;
  assign n18425 = n18422 | n18423;
  assign n18426 = ~n18424 & n18425;
  assign n18427 = n18409 | n18426;
  assign n18428 = n18409 & n18426;
  assign n18429 = n18427 & ~n18428;
  assign n18430 = n18408 & n18429;
  assign n18431 = n18408 | n18429;
  assign n18432 = ~n18430 & n18431;
  assign n18433 = x113 & x148;
  assign n18434 = n18432 | n18433;
  assign n18435 = n18432 & n18433;
  assign n18436 = n18434 & ~n18435;
  assign n18437 = ~n18404 & n18436;
  assign n18438 = n18404 & ~n18436;
  assign n18439 = n18437 | n18438;
  assign n18440 = x112 & x149;
  assign n18441 = n18439 & n18440;
  assign n18442 = n18439 | n18440;
  assign n18443 = ~n18441 & n18442;
  assign n18444 = x114 & x148;
  assign n29529 = n18390 | n18422;
  assign n29530 = n18393 | n29529;
  assign n18446 = n18377 | n18390;
  assign n18447 = n18391 & n18422;
  assign n18448 = n18446 & n18447;
  assign n18449 = n18423 & ~n18448;
  assign n18450 = n29530 & n18449;
  assign n29531 = n18429 | n18450;
  assign n29532 = (n18408 & n18450) | (n18408 & n29531) | (n18450 & n29531);
  assign n29533 = n18382 & n18415;
  assign n29534 = (n18385 & n18415) | (n18385 & n29533) | (n18415 & n29533);
  assign n34721 = n18382 & n18416;
  assign n34722 = (n18415 & n18416) | (n18415 & n34721) | (n18416 & n34721);
  assign n29538 = (n18385 & n18416) | (n18385 & n34722) | (n18416 & n34722);
  assign n18455 = ~n29534 & n29538;
  assign n18457 = x118 & x144;
  assign n18458 = x117 & x145;
  assign n18459 = n18457 | n18458;
  assign n18460 = n18457 & n18458;
  assign n18461 = n18459 & ~n18460;
  assign n18462 = n18413 | n18461;
  assign n29539 = n18462 | n29533;
  assign n29540 = n18415 | n18462;
  assign n29541 = (n18385 & n29539) | (n18385 & n29540) | (n29539 & n29540);
  assign n18466 = n18414 & n18461;
  assign n18464 = n18382 | n18413;
  assign n29542 = n18464 & n18466;
  assign n29543 = (n18385 & n18466) | (n18385 & n29542) | (n18466 & n29542);
  assign n18468 = n29541 & ~n29543;
  assign n18469 = x116 & x146;
  assign n18470 = n18468 | n18469;
  assign n18471 = n18468 & n18469;
  assign n18472 = n18470 & ~n18471;
  assign n29544 = n18455 | n18472;
  assign n29545 = n18448 | n29544;
  assign n29546 = n18455 & n18472;
  assign n29547 = (n18448 & n18472) | (n18448 & n29546) | (n18472 & n29546);
  assign n18475 = n29545 & ~n29547;
  assign n18476 = x115 & x147;
  assign n18477 = n18475 & n18476;
  assign n18478 = n18475 | n18476;
  assign n18479 = ~n18477 & n18478;
  assign n18480 = n29532 & n18479;
  assign n18481 = n29532 | n18479;
  assign n18482 = ~n18480 & n18481;
  assign n18483 = n18444 | n18482;
  assign n18484 = n18444 & n18482;
  assign n18485 = n18483 & ~n18484;
  assign n18486 = n18404 | n18435;
  assign n18487 = n18434 & n18486;
  assign n18488 = n18485 & ~n18487;
  assign n18489 = ~n18485 & n18487;
  assign n18490 = n18488 | n18489;
  assign n18491 = x113 & x149;
  assign n18492 = n18490 | n18491;
  assign n18493 = n18490 & n18491;
  assign n18494 = n18492 & ~n18493;
  assign n18495 = ~n18441 & n18494;
  assign n18496 = n18441 & ~n18494;
  assign n18497 = n18495 | n18496;
  assign n18498 = x112 & x150;
  assign n18499 = n18497 & n18498;
  assign n18500 = n18497 | n18498;
  assign n18501 = ~n18499 & n18500;
  assign n18502 = n18441 | n18493;
  assign n18503 = n18492 & n18502;
  assign n29548 = n18483 & n18484;
  assign n29549 = (n18483 & n18487) | (n18483 & n29548) | (n18487 & n29548);
  assign n18506 = n18477 | n18480;
  assign n18509 = x119 & x144;
  assign n18510 = x118 & x145;
  assign n18511 = n18509 & n18510;
  assign n18512 = n18509 | n18510;
  assign n18513 = ~n18511 & n18512;
  assign n18514 = x117 & x146;
  assign n18515 = n18513 & n18514;
  assign n18516 = n18513 | n18514;
  assign n18517 = ~n18515 & n18516;
  assign n29550 = ~n18460 & n18517;
  assign n29551 = ~n29543 & n29550;
  assign n29552 = n18460 & ~n18517;
  assign n29553 = (~n18517 & n29543) | (~n18517 & n29552) | (n29543 & n29552);
  assign n18520 = n29551 | n29553;
  assign n18521 = x116 & x147;
  assign n18522 = n18520 & n18521;
  assign n18523 = n18520 | n18521;
  assign n18524 = ~n18522 & n18523;
  assign n29554 = n18471 | n18524;
  assign n29555 = n29547 | n29554;
  assign n29556 = n18471 & n18524;
  assign n29557 = (n18524 & n29547) | (n18524 & n29556) | (n29547 & n29556);
  assign n18527 = n29555 & ~n29557;
  assign n18528 = x115 & x148;
  assign n18529 = n18527 | n18528;
  assign n18530 = n18527 & n18528;
  assign n18531 = n18529 & ~n18530;
  assign n18532 = n18506 | n18531;
  assign n18533 = n18506 & n18531;
  assign n18534 = n18532 & ~n18533;
  assign n18535 = n29549 & n18534;
  assign n18536 = n29549 | n18534;
  assign n18537 = ~n18535 & n18536;
  assign n18538 = x114 & x149;
  assign n18539 = n18537 & n18538;
  assign n18540 = n18537 | n18538;
  assign n18541 = ~n18539 & n18540;
  assign n18542 = n18503 & n18541;
  assign n18543 = n18503 | n18541;
  assign n18544 = ~n18542 & n18543;
  assign n18545 = x113 & x150;
  assign n18546 = n18544 | n18545;
  assign n18547 = n18544 & n18545;
  assign n18548 = n18546 & ~n18547;
  assign n18549 = ~n18499 & n18548;
  assign n18550 = n18499 & ~n18548;
  assign n18551 = n18549 | n18550;
  assign n18552 = x112 & x151;
  assign n18553 = n18551 & n18552;
  assign n18554 = n18551 | n18552;
  assign n18555 = ~n18553 & n18554;
  assign n18556 = x113 & x151;
  assign n18557 = n18499 | n18547;
  assign n18558 = n18546 & n18557;
  assign n29558 = n18477 | n18527;
  assign n29559 = n18480 | n29558;
  assign n18560 = n29532 | n18477;
  assign n18561 = n18478 & n18527;
  assign n29560 = n18528 & ~n18561;
  assign n29561 = (n18528 & ~n18560) | (n18528 & n29560) | (~n18560 & n29560);
  assign n18564 = n29559 & n29561;
  assign n29562 = n18534 | n18564;
  assign n29563 = (n18564 & n29549) | (n18564 & n29562) | (n29549 & n29562);
  assign n29564 = n18471 | n18520;
  assign n29565 = n29547 | n29564;
  assign n18568 = n18470 & n18520;
  assign n29566 = n18455 | n18471;
  assign n29568 = n18568 & n29566;
  assign n29569 = (n18448 & n18568) | (n18448 & n29568) | (n18568 & n29568);
  assign n18570 = n18521 & ~n29569;
  assign n18571 = n29565 & n18570;
  assign n29570 = n18561 | n18571;
  assign n29571 = (n18560 & n18571) | (n18560 & n29570) | (n18571 & n29570);
  assign n29572 = n18460 & n18513;
  assign n29573 = (n18513 & n29543) | (n18513 & n29572) | (n29543 & n29572);
  assign n34723 = n18460 & n18514;
  assign n34724 = (n18513 & n18514) | (n18513 & n34723) | (n18514 & n34723);
  assign n29577 = (n18514 & n29543) | (n18514 & n34724) | (n29543 & n34724);
  assign n18576 = ~n29573 & n29577;
  assign n18578 = x120 & x144;
  assign n18579 = x119 & x145;
  assign n18580 = n18578 | n18579;
  assign n18581 = n18578 & n18579;
  assign n18582 = n18580 & ~n18581;
  assign n18583 = n18511 | n18582;
  assign n29578 = n18583 | n29572;
  assign n29579 = n18513 | n18583;
  assign n29580 = (n29543 & n29578) | (n29543 & n29579) | (n29578 & n29579);
  assign n18585 = n18512 & n18582;
  assign n29581 = n18460 | n18511;
  assign n29583 = n18585 & n29581;
  assign n29584 = (n18585 & n29543) | (n18585 & n29583) | (n29543 & n29583);
  assign n18588 = n29580 & ~n29584;
  assign n18589 = x118 & x146;
  assign n18590 = n18588 | n18589;
  assign n18591 = n18588 & n18589;
  assign n18592 = n18590 & ~n18591;
  assign n29585 = ~n18576 & n18592;
  assign n29586 = ~n29569 & n29585;
  assign n29587 = n18576 & ~n18592;
  assign n29588 = (~n18592 & n29569) | (~n18592 & n29587) | (n29569 & n29587);
  assign n18595 = n29586 | n29588;
  assign n18596 = x117 & x147;
  assign n18597 = x116 & x148;
  assign n18598 = n18596 | n18597;
  assign n18599 = n18596 & n18597;
  assign n18600 = n18598 & ~n18599;
  assign n18601 = n18595 | n18600;
  assign n18602 = n18595 & n18600;
  assign n18603 = n18601 & ~n18602;
  assign n18604 = n29571 | n18603;
  assign n18605 = n29571 & n18603;
  assign n18606 = n18604 & ~n18605;
  assign n18607 = n29563 & n18606;
  assign n18608 = n18564 | n18606;
  assign n18609 = n18535 | n18608;
  assign n18610 = ~n18607 & n18609;
  assign n18611 = x115 & x149;
  assign n18612 = n18610 | n18611;
  assign n34725 = n18564 & n18611;
  assign n34726 = (n18606 & n18611) | (n18606 & n34725) | (n18611 & n34725);
  assign n29590 = (n18535 & n18611) | (n18535 & n34726) | (n18611 & n34726);
  assign n18614 = ~n18607 & n29590;
  assign n18615 = n18612 & ~n18614;
  assign n18616 = n18539 | n18542;
  assign n18617 = n18615 & ~n18616;
  assign n18618 = ~n18615 & n18616;
  assign n18619 = n18617 | n18618;
  assign n18620 = x114 & x150;
  assign n18621 = n18619 | n18620;
  assign n18622 = n18619 & n18620;
  assign n18623 = n18621 & ~n18622;
  assign n18624 = ~n18558 & n18623;
  assign n18625 = n18558 & ~n18623;
  assign n18626 = n18624 | n18625;
  assign n18627 = n18556 & ~n18626;
  assign n18628 = ~n18556 & n18626;
  assign n18629 = n18627 | n18628;
  assign n18630 = ~n18553 & n18629;
  assign n18631 = n18553 & ~n18629;
  assign n18632 = n18630 | n18631;
  assign n18633 = x112 & x152;
  assign n18634 = n18632 & n18633;
  assign n18635 = n18632 | n18633;
  assign n18636 = ~n18634 & n18635;
  assign n18637 = n18539 | n18614;
  assign n29591 = n18612 & n18637;
  assign n29592 = (n18542 & n18612) | (n18542 & n29591) | (n18612 & n29591);
  assign n18640 = n18595 & n18596;
  assign n18641 = n18595 | n18596;
  assign n18642 = ~n18640 & n18641;
  assign n18643 = n29571 | n18642;
  assign n29593 = n18597 & ~n18642;
  assign n29594 = (n18597 & ~n29571) | (n18597 & n29593) | (~n29571 & n29593);
  assign n18646 = n18643 & n29594;
  assign n29595 = n18606 | n18646;
  assign n29596 = (n18646 & n29563) | (n18646 & n29595) | (n29563 & n29595);
  assign n29597 = n18640 | n18642;
  assign n29598 = (n18640 & n29571) | (n18640 & n29597) | (n29571 & n29597);
  assign n29599 = n18576 & n18590;
  assign n29600 = (n18590 & n29569) | (n18590 & n29599) | (n29569 & n29599);
  assign n18650 = x119 & x146;
  assign n18656 = x121 & x144;
  assign n18657 = x120 & x145;
  assign n18658 = n18656 & n18657;
  assign n18659 = n18656 | n18657;
  assign n18660 = ~n18658 & n18659;
  assign n18651 = n18458 | n18579;
  assign n18652 = n18457 & n18651;
  assign n34727 = n18581 | n18652;
  assign n34728 = (n18581 & n18585) | (n18581 & n34727) | (n18585 & n34727);
  assign n34731 = n18660 & n34728;
  assign n34729 = n18512 | n18581;
  assign n34730 = (n18581 & n18582) | (n18581 & n34729) | (n18582 & n34729);
  assign n34732 = n18660 & n34730;
  assign n34733 = (n29543 & n34731) | (n29543 & n34732) | (n34731 & n34732);
  assign n34734 = n18660 | n34728;
  assign n34735 = n18660 | n34730;
  assign n34736 = (n29543 & n34734) | (n29543 & n34735) | (n34734 & n34735);
  assign n18663 = ~n34733 & n34736;
  assign n18664 = n18650 & n18663;
  assign n18665 = n18650 | n18663;
  assign n18666 = ~n18664 & n18665;
  assign n18667 = n18591 | n18666;
  assign n18668 = n29600 | n18667;
  assign n29606 = n18576 | n18591;
  assign n29607 = n29569 | n29606;
  assign n18670 = n18590 & n18666;
  assign n18671 = n29607 & n18670;
  assign n18672 = n18668 & ~n18671;
  assign n18673 = x118 & x147;
  assign n18674 = n18672 & n18673;
  assign n18675 = n18672 | n18673;
  assign n18676 = ~n18674 & n18675;
  assign n18677 = x117 & x148;
  assign n18678 = n18676 & n18677;
  assign n18679 = n18676 | n18677;
  assign n18680 = ~n18678 & n18679;
  assign n18681 = n29598 | n18680;
  assign n18682 = n29598 & n18680;
  assign n18683 = n18681 & ~n18682;
  assign n18684 = x116 & x149;
  assign n18685 = n18683 | n18684;
  assign n18686 = n18683 & n18684;
  assign n18687 = n18685 & ~n18686;
  assign n18688 = ~n29596 & n18687;
  assign n18689 = n29596 & ~n18687;
  assign n18690 = n18688 | n18689;
  assign n18691 = n29592 & ~n18690;
  assign n18692 = ~n29592 & n18690;
  assign n18693 = n18691 | n18692;
  assign n18694 = x115 & x150;
  assign n18695 = n18693 | n18694;
  assign n18696 = n18693 & n18694;
  assign n18697 = n18695 & ~n18696;
  assign n18698 = n18558 | n18622;
  assign n18699 = n18621 & n18698;
  assign n18700 = n18697 & ~n18699;
  assign n18701 = ~n18697 & n18699;
  assign n18702 = n18700 | n18701;
  assign n18703 = x114 & x151;
  assign n18704 = n18702 | n18703;
  assign n18705 = n18702 & n18703;
  assign n18706 = n18704 & ~n18705;
  assign n29608 = n18633 & n18706;
  assign n29609 = n18632 & n29608;
  assign n29610 = n18633 | n18706;
  assign n29611 = (n18632 & n18706) | (n18632 & n29610) | (n18706 & n29610);
  assign n18709 = ~n29609 & n29611;
  assign n29614 = n18552 | n18556;
  assign n29615 = (n18551 & n18556) | (n18551 & n29614) | (n18556 & n29614);
  assign n29612 = n18552 & n18556;
  assign n29613 = n18551 & n29612;
  assign n29616 = n29613 & n29615;
  assign n29617 = (n18626 & n29615) | (n18626 & n29616) | (n29615 & n29616);
  assign n18714 = x113 & x152;
  assign n18715 = n29617 & ~n18714;
  assign n18716 = ~n29617 & n18714;
  assign n18717 = n18715 | n18716;
  assign n18718 = ~n18709 & n18717;
  assign n18719 = n18709 & ~n18717;
  assign n18720 = n18718 | n18719;
  assign n18721 = x112 & x153;
  assign n18722 = n18720 & n18721;
  assign n18723 = n18720 | n18721;
  assign n18724 = ~n18722 & n18723;
  assign n18728 = n29596 & n18683;
  assign n29620 = (n18684 & n18686) | (n18684 & n29596) | (n18686 & n29596);
  assign n18731 = ~n18728 & n29620;
  assign n29621 = n18690 | n18731;
  assign n29622 = (n18731 & n29592) | (n18731 & n29621) | (n29592 & n29621);
  assign n18733 = n29598 | n18676;
  assign n18734 = n29571 | n18640;
  assign n18735 = n18641 & n18676;
  assign n18736 = n18734 & n18735;
  assign n18737 = n18677 & ~n18736;
  assign n18738 = n18733 & n18737;
  assign n29623 = n18683 | n18738;
  assign n29624 = (n18738 & n29596) | (n18738 & n29623) | (n29596 & n29623);
  assign n37285 = n18590 | n18664;
  assign n37286 = (n18664 & n18666) | (n18664 & n37285) | (n18666 & n37285);
  assign n34738 = (n18664 & n29607) | (n18664 & n37286) | (n29607 & n37286);
  assign n18743 = x122 & x144;
  assign n18744 = x121 & x145;
  assign n18745 = n18743 | n18744;
  assign n18746 = n18743 & n18744;
  assign n18747 = n18745 & ~n18746;
  assign n18748 = n18659 & n18747;
  assign n34739 = n18658 & n18659;
  assign n34740 = n18747 & n34739;
  assign n34741 = (n18748 & n34728) | (n18748 & n34740) | (n34728 & n34740);
  assign n34742 = (n18748 & n34730) | (n18748 & n34740) | (n34730 & n34740);
  assign n34743 = (n29543 & n34741) | (n29543 & n34742) | (n34741 & n34742);
  assign n18750 = n18658 | n18747;
  assign n29627 = n18660 | n18750;
  assign n34744 = (n18750 & n29627) | (n18750 & n34728) | (n29627 & n34728);
  assign n34745 = (n18750 & n29627) | (n18750 & n34730) | (n29627 & n34730);
  assign n34746 = (n29543 & n34744) | (n29543 & n34745) | (n34744 & n34745);
  assign n18752 = ~n34743 & n34746;
  assign n18753 = x120 & x146;
  assign n18754 = x119 & x147;
  assign n18755 = ~n18753 & n18754;
  assign n18756 = n18753 & ~n18754;
  assign n18757 = n18755 | n18756;
  assign n18758 = n18752 & ~n18757;
  assign n18759 = ~n18752 & n18757;
  assign n18760 = n18758 | n18759;
  assign n18761 = x118 & x148;
  assign n18762 = ~n18760 & n18761;
  assign n18763 = n18760 & ~n18761;
  assign n18764 = n18762 | n18763;
  assign n18765 = n34738 | n18764;
  assign n18766 = n34738 & n18764;
  assign n18767 = n18765 & ~n18766;
  assign n18768 = x117 & x149;
  assign n18769 = n18767 & ~n18768;
  assign n18770 = ~n18767 & n18768;
  assign n18771 = n18769 | n18770;
  assign n34747 = n18674 | n18771;
  assign n34748 = n18736 | n34747;
  assign n34749 = n18674 & n18771;
  assign n34750 = (n18736 & n18771) | (n18736 & n34749) | (n18771 & n34749);
  assign n18774 = n34748 & ~n34750;
  assign n18775 = x116 & x150;
  assign n18776 = n18774 & ~n18775;
  assign n18777 = ~n18774 & n18775;
  assign n18778 = n18776 | n18777;
  assign n18779 = n29624 | n18778;
  assign n18780 = n29624 & n18778;
  assign n18781 = n18779 & ~n18780;
  assign n18782 = n29622 | n18781;
  assign n18783 = n29622 & n18781;
  assign n18784 = n18782 & ~n18783;
  assign n29618 = n18621 | n18696;
  assign n29619 = (n18696 & n18698) | (n18696 & n29618) | (n18698 & n29618);
  assign n29629 = n18695 | n18784;
  assign n29630 = (n18784 & n29619) | (n18784 & n29629) | (n29619 & n29629);
  assign n18786 = n18695 & n18784;
  assign n18787 = n29619 & n18786;
  assign n18788 = n29630 & ~n18787;
  assign n18789 = x115 & x151;
  assign n18790 = n18788 & ~n18789;
  assign n18791 = ~n18788 & n18789;
  assign n18792 = n18790 | n18791;
  assign n18793 = n18705 | n29617;
  assign n18794 = n18704 & n18793;
  assign n18795 = n18792 & ~n18794;
  assign n18796 = ~n18792 & n18794;
  assign n18797 = n18795 | n18796;
  assign n18798 = x114 & x152;
  assign n18799 = n18797 | n18798;
  assign n18800 = n18797 & n18798;
  assign n18801 = n18799 & ~n18800;
  assign n29631 = n18633 & n18714;
  assign n29632 = n18632 & n29631;
  assign n18803 = n18706 & ~n29617;
  assign n18804 = ~n18706 & n29617;
  assign n18805 = n18803 | n18804;
  assign n18806 = n29632 | n18805;
  assign n29633 = n18633 | n18714;
  assign n29634 = (n18632 & n18714) | (n18632 & n29633) | (n18714 & n29633);
  assign n18808 = n18806 & n29634;
  assign n18809 = n18801 & n18808;
  assign n18810 = n18801 | n18808;
  assign n18811 = ~n18809 & n18810;
  assign n18812 = x113 & x153;
  assign n18813 = n18811 | n18812;
  assign n18814 = n18811 & n18812;
  assign n18815 = n18813 & ~n18814;
  assign n18816 = n18722 & ~n18815;
  assign n18817 = ~n18722 & n18815;
  assign n18818 = n18816 | n18817;
  assign n18819 = x112 & x154;
  assign n18820 = n18818 & n18819;
  assign n18821 = n18818 | n18819;
  assign n18822 = ~n18820 & n18821;
  assign n18823 = x115 & x152;
  assign n18824 = n18788 | n18789;
  assign n18825 = n18788 & n18789;
  assign n29635 = n18704 | n18825;
  assign n29636 = (n18793 & n18825) | (n18793 & n29635) | (n18825 & n29635);
  assign n18827 = n18824 & n29636;
  assign n18828 = x116 & x151;
  assign n29641 = n18664 | n18760;
  assign n34751 = n18670 | n29641;
  assign n34752 = (n29607 & n29641) | (n29607 & n34751) | (n29641 & n34751);
  assign n29643 = n18664 & n18760;
  assign n34753 = (n18670 & n18760) | (n18670 & n29643) | (n18760 & n29643);
  assign n34754 = n18760 & n29643;
  assign n34755 = (n29607 & n34753) | (n29607 & n34754) | (n34753 & n34754);
  assign n18835 = n34752 & ~n34755;
  assign n29645 = n18674 & n18835;
  assign n29646 = (n18736 & n18835) | (n18736 & n29645) | (n18835 & n29645);
  assign n34756 = n18761 & n18835;
  assign n34757 = (n18674 & n18761) | (n18674 & n34756) | (n18761 & n34756);
  assign n29650 = (n18736 & n18761) | (n18736 & n34757) | (n18761 & n34757);
  assign n18839 = ~n29646 & n29650;
  assign n29637 = n18674 | n18767;
  assign n29638 = n18736 | n29637;
  assign n29639 = n18674 & n18767;
  assign n29640 = (n18736 & n18767) | (n18736 & n29639) | (n18767 & n29639);
  assign n18831 = n29638 & ~n29640;
  assign n29651 = n18831 | n18839;
  assign n29652 = (n18839 & n29624) | (n18839 & n29651) | (n29624 & n29651);
  assign n18841 = n18752 & n18753;
  assign n18845 = x121 & x146;
  assign n18847 = x123 & x144;
  assign n18848 = x122 & x145;
  assign n18849 = n18847 & n18848;
  assign n18850 = n18847 | n18848;
  assign n18851 = ~n18849 & n18850;
  assign n34760 = n18659 | n18746;
  assign n34761 = (n18746 & n18747) | (n18746 & n34760) | (n18747 & n34760);
  assign n29659 = n18851 & n34761;
  assign n34758 = n18746 & n18851;
  assign n34759 = (n18851 & n34740) | (n18851 & n34758) | (n34740 & n34758);
  assign n34762 = (n29659 & n34728) | (n29659 & n34759) | (n34728 & n34759);
  assign n34763 = (n29659 & n34730) | (n29659 & n34759) | (n34730 & n34759);
  assign n34764 = (n29543 & n34762) | (n29543 & n34763) | (n34762 & n34763);
  assign n29662 = n18851 | n34761;
  assign n34765 = n18746 | n18851;
  assign n34766 = n34740 | n34765;
  assign n34767 = (n29662 & n34728) | (n29662 & n34766) | (n34728 & n34766);
  assign n34768 = (n29662 & n34730) | (n29662 & n34766) | (n34730 & n34766);
  assign n34769 = (n29543 & n34767) | (n29543 & n34768) | (n34767 & n34768);
  assign n18854 = ~n34764 & n34769;
  assign n18855 = n18845 | n18854;
  assign n18856 = n18845 & n18854;
  assign n18857 = n18855 & ~n18856;
  assign n18858 = ~n18841 & n18857;
  assign n18842 = n18752 | n18753;
  assign n18843 = ~n18841 & n18842;
  assign n29653 = n18664 & n18843;
  assign n29664 = n18858 & ~n29653;
  assign n29665 = ~n18843 & n18858;
  assign n29666 = (~n18671 & n29664) | (~n18671 & n29665) | (n29664 & n29665);
  assign n18861 = n18842 & ~n18857;
  assign n29667 = n18664 | n18841;
  assign n29669 = n18861 & n29667;
  assign n29670 = (n18671 & n18861) | (n18671 & n29669) | (n18861 & n29669);
  assign n18863 = n29666 | n29670;
  assign n18864 = x120 & x147;
  assign n18865 = n18863 | n18864;
  assign n18866 = n18863 & n18864;
  assign n18867 = n18865 & ~n18866;
  assign n18868 = x119 & x148;
  assign n18869 = n18867 & n18868;
  assign n18870 = n18867 | n18868;
  assign n18871 = ~n18869 & n18870;
  assign n34770 = (n18670 & n18843) | (n18670 & n29653) | (n18843 & n29653);
  assign n34771 = n18843 & n29653;
  assign n34772 = (n29607 & n34770) | (n29607 & n34771) | (n34770 & n34771);
  assign n29671 = n18664 | n18843;
  assign n34773 = n18670 | n29671;
  assign n34774 = (n29607 & n29671) | (n29607 & n34773) | (n29671 & n34773);
  assign n18873 = ~n34772 & n34774;
  assign n18874 = n18754 & n18873;
  assign n29673 = n18874 | n29645;
  assign n29674 = n18835 | n18874;
  assign n29675 = (n18736 & n29673) | (n18736 & n29674) | (n29673 & n29674);
  assign n18876 = n18871 | n29675;
  assign n18877 = n18871 & n29675;
  assign n18878 = n18876 & ~n18877;
  assign n18879 = x118 & x149;
  assign n18880 = n18878 | n18879;
  assign n18881 = n18878 & n18879;
  assign n18882 = n18880 & ~n18881;
  assign n18883 = n29652 | n18882;
  assign n18884 = n29652 & n18882;
  assign n18885 = n18883 & ~n18884;
  assign n18886 = x117 & x150;
  assign n18887 = n18885 | n18886;
  assign n18888 = n18885 & n18886;
  assign n18889 = n18887 & ~n18888;
  assign n18894 = n29624 | n18831;
  assign n29676 = n18768 & ~n18831;
  assign n29677 = (n18768 & ~n29624) | (n18768 & n29676) | (~n29624 & n29676);
  assign n18896 = n18894 & n29677;
  assign n18890 = n29624 | n18774;
  assign n18891 = n29624 & n18774;
  assign n18892 = n18890 & ~n18891;
  assign n29678 = n18892 | n18896;
  assign n29679 = (n18896 & n29622) | (n18896 & n29678) | (n29622 & n29678);
  assign n18898 = n18889 | n29679;
  assign n18899 = n18889 & n29679;
  assign n18900 = n18898 & ~n18899;
  assign n18901 = n29622 | n18892;
  assign n29680 = n18775 & ~n18892;
  assign n29681 = (n18775 & ~n29622) | (n18775 & n29680) | (~n29622 & n29680);
  assign n18903 = n18901 & n29681;
  assign n29682 = n18786 | n18903;
  assign n29683 = (n18903 & n29619) | (n18903 & n29682) | (n29619 & n29682);
  assign n18905 = n18900 | n29683;
  assign n18906 = n18900 & n29683;
  assign n18907 = n18905 & ~n18906;
  assign n18908 = n18828 & n18907;
  assign n18909 = n18828 | n18907;
  assign n18910 = ~n18908 & n18909;
  assign n18911 = n18827 & n18910;
  assign n18912 = n18827 | n18910;
  assign n18913 = ~n18911 & n18912;
  assign n18914 = n18823 | n18913;
  assign n18915 = n18823 & n18913;
  assign n18916 = n18914 & ~n18915;
  assign n18917 = n18800 | n18808;
  assign n18918 = n18799 & n18917;
  assign n18919 = n18916 & ~n18918;
  assign n18920 = ~n18916 & n18918;
  assign n18921 = n18919 | n18920;
  assign n18922 = x114 & x153;
  assign n18923 = n18921 | n18922;
  assign n18924 = n18921 & n18922;
  assign n18925 = n18923 & ~n18924;
  assign n29686 = n18721 & n18812;
  assign n29687 = n18720 & n29686;
  assign n29684 = n18721 | n18812;
  assign n29685 = (n18720 & n18812) | (n18720 & n29684) | (n18812 & n29684);
  assign n29688 = n29685 | n29687;
  assign n29689 = (n18811 & n29687) | (n18811 & n29688) | (n29687 & n29688);
  assign n18930 = n18925 & ~n29689;
  assign n18931 = ~n18925 & n29689;
  assign n18932 = n18930 | n18931;
  assign n18933 = x113 & x154;
  assign n18934 = n18932 & n18933;
  assign n18935 = n18932 | n18933;
  assign n18936 = ~n18934 & n18935;
  assign n18937 = ~n18820 & n18936;
  assign n18938 = n18820 & ~n18936;
  assign n18939 = n18937 | n18938;
  assign n18940 = x112 & x155;
  assign n18941 = n18939 & n18940;
  assign n18942 = n18939 | n18940;
  assign n18943 = ~n18941 & n18942;
  assign n18944 = n18924 | n29689;
  assign n18946 = x114 & x154;
  assign n34775 = n18922 & n18946;
  assign n34776 = (n18921 & n18946) | (n18921 & n34775) | (n18946 & n34775);
  assign n29691 = n18944 & n34776;
  assign n34777 = n18922 | n18946;
  assign n34778 = n18921 | n34777;
  assign n29693 = (n18944 & n18946) | (n18944 & n34778) | (n18946 & n34778);
  assign n18949 = ~n29691 & n29693;
  assign n18950 = x116 & x152;
  assign n29694 = n18908 | n18910;
  assign n29695 = (n18827 & n18908) | (n18827 & n29694) | (n18908 & n29694);
  assign n18952 = x117 & x151;
  assign n29696 = n18878 & n29651;
  assign n29697 = n18839 & n18878;
  assign n29698 = (n29624 & n29696) | (n29624 & n29697) | (n29696 & n29697);
  assign n29699 = n18867 | n29674;
  assign n29700 = n18867 | n29673;
  assign n29701 = (n18736 & n29699) | (n18736 & n29700) | (n29699 & n29700);
  assign n29702 = n18867 & n29674;
  assign n29703 = n18867 & n29673;
  assign n29704 = (n18736 & n29702) | (n18736 & n29703) | (n29702 & n29703);
  assign n18956 = n18868 & ~n29704;
  assign n18957 = n29701 & n18956;
  assign n18958 = n29698 | n18957;
  assign n18962 = x122 & x146;
  assign n18964 = x124 & x144;
  assign n18965 = x123 & x145;
  assign n18966 = n18964 & ~n18965;
  assign n18967 = ~n18964 & n18965;
  assign n18968 = n18966 | n18967;
  assign n29707 = n18849 & n18968;
  assign n29708 = (n18968 & n34764) | (n18968 & n29707) | (n34764 & n29707);
  assign n29709 = n18849 | n18968;
  assign n29710 = n34764 | n29709;
  assign n18971 = ~n29708 & n29710;
  assign n18972 = n18962 & n18971;
  assign n18973 = n18962 | n18971;
  assign n18974 = ~n18972 & n18973;
  assign n18959 = n18842 & n18857;
  assign n29705 = n18959 & n29667;
  assign n29711 = n18856 & n18974;
  assign n34779 = (n18974 & n29705) | (n18974 & n29711) | (n29705 & n29711);
  assign n34780 = (n18959 & n18974) | (n18959 & n29711) | (n18974 & n29711);
  assign n34781 = (n18671 & n34779) | (n18671 & n34780) | (n34779 & n34780);
  assign n29713 = n18856 | n18974;
  assign n34782 = n29705 | n29713;
  assign n34783 = n18959 | n29713;
  assign n34784 = (n18671 & n34782) | (n18671 & n34783) | (n34782 & n34783);
  assign n18977 = ~n34781 & n34784;
  assign n18978 = x121 & x147;
  assign n18979 = n18977 & n18978;
  assign n18980 = n18977 | n18978;
  assign n18981 = ~n18979 & n18980;
  assign n18982 = x120 & x148;
  assign n18983 = n18981 & n18982;
  assign n18984 = n18981 | n18982;
  assign n18985 = ~n18983 & n18984;
  assign n29715 = n18674 | n18874;
  assign n29716 = n18736 | n29715;
  assign n18987 = n18754 | n18873;
  assign n34785 = n18866 | n18987;
  assign n34786 = (n18866 & n18867) | (n18866 & n34785) | (n18867 & n34785);
  assign n29718 = (n18866 & n29716) | (n18866 & n34786) | (n29716 & n34786);
  assign n18991 = n18985 | n29718;
  assign n18992 = n18985 & n29718;
  assign n18993 = n18991 & ~n18992;
  assign n18994 = x119 & x149;
  assign n18995 = n18993 | n18994;
  assign n18996 = n18993 & n18994;
  assign n18997 = n18995 & ~n18996;
  assign n18998 = n18958 | n18997;
  assign n18999 = n18958 & n18997;
  assign n19000 = n18998 & ~n18999;
  assign n19001 = x118 & x150;
  assign n19002 = n19000 | n19001;
  assign n19003 = n19000 & n19001;
  assign n19004 = n19002 & ~n19003;
  assign n29719 = n18885 & n29678;
  assign n29720 = n18885 & n18896;
  assign n29721 = (n29622 & n29719) | (n29622 & n29720) | (n29719 & n29720);
  assign n29722 = n18878 | n29651;
  assign n29723 = n18839 | n18878;
  assign n29724 = (n29624 & n29722) | (n29624 & n29723) | (n29722 & n29723);
  assign n19007 = n18879 & ~n29698;
  assign n19008 = n29724 & n19007;
  assign n19009 = n29721 | n19008;
  assign n19010 = n19004 | n19009;
  assign n19011 = n19004 & n19009;
  assign n19012 = n19010 & ~n19011;
  assign n29725 = n18885 | n29678;
  assign n29726 = n18885 | n18896;
  assign n29727 = (n29622 & n29725) | (n29622 & n29726) | (n29725 & n29726);
  assign n19014 = n18886 & ~n29721;
  assign n19015 = n29727 & n19014;
  assign n29728 = n18900 | n19015;
  assign n29730 = n19012 | n29728;
  assign n29731 = n19012 | n19015;
  assign n29732 = (n29683 & n29730) | (n29683 & n29731) | (n29730 & n29731);
  assign n29733 = n19012 & n29728;
  assign n29734 = n19012 & n19015;
  assign n29735 = (n29683 & n29733) | (n29683 & n29734) | (n29733 & n29734);
  assign n19019 = n29732 & ~n29735;
  assign n19020 = n18952 & n19019;
  assign n19021 = n18952 | n19019;
  assign n19022 = ~n19020 & n19021;
  assign n19023 = n29695 & n19022;
  assign n19024 = n29695 | n19022;
  assign n19025 = ~n19023 & n19024;
  assign n19026 = n18950 | n19025;
  assign n19027 = n18950 & n19025;
  assign n19028 = n19026 & ~n19027;
  assign n29736 = n18914 & n18915;
  assign n29737 = (n18914 & n18918) | (n18914 & n29736) | (n18918 & n29736);
  assign n19031 = n19028 & ~n29737;
  assign n19032 = ~n19028 & n29737;
  assign n19033 = n19031 | n19032;
  assign n19034 = x115 & x153;
  assign n19035 = n19033 | n19034;
  assign n19036 = n19033 & n19034;
  assign n19037 = n19035 & ~n19036;
  assign n19038 = ~n18949 & n19037;
  assign n19039 = n18949 & ~n19037;
  assign n19040 = n19038 | n19039;
  assign n19041 = n18820 | n18934;
  assign n19042 = n18935 & n19041;
  assign n19043 = n19040 & ~n19042;
  assign n19044 = ~n19040 & n19042;
  assign n19045 = n19043 | n19044;
  assign n19046 = x113 & x155;
  assign n19047 = n19045 | n19046;
  assign n19048 = n19045 & n19046;
  assign n19049 = n19047 & ~n19048;
  assign n19050 = ~n18941 & n19049;
  assign n19051 = n18941 & ~n19049;
  assign n19052 = n19050 | n19051;
  assign n19053 = x112 & x156;
  assign n19054 = n19052 & n19053;
  assign n19055 = n19052 | n19053;
  assign n19056 = ~n19054 & n19055;
  assign n18945 = n18923 & n18944;
  assign n29738 = n19035 & n19036;
  assign n29739 = (n18945 & n19035) | (n18945 & n29738) | (n19035 & n29738);
  assign n19059 = x115 & x154;
  assign n19060 = n29739 & n19059;
  assign n19061 = n29739 | n19059;
  assign n19062 = ~n19060 & n19061;
  assign n19063 = x117 & x152;
  assign n19065 = x118 & x151;
  assign n29742 = n18957 & n18993;
  assign n29743 = (n18993 & n29698) | (n18993 & n29742) | (n29698 & n29742);
  assign n34787 = n18981 & n34786;
  assign n34788 = n18866 & n18981;
  assign n34789 = (n29716 & n34787) | (n29716 & n34788) | (n34787 & n34788);
  assign n34790 = (n18982 & n18983) | (n18982 & n34786) | (n18983 & n34786);
  assign n37727 = n18864 & n18982;
  assign n37728 = n18863 & n37727;
  assign n37288 = (n18981 & n18982) | (n18981 & n37728) | (n18982 & n37728);
  assign n34792 = (n29716 & n34790) | (n29716 & n37288) | (n34790 & n37288);
  assign n19070 = ~n34789 & n34792;
  assign n19071 = n29743 | n19070;
  assign n19094 = x122 & x147;
  assign n29706 = (n18671 & n18959) | (n18671 & n29705) | (n18959 & n29705);
  assign n19075 = x125 & x144;
  assign n19076 = x124 & x145;
  assign n19077 = n19075 & n19076;
  assign n19078 = n19075 | n19076;
  assign n19079 = ~n19077 & n19078;
  assign n19080 = x123 & x146;
  assign n19081 = n19079 & n19080;
  assign n19082 = n19079 | n19080;
  assign n19083 = ~n19081 & n19082;
  assign n19073 = n18964 & n18965;
  assign n34793 = n18849 | n19073;
  assign n34794 = (n18968 & n19073) | (n18968 & n34793) | (n19073 & n34793);
  assign n29750 = n19083 & ~n34794;
  assign n29748 = n18968 | n19073;
  assign n29751 = n19083 & ~n29748;
  assign n29752 = (~n34764 & n29750) | (~n34764 & n29751) | (n29750 & n29751);
  assign n29753 = ~n19083 & n34794;
  assign n29754 = ~n19083 & n29748;
  assign n29755 = (n34764 & n29753) | (n34764 & n29754) | (n29753 & n29754);
  assign n19086 = n29752 | n29755;
  assign n19087 = n18972 | n19086;
  assign n29756 = n19087 | n29711;
  assign n29757 = n18974 | n19087;
  assign n29758 = (n29706 & n29756) | (n29706 & n29757) | (n29756 & n29757);
  assign n19091 = n18973 & n19086;
  assign n19089 = n18856 | n18972;
  assign n29759 = n19089 & n19091;
  assign n34795 = (n19091 & n29705) | (n19091 & n29759) | (n29705 & n29759);
  assign n34796 = (n18959 & n19091) | (n18959 & n29759) | (n19091 & n29759);
  assign n34797 = (n18671 & n34795) | (n18671 & n34796) | (n34795 & n34796);
  assign n34798 = ~n19094 & n34797;
  assign n34799 = (n19094 & n29758) | (n19094 & ~n34798) | (n29758 & ~n34798);
  assign n29761 = n19094 & ~n29759;
  assign n34800 = ~n19086 & n19094;
  assign n34801 = (~n18973 & n19094) | (~n18973 & n34800) | (n19094 & n34800);
  assign n29763 = (~n29706 & n29761) | (~n29706 & n34801) | (n29761 & n34801);
  assign n19097 = n29758 & n29763;
  assign n19099 = x121 & x148;
  assign n29764 = ~n19097 & n19099;
  assign n29765 = n34799 & n29764;
  assign n29766 = n19097 & ~n19099;
  assign n29767 = (n34799 & n19099) | (n34799 & ~n29766) | (n19099 & ~n29766);
  assign n19102 = ~n29765 & n29767;
  assign n29745 = n18979 | n18981;
  assign n29768 = n19102 & ~n29745;
  assign n29769 = ~n18979 & n19102;
  assign n29770 = (~n29718 & n29768) | (~n29718 & n29769) | (n29768 & n29769);
  assign n29771 = ~n19102 & n29745;
  assign n29772 = n18979 & ~n19102;
  assign n29773 = (n29718 & n29771) | (n29718 & n29772) | (n29771 & n29772);
  assign n19105 = n29770 | n29773;
  assign n19106 = x120 & x149;
  assign n19107 = n19105 | n19106;
  assign n19108 = n19105 & n19106;
  assign n19109 = n19107 & ~n19108;
  assign n19110 = n19071 | n19109;
  assign n19111 = n19071 & n19109;
  assign n19112 = n19110 & ~n19111;
  assign n19113 = x119 & x150;
  assign n19114 = n19112 | n19113;
  assign n19115 = n19112 & n19113;
  assign n19116 = n19114 & ~n19115;
  assign n29774 = n19000 & n19008;
  assign n29775 = (n19000 & n29721) | (n19000 & n29774) | (n29721 & n29774);
  assign n29776 = n18957 | n18993;
  assign n29777 = n29698 | n29776;
  assign n19119 = n18994 & ~n29743;
  assign n19120 = n29777 & n19119;
  assign n19121 = n29775 | n19120;
  assign n19122 = n19116 | n19121;
  assign n19123 = n19116 & n19121;
  assign n19124 = n19122 & ~n19123;
  assign n29778 = n19000 | n19008;
  assign n29779 = n29721 | n29778;
  assign n19126 = n19001 & ~n29775;
  assign n19127 = n29779 & n19126;
  assign n29780 = n19124 & n19127;
  assign n29781 = (n19124 & n29735) | (n19124 & n29780) | (n29735 & n29780);
  assign n29782 = n19124 | n19127;
  assign n29783 = n29735 | n29782;
  assign n19131 = ~n29781 & n29783;
  assign n19132 = n19065 & n19131;
  assign n19133 = n19065 | n19131;
  assign n19134 = ~n19132 & n19133;
  assign n29740 = n19020 | n19022;
  assign n29784 = n19134 & n29740;
  assign n29785 = n19020 & n19134;
  assign n29786 = (n29695 & n29784) | (n29695 & n29785) | (n29784 & n29785);
  assign n29787 = n19134 | n29740;
  assign n29788 = n19020 | n19134;
  assign n29789 = (n29695 & n29787) | (n29695 & n29788) | (n29787 & n29788);
  assign n19137 = ~n29786 & n29789;
  assign n19138 = n19063 | n19137;
  assign n19139 = n19063 & n19137;
  assign n19140 = n19138 & ~n19139;
  assign n29790 = n19026 & n19027;
  assign n29791 = (n19026 & n29737) | (n19026 & n29790) | (n29737 & n29790);
  assign n19143 = n19140 & ~n29791;
  assign n19144 = ~n19140 & n29791;
  assign n19145 = n19143 | n19144;
  assign n19146 = x116 & x153;
  assign n19147 = n19145 | n19146;
  assign n19148 = n19145 & n19146;
  assign n19149 = n19147 & ~n19148;
  assign n19150 = ~n19062 & n19149;
  assign n19151 = n19062 & ~n19149;
  assign n19152 = n19150 | n19151;
  assign n19153 = ~n18945 & n19037;
  assign n19154 = n18945 & ~n19037;
  assign n19155 = n19153 | n19154;
  assign n19158 = n18946 | n19155;
  assign n19156 = n18946 & n19155;
  assign n29792 = n19156 & n19158;
  assign n29793 = (n19042 & n19158) | (n19042 & n29792) | (n19158 & n29792);
  assign n19160 = n19152 & ~n29793;
  assign n19161 = ~n19152 & n29793;
  assign n19162 = n19160 | n19161;
  assign n19163 = x114 & x155;
  assign n19164 = n19162 | n19163;
  assign n19165 = n19162 & n19163;
  assign n19166 = n19164 & ~n19165;
  assign n19167 = n18941 | n19048;
  assign n19168 = n19047 & n19167;
  assign n19169 = n19166 & ~n19168;
  assign n19170 = ~n19166 & n19168;
  assign n19171 = n19169 | n19170;
  assign n19172 = x113 & x156;
  assign n19173 = n19171 & ~n19172;
  assign n19174 = ~n19171 & n19172;
  assign n19175 = n19173 | n19174;
  assign n19176 = ~n19054 & n19175;
  assign n19177 = n19054 & ~n19175;
  assign n19178 = n19176 | n19177;
  assign n19179 = x112 & x157;
  assign n19180 = n19178 & n19179;
  assign n19181 = n19178 | n19179;
  assign n19182 = ~n19180 & n19181;
  assign n19183 = x114 & x156;
  assign n29794 = n19164 & n19165;
  assign n29795 = (n19164 & n19168) | (n19164 & n29794) | (n19168 & n29794);
  assign n29796 = n19138 & n19139;
  assign n29797 = (n19138 & n29791) | (n19138 & n29796) | (n29791 & n29796);
  assign n29798 = n19112 & n19120;
  assign n29799 = (n19112 & n29775) | (n19112 & n29798) | (n29775 & n29798);
  assign n29800 = n19070 & n19105;
  assign n29801 = (n19105 & n29743) | (n19105 & n29800) | (n29743 & n29800);
  assign n34802 = n19070 & n19106;
  assign n34803 = (n19105 & n19106) | (n19105 & n34802) | (n19106 & n34802);
  assign n29805 = (n19106 & n29743) | (n19106 & n34803) | (n29743 & n34803);
  assign n19193 = ~n29801 & n29805;
  assign n19098 = n34799 & ~n19097;
  assign n29806 = n19098 | n29745;
  assign n29807 = n18979 | n19098;
  assign n29808 = (n29718 & n29806) | (n29718 & n29807) | (n29806 & n29807);
  assign n19196 = n18866 | n18979;
  assign n18988 = n18867 & n18987;
  assign n29809 = n18988 | n19196;
  assign n29810 = (n19196 & n29716) | (n19196 & n29809) | (n29716 & n29809);
  assign n19198 = n18980 & ~n19097;
  assign n34804 = n19099 & ~n34799;
  assign n34805 = (n19099 & ~n19198) | (n19099 & n34804) | (~n19198 & n34804);
  assign n29812 = (n19099 & ~n29810) | (n19099 & n34805) | (~n29810 & n34805);
  assign n19202 = n29808 & n29812;
  assign n29813 = n19202 | n29800;
  assign n29814 = n19105 | n19202;
  assign n29815 = (n29743 & n29813) | (n29743 & n29814) | (n29813 & n29814);
  assign n19204 = x121 & x149;
  assign n19205 = x122 & x148;
  assign n19213 = x126 & x144;
  assign n19214 = x125 & x145;
  assign n19215 = n19213 | n19214;
  assign n19216 = n19213 & n19214;
  assign n19217 = n19215 & ~n19216;
  assign n19218 = n19078 & n19217;
  assign n29830 = n19077 | n34794;
  assign n29833 = n19218 & n29830;
  assign n34812 = n19073 | n19077;
  assign n34813 = n18968 | n34812;
  assign n29834 = n19218 & n34813;
  assign n29835 = (n34764 & n29833) | (n34764 & n29834) | (n29833 & n29834);
  assign n19220 = n19077 | n19217;
  assign n29818 = n19079 & n34794;
  assign n29836 = n19220 | n29818;
  assign n29819 = n19079 & n29748;
  assign n29837 = n19220 | n29819;
  assign n29838 = (n34764 & n29836) | (n34764 & n29837) | (n29836 & n29837);
  assign n19222 = ~n29835 & n29838;
  assign n19223 = x124 & x146;
  assign n19224 = n19222 & n19223;
  assign n19225 = n19222 | n19223;
  assign n19226 = ~n19224 & n19225;
  assign n29820 = (n34764 & n29818) | (n34764 & n29819) | (n29818 & n29819);
  assign n34808 = (n19080 & n19081) | (n19080 & n34794) | (n19081 & n34794);
  assign n34809 = (n19080 & n19081) | (n19080 & n29748) | (n19081 & n29748);
  assign n29826 = (n34764 & n34808) | (n34764 & n34809) | (n34808 & n34809);
  assign n19210 = ~n29820 & n29826;
  assign n37289 = n19210 & n19226;
  assign n37290 = (n19226 & n29759) | (n19226 & n37289) | (n29759 & n37289);
  assign n34810 = n19086 | n19210;
  assign n34811 = (n18973 & n19210) | (n18973 & n34810) | (n19210 & n34810);
  assign n34815 = n19226 & n34811;
  assign n34816 = (n29706 & n37290) | (n29706 & n34815) | (n37290 & n34815);
  assign n37291 = n19210 | n19226;
  assign n37292 = n29759 | n37291;
  assign n34818 = n19226 | n34811;
  assign n34819 = (n29706 & n37292) | (n29706 & n34818) | (n37292 & n34818);
  assign n19229 = ~n34816 & n34819;
  assign n19230 = x123 & x147;
  assign n19231 = n19229 & n19230;
  assign n19232 = n19229 | n19230;
  assign n19233 = ~n19231 & n19232;
  assign n34806 = n19097 | n34799;
  assign n34807 = (n19097 & n19198) | (n19097 & n34806) | (n19198 & n34806);
  assign n34820 = n19233 & n34807;
  assign n34821 = n19097 & n19233;
  assign n34822 = (n29810 & n34820) | (n29810 & n34821) | (n34820 & n34821);
  assign n34823 = n19233 | n34807;
  assign n34824 = n19097 | n19233;
  assign n34825 = (n29810 & n34823) | (n29810 & n34824) | (n34823 & n34824);
  assign n19236 = ~n34822 & n34825;
  assign n19237 = n19205 & n19236;
  assign n19238 = n19205 | n19236;
  assign n19239 = ~n19237 & n19238;
  assign n19240 = n19204 & n19239;
  assign n19241 = n19204 | n19239;
  assign n19242 = ~n19240 & n19241;
  assign n19243 = n29815 | n19242;
  assign n19244 = n29815 & n19242;
  assign n19245 = n19243 & ~n19244;
  assign n34826 = n19193 | n19245;
  assign n34827 = n29799 | n34826;
  assign n34828 = n19193 & n19245;
  assign n34829 = (n19245 & n29799) | (n19245 & n34828) | (n29799 & n34828);
  assign n19248 = n34827 & ~n34829;
  assign n19249 = x120 & x150;
  assign n19250 = x119 & x151;
  assign n19251 = n19249 & n19250;
  assign n19252 = n19249 | n19250;
  assign n19253 = ~n19251 & n19252;
  assign n19254 = n19248 & n19253;
  assign n19255 = n19248 | n19253;
  assign n19256 = ~n19254 & n19255;
  assign n29839 = n19112 | n19120;
  assign n29840 = n29775 | n29839;
  assign n19258 = n19113 & ~n29799;
  assign n19259 = n29840 & n19258;
  assign n19260 = n29781 | n19259;
  assign n19261 = n19256 | n19260;
  assign n19262 = n19256 & n19260;
  assign n19263 = n19261 & ~n19262;
  assign n29841 = n19132 | n19263;
  assign n29842 = n29786 | n29841;
  assign n29843 = n19132 & n19263;
  assign n29844 = (n19263 & n29786) | (n19263 & n29843) | (n29786 & n29843);
  assign n19266 = n29842 & ~n29844;
  assign n19267 = x118 & x152;
  assign n19268 = x117 & x153;
  assign n19269 = n19267 & n19268;
  assign n19270 = n19267 | n19268;
  assign n19271 = ~n19269 & n19270;
  assign n19272 = n19266 & n19271;
  assign n19273 = n19266 | n19271;
  assign n19274 = ~n19272 & n19273;
  assign n19275 = n29797 & n19274;
  assign n19276 = n29797 | n19274;
  assign n19277 = ~n19275 & n19276;
  assign n19278 = x116 & x154;
  assign n19279 = ~n19277 & n19278;
  assign n19280 = n19277 & ~n19278;
  assign n19281 = n19279 | n19280;
  assign n29845 = n19147 & n19148;
  assign n29846 = (n19147 & n29739) | (n19147 & n29845) | (n29739 & n29845);
  assign n19284 = n19281 & ~n29846;
  assign n19285 = ~n19281 & n29846;
  assign n19286 = n19284 | n19285;
  assign n19287 = x115 & x155;
  assign n19288 = n19286 & ~n19287;
  assign n19289 = ~n19286 & n19287;
  assign n19290 = n19288 | n19289;
  assign n19291 = ~n29739 & n19149;
  assign n19292 = n29739 & ~n19149;
  assign n19293 = n19291 | n19292;
  assign n19296 = n19059 | n19293;
  assign n19294 = n19059 & n19293;
  assign n29847 = n19294 & n19296;
  assign n29848 = (n19296 & n29793) | (n19296 & n29847) | (n29793 & n29847);
  assign n19298 = n19290 & ~n29848;
  assign n19299 = ~n19290 & n29848;
  assign n19300 = n19298 | n19299;
  assign n19301 = n29795 & n19300;
  assign n19302 = n29795 | n19300;
  assign n19303 = ~n19301 & n19302;
  assign n19304 = n19183 | n19303;
  assign n19305 = n19183 & n19303;
  assign n19306 = n19304 & ~n19305;
  assign n29849 = n19053 & n19172;
  assign n29850 = n19052 & n29849;
  assign n19308 = n19171 | n29850;
  assign n29851 = n19053 | n19172;
  assign n29852 = (n19052 & n19172) | (n19052 & n29851) | (n19172 & n29851);
  assign n19310 = n19308 & n29852;
  assign n19311 = n19306 & ~n19310;
  assign n19312 = ~n19306 & n19310;
  assign n19313 = n19311 | n19312;
  assign n19314 = x113 & x157;
  assign n19315 = n19313 | n19314;
  assign n19316 = n19313 & n19314;
  assign n19317 = n19315 & ~n19316;
  assign n19318 = ~n19180 & n19317;
  assign n19319 = n19180 & ~n19317;
  assign n19320 = n19318 | n19319;
  assign n19321 = x112 & x158;
  assign n19322 = n19320 & n19321;
  assign n19323 = n19320 | n19321;
  assign n19324 = ~n19322 & n19323;
  assign n19325 = x113 & x158;
  assign n19326 = n19180 | n19316;
  assign n19327 = n19315 & n19326;
  assign n19328 = x115 & x156;
  assign n19334 = n19266 & n19267;
  assign n19335 = n19266 | n19267;
  assign n19336 = ~n19334 & n19335;
  assign n29857 = n19334 | n19336;
  assign n29858 = (n19334 & n29797) | (n19334 & n29857) | (n29797 & n29857);
  assign n19194 = n29799 | n19193;
  assign n19339 = n19245 | n19249;
  assign n19340 = n19245 & n19249;
  assign n19341 = n19339 & ~n19340;
  assign n19342 = n19194 | n19341;
  assign n19343 = n19194 & n19341;
  assign n19344 = n19342 & ~n19343;
  assign n34830 = n19259 & n19344;
  assign n34831 = (n19344 & n29781) | (n19344 & n34830) | (n29781 & n34830);
  assign n29859 = n19250 & n19344;
  assign n29860 = (n19250 & n19260) | (n19250 & n29859) | (n19260 & n29859);
  assign n19348 = ~n34831 & n29860;
  assign n29861 = n19348 | n29843;
  assign n29862 = n19263 | n19348;
  assign n29863 = (n29786 & n29861) | (n29786 & n29862) | (n29861 & n29862);
  assign n34833 = n19237 | n19239;
  assign n34834 = (n19237 & n29815) | (n19237 & n34833) | (n29815 & n34833);
  assign n19358 = x127 & x144;
  assign n19359 = x126 & x145;
  assign n19360 = n19358 & n19359;
  assign n19361 = n19358 | n19359;
  assign n19362 = ~n19360 & n19361;
  assign n19363 = x125 & x146;
  assign n19364 = n19362 | n19363;
  assign n19365 = n19362 & n19363;
  assign n19366 = n19364 & ~n19365;
  assign n29867 = n19216 | n29834;
  assign n34837 = n19366 | n29867;
  assign n37293 = n19078 | n19216;
  assign n37294 = (n19216 & n19217) | (n19216 & n37293) | (n19217 & n37293);
  assign n34836 = (n19216 & n29830) | (n19216 & n37294) | (n29830 & n37294);
  assign n34838 = n19366 | n34836;
  assign n34839 = (n34764 & n34837) | (n34764 & n34838) | (n34837 & n34838);
  assign n34840 = n19366 & n29867;
  assign n34841 = n19366 & n34836;
  assign n34842 = (n34764 & n34840) | (n34764 & n34841) | (n34840 & n34841);
  assign n19369 = n34839 & ~n34842;
  assign n19370 = n19225 & n19369;
  assign n29827 = n19210 | n29759;
  assign n29869 = n19224 & n19370;
  assign n34843 = (n19370 & n29827) | (n19370 & n29869) | (n29827 & n29869);
  assign n34844 = (n19370 & n29869) | (n19370 & n34811) | (n29869 & n34811);
  assign n34845 = (n29706 & n34843) | (n29706 & n34844) | (n34843 & n34844);
  assign n19372 = n19224 | n19369;
  assign n29871 = n19226 | n19372;
  assign n34846 = (n19372 & n29827) | (n19372 & n29871) | (n29827 & n29871);
  assign n34847 = (n19372 & n29871) | (n19372 & n34811) | (n29871 & n34811);
  assign n34848 = (n29706 & n34846) | (n29706 & n34847) | (n34846 & n34847);
  assign n19374 = ~n34845 & n34848;
  assign n19375 = x124 & x147;
  assign n19376 = n19374 & n19375;
  assign n19377 = n19374 | n19375;
  assign n19378 = ~n19376 & n19377;
  assign n19379 = n19231 | n19378;
  assign n29817 = (n19097 & n29810) | (n19097 & n34807) | (n29810 & n34807);
  assign n29873 = n19233 | n19379;
  assign n29874 = (n19379 & n29817) | (n19379 & n29873) | (n29817 & n29873);
  assign n19385 = x123 & x148;
  assign n19382 = n19232 & n19378;
  assign n34849 = n19231 & n19232;
  assign n34850 = n19378 & n34849;
  assign n34851 = (n19382 & n34807) | (n19382 & n34850) | (n34807 & n34850);
  assign n34852 = (n19097 & n19382) | (n19097 & n34850) | (n19382 & n34850);
  assign n34853 = (n29810 & n34851) | (n29810 & n34852) | (n34851 & n34852);
  assign n34854 = n19385 | n34853;
  assign n34855 = n29874 & ~n34854;
  assign n34856 = n19385 & n34853;
  assign n34857 = (n19385 & ~n29874) | (n19385 & n34856) | (~n29874 & n34856);
  assign n19388 = n34855 | n34857;
  assign n19389 = x122 & x149;
  assign n19390 = n19388 & n19389;
  assign n19391 = n19388 | n19389;
  assign n19392 = ~n19390 & n19391;
  assign n19393 = n34834 | n19392;
  assign n19394 = n34834 & n19392;
  assign n19395 = n19393 & ~n19394;
  assign n19350 = n29815 & n19239;
  assign n34832 = (n19204 & n19240) | (n19204 & n29815) | (n19240 & n29815);
  assign n19353 = ~n19350 & n34832;
  assign n29864 = n19245 | n19353;
  assign n34858 = n19395 | n29864;
  assign n34859 = n19353 | n19395;
  assign n34860 = (n19194 & n34858) | (n19194 & n34859) | (n34858 & n34859);
  assign n34861 = n19395 & n29864;
  assign n34862 = n19353 & n19395;
  assign n34863 = (n19194 & n34861) | (n19194 & n34862) | (n34861 & n34862);
  assign n19398 = n34860 & ~n34863;
  assign n19399 = x121 & x150;
  assign n19400 = x120 & x151;
  assign n19401 = n19399 & n19400;
  assign n19402 = n19399 | n19400;
  assign n19403 = ~n19401 & n19402;
  assign n19404 = n19398 & n19403;
  assign n19405 = n19398 | n19403;
  assign n19406 = ~n19404 & n19405;
  assign n19407 = n19248 & n19249;
  assign n29877 = n19344 | n19407;
  assign n29878 = (n19260 & n19407) | (n19260 & n29877) | (n19407 & n29877);
  assign n19409 = n19406 | n29878;
  assign n19410 = n19406 & n29878;
  assign n19411 = n19409 & ~n19410;
  assign n19412 = n29863 | n19411;
  assign n19413 = n29863 & n19411;
  assign n19414 = n19412 & ~n19413;
  assign n19415 = x119 & x152;
  assign n19416 = x118 & x153;
  assign n19417 = n19415 & n19416;
  assign n19418 = n19415 | n19416;
  assign n19419 = ~n19417 & n19418;
  assign n19420 = n19414 & n19419;
  assign n19421 = n19414 | n19419;
  assign n19422 = ~n19420 & n19421;
  assign n19423 = n29858 | n19422;
  assign n19424 = n29858 & n19422;
  assign n19425 = n19423 & ~n19424;
  assign n19426 = x117 & x154;
  assign n19427 = n19425 | n19426;
  assign n19428 = n19425 & n19426;
  assign n19429 = n19427 & ~n19428;
  assign n19431 = n29797 | n19336;
  assign n29879 = n19268 & ~n19336;
  assign n29880 = (n19268 & ~n29797) | (n19268 & n29879) | (~n29797 & n29879);
  assign n19433 = n19431 & n29880;
  assign n29881 = n19277 | n19433;
  assign n29882 = (n19433 & n29846) | (n19433 & n29881) | (n29846 & n29881);
  assign n19435 = ~n19429 & n29882;
  assign n19436 = n19429 & ~n29882;
  assign n19437 = n19435 | n19436;
  assign n19438 = x116 & x155;
  assign n19439 = n19437 & n19438;
  assign n19440 = n19437 | n19438;
  assign n19441 = ~n19439 & n19440;
  assign n19442 = n19277 | n29846;
  assign n29883 = (n19278 & n19279) | (n19278 & ~n29846) | (n19279 & ~n29846);
  assign n19444 = n19442 & n29883;
  assign n29884 = n19286 | n19444;
  assign n29885 = (n19444 & n29848) | (n19444 & n29884) | (n29848 & n29884);
  assign n19446 = ~n19441 & n29885;
  assign n19447 = n19441 & ~n29885;
  assign n19448 = n19446 | n19447;
  assign n19329 = n19286 & n29848;
  assign n29853 = n19286 & n19287;
  assign n29854 = (n19287 & n29848) | (n19287 & n29853) | (n29848 & n29853);
  assign n19332 = ~n19329 & n29854;
  assign n29855 = n19300 | n19332;
  assign n29886 = n19448 & n29855;
  assign n29887 = n19332 & n19448;
  assign n29888 = (n29795 & n29886) | (n29795 & n29887) | (n29886 & n29887);
  assign n29889 = n19448 | n29855;
  assign n29890 = n19332 | n19448;
  assign n29891 = (n29795 & n29889) | (n29795 & n29890) | (n29889 & n29890);
  assign n19451 = ~n29888 & n29891;
  assign n19452 = n19328 | n19451;
  assign n19453 = n19328 & n19451;
  assign n19454 = n19452 & ~n19453;
  assign n19455 = n19305 | n19310;
  assign n19456 = n19304 & n19455;
  assign n19457 = n19454 & ~n19456;
  assign n19458 = ~n19454 & n19456;
  assign n19459 = n19457 | n19458;
  assign n19460 = x114 & x157;
  assign n19461 = n19459 | n19460;
  assign n19462 = n19459 & n19460;
  assign n19463 = n19461 & ~n19462;
  assign n19464 = ~n19327 & n19463;
  assign n19465 = n19327 & ~n19463;
  assign n19466 = n19464 | n19465;
  assign n19467 = n19325 & ~n19466;
  assign n19468 = ~n19325 & n19466;
  assign n19469 = n19467 | n19468;
  assign n19470 = ~n19322 & n19469;
  assign n19471 = n19322 & ~n19469;
  assign n19472 = n19470 | n19471;
  assign n19473 = x112 & x159;
  assign n19474 = n19472 & n19473;
  assign n19475 = n19472 | n19473;
  assign n19476 = ~n19474 & n19475;
  assign n29892 = n19461 & n19462;
  assign n29893 = (n19327 & n19461) | (n19327 & n29892) | (n19461 & n29892);
  assign n19479 = x114 & x158;
  assign n19480 = n29893 & n19479;
  assign n19481 = n29893 | n19479;
  assign n19482 = ~n19480 & n19481;
  assign n19483 = x116 & x156;
  assign n19489 = n19414 & n19415;
  assign n19490 = n19414 | n19415;
  assign n19491 = ~n19489 & n19490;
  assign n29900 = n19489 | n19491;
  assign n29901 = (n19489 & n29858) | (n19489 & n29900) | (n29858 & n29900);
  assign n29865 = (n19194 & n19353) | (n19194 & n29864) | (n19353 & n29864);
  assign n34864 = n19385 & ~n34853;
  assign n34865 = n29874 & n34864;
  assign n37295 = n19237 | n34865;
  assign n37296 = (n19388 & n34865) | (n19388 & n37295) | (n34865 & n37295);
  assign n34867 = n19388 | n34865;
  assign n34868 = (n19350 & n37296) | (n19350 & n34867) | (n37296 & n34867);
  assign n19512 = x125 & x147;
  assign n19515 = x128 & x144;
  assign n19516 = x127 & x145;
  assign n19517 = n19515 & n19516;
  assign n19518 = n19515 | n19516;
  assign n19519 = ~n19517 & n19518;
  assign n29912 = n19360 | n19362;
  assign n29914 = n19519 | n29912;
  assign n29915 = n19360 | n19519;
  assign n34869 = (n29867 & n29914) | (n29867 & n29915) | (n29914 & n29915);
  assign n34870 = (n29914 & n29915) | (n29914 & n34836) | (n29915 & n34836);
  assign n34871 = (n34764 & n34869) | (n34764 & n34870) | (n34869 & n34870);
  assign n29917 = n19519 & n29912;
  assign n29918 = n19360 & n19519;
  assign n34872 = (n29867 & n29917) | (n29867 & n29918) | (n29917 & n29918);
  assign n34873 = (n29917 & n29918) | (n29917 & n34836) | (n29918 & n34836);
  assign n34874 = (n34764 & n34872) | (n34764 & n34873) | (n34872 & n34873);
  assign n19522 = n34871 & ~n34874;
  assign n19523 = x126 & x146;
  assign n19524 = n19522 & n19523;
  assign n19525 = n19522 | n19523;
  assign n19526 = ~n19524 & n19525;
  assign n37297 = n19216 | n19362;
  assign n37298 = n29834 | n37297;
  assign n37299 = n19362 | n37294;
  assign n37300 = (n29830 & n37297) | (n29830 & n37299) | (n37297 & n37299);
  assign n34877 = (n34764 & n37298) | (n34764 & n37300) | (n37298 & n37300);
  assign n37729 = ~n19216 & n19363;
  assign n37730 = (~n19362 & n19363) | (~n19362 & n37729) | (n19363 & n37729);
  assign n29920 = ~n19362 & n19363;
  assign n37303 = (~n29834 & n37730) | (~n29834 & n29920) | (n37730 & n29920);
  assign n37304 = (n19363 & n29920) | (n19363 & ~n37294) | (n29920 & ~n37294);
  assign n37305 = (~n29830 & n37730) | (~n29830 & n37304) | (n37730 & n37304);
  assign n34880 = (~n34764 & n37303) | (~n34764 & n37305) | (n37303 & n37305);
  assign n19529 = n34877 & n34880;
  assign n34881 = n19224 | n19529;
  assign n34882 = (n19370 & n19529) | (n19370 & n34881) | (n19529 & n34881);
  assign n29925 = n19526 & n34882;
  assign n34883 = n19369 | n19529;
  assign n34884 = (n19225 & n19529) | (n19225 & n34883) | (n19529 & n34883);
  assign n29926 = n19526 & n34884;
  assign n34885 = (n29827 & n29925) | (n29827 & n29926) | (n29925 & n29926);
  assign n34886 = (n29925 & n29926) | (n29925 & n34811) | (n29926 & n34811);
  assign n34887 = (n29706 & n34885) | (n29706 & n34886) | (n34885 & n34886);
  assign n29928 = n19526 | n34882;
  assign n29929 = n19526 | n34884;
  assign n34888 = (n29827 & n29928) | (n29827 & n29929) | (n29928 & n29929);
  assign n34889 = (n29928 & n29929) | (n29928 & n34811) | (n29929 & n34811);
  assign n34890 = (n29706 & n34888) | (n29706 & n34889) | (n34888 & n34889);
  assign n19533 = ~n34887 & n34890;
  assign n19534 = n19512 & n19533;
  assign n19535 = n19512 | n19533;
  assign n19536 = ~n19534 & n19535;
  assign n29931 = n19376 & n19536;
  assign n29932 = (n19536 & n34853) | (n19536 & n29931) | (n34853 & n29931);
  assign n29933 = n19376 | n19536;
  assign n29934 = n34853 | n29933;
  assign n19540 = ~n29932 & n29934;
  assign n19541 = x124 & x148;
  assign n19542 = n19540 & n19541;
  assign n19543 = n19540 | n19541;
  assign n19544 = ~n19542 & n19543;
  assign n19545 = x123 & x149;
  assign n19546 = n19544 & n19545;
  assign n19547 = n19544 | n19545;
  assign n19548 = ~n19546 & n19547;
  assign n19549 = n34868 | n19548;
  assign n19550 = n34868 & n19548;
  assign n19551 = n19549 & ~n19550;
  assign n29906 = n19237 & n19388;
  assign n29907 = (n19350 & n19388) | (n19350 & n29906) | (n19388 & n29906);
  assign n37731 = n19205 & n19389;
  assign n37732 = n19236 & n37731;
  assign n37307 = (n19388 & n19389) | (n19388 & n37732) | (n19389 & n37732);
  assign n34892 = (n19350 & n19389) | (n19350 & n37307) | (n19389 & n37307);
  assign n19508 = ~n29907 & n34892;
  assign n29910 = n19395 | n19508;
  assign n29935 = n19551 | n29910;
  assign n29936 = n19508 | n19551;
  assign n29937 = (n29865 & n29935) | (n29865 & n29936) | (n29935 & n29936);
  assign n29938 = n19551 & n29910;
  assign n29939 = n19508 & n19551;
  assign n29940 = (n29865 & n29938) | (n29865 & n29939) | (n29938 & n29939);
  assign n19554 = n29937 & ~n29940;
  assign n19555 = x122 & x150;
  assign n19556 = x121 & x151;
  assign n19557 = n19555 & n19556;
  assign n19558 = n19555 | n19556;
  assign n19559 = ~n19557 & n19558;
  assign n19560 = n19554 & n19559;
  assign n19561 = n19554 | n19559;
  assign n19562 = ~n19560 & n19561;
  assign n19563 = n19398 & n19399;
  assign n19494 = n19395 | n19399;
  assign n19495 = n19395 & n19399;
  assign n19496 = n19494 & ~n19495;
  assign n19497 = n29865 | n19496;
  assign n19498 = n29865 & n19496;
  assign n19499 = n19497 & ~n19498;
  assign n29941 = n19499 | n19563;
  assign n29942 = (n19563 & n29878) | (n19563 & n29941) | (n29878 & n29941);
  assign n19565 = n19562 | n29942;
  assign n19566 = n19562 & n29942;
  assign n19567 = n19565 & ~n19566;
  assign n34893 = n19499 & n29877;
  assign n34894 = n19407 & n19499;
  assign n34895 = (n19260 & n34893) | (n19260 & n34894) | (n34893 & n34894);
  assign n29902 = n19400 & n19499;
  assign n29903 = (n19400 & n29878) | (n19400 & n29902) | (n29878 & n29902);
  assign n19503 = ~n34895 & n29903;
  assign n29904 = n19411 | n19503;
  assign n29943 = n19567 | n29904;
  assign n29944 = n19503 | n19567;
  assign n29945 = (n29863 & n29943) | (n29863 & n29944) | (n29943 & n29944);
  assign n29946 = n19567 & n29904;
  assign n29947 = n19503 & n19567;
  assign n29948 = (n29863 & n29946) | (n29863 & n29947) | (n29946 & n29947);
  assign n19570 = n29945 & ~n29948;
  assign n19571 = x120 & x152;
  assign n19572 = x119 & x153;
  assign n19573 = n19571 & n19572;
  assign n19574 = n19571 | n19572;
  assign n19575 = ~n19573 & n19574;
  assign n19576 = n19570 & n19575;
  assign n19577 = n19570 | n19575;
  assign n19578 = ~n19576 & n19577;
  assign n19579 = n29901 | n19578;
  assign n19580 = n29901 & n19578;
  assign n19581 = n19579 & ~n19580;
  assign n19582 = x118 & x154;
  assign n19583 = n19581 | n19582;
  assign n19584 = n19581 & n19582;
  assign n19585 = n19583 & ~n19584;
  assign n29949 = n19425 & n29881;
  assign n29950 = n19425 & n19433;
  assign n29951 = (n29846 & n29949) | (n29846 & n29950) | (n29949 & n29950);
  assign n19587 = n29858 | n19491;
  assign n29952 = n19416 & ~n19491;
  assign n29953 = (n19416 & ~n29858) | (n19416 & n29952) | (~n29858 & n29952);
  assign n19589 = n19587 & n29953;
  assign n19590 = n29951 | n19589;
  assign n19591 = ~n19585 & n19590;
  assign n19592 = n19585 & ~n19590;
  assign n19593 = n19591 | n19592;
  assign n19594 = x117 & x155;
  assign n19595 = n19593 & n19594;
  assign n19596 = n19593 | n19594;
  assign n19597 = ~n19595 & n19596;
  assign n29897 = n19437 & n29884;
  assign n29898 = n19437 & n19444;
  assign n29899 = (n29848 & n29897) | (n29848 & n29898) | (n29897 & n29898);
  assign n29954 = n19425 | n29881;
  assign n29955 = n19425 | n19433;
  assign n29956 = (n29846 & n29954) | (n29846 & n29955) | (n29954 & n29955);
  assign n19599 = n19426 & ~n29951;
  assign n19600 = n29956 & n19599;
  assign n19601 = n29899 | n19600;
  assign n19602 = ~n19597 & n19601;
  assign n19603 = n19597 & ~n19601;
  assign n19604 = n19602 | n19603;
  assign n29894 = n19437 | n29884;
  assign n29895 = n19437 | n19444;
  assign n29896 = (n29848 & n29894) | (n29848 & n29895) | (n29894 & n29895);
  assign n19486 = n19438 & ~n29899;
  assign n19487 = n29896 & n19486;
  assign n29957 = n19487 & n19604;
  assign n29958 = (n19604 & n29888) | (n19604 & n29957) | (n29888 & n29957);
  assign n29959 = n19487 | n19604;
  assign n29960 = n29888 | n29959;
  assign n19607 = ~n29958 & n29960;
  assign n19608 = n19483 | n19607;
  assign n19609 = n19483 & n19607;
  assign n19610 = n19608 & ~n19609;
  assign n29961 = n19304 | n19453;
  assign n29962 = (n19453 & n19455) | (n19453 & n29961) | (n19455 & n29961);
  assign n19612 = n19452 & n29962;
  assign n19613 = n19610 & ~n19612;
  assign n19614 = ~n19610 & n19612;
  assign n19615 = n19613 | n19614;
  assign n19616 = x115 & x157;
  assign n19617 = n19615 | n19616;
  assign n19618 = n19615 & n19616;
  assign n19619 = n19617 & ~n19618;
  assign n19620 = ~n19482 & n19619;
  assign n19621 = n19482 & ~n19619;
  assign n19622 = n19620 | n19621;
  assign n29963 = n19321 & n19325;
  assign n29964 = n19320 & n29963;
  assign n19624 = n19466 | n29964;
  assign n29965 = n19321 | n19325;
  assign n29966 = (n19320 & n19325) | (n19320 & n29965) | (n19325 & n29965);
  assign n19626 = n19624 & n29966;
  assign n19627 = n19622 & ~n19626;
  assign n19628 = ~n19622 & n19626;
  assign n19629 = n19627 | n19628;
  assign n19630 = x113 & x159;
  assign n19631 = n19629 | n19630;
  assign n19632 = n19629 & n19630;
  assign n19633 = n19631 & ~n19632;
  assign n19634 = ~n19474 & n19633;
  assign n19635 = n19474 & ~n19633;
  assign n19636 = n19634 | n19635;
  assign n19637 = x112 & x160;
  assign n19638 = n19636 & n19637;
  assign n19639 = n19636 | n19637;
  assign n19640 = ~n19638 & n19639;
  assign n29967 = n19617 & n19618;
  assign n29968 = (n19617 & n29893) | (n19617 & n29967) | (n29893 & n29967);
  assign n19643 = x115 & x158;
  assign n19644 = n29968 & n19643;
  assign n19645 = n29968 | n19643;
  assign n19646 = ~n19644 & n19645;
  assign n19647 = x117 & x156;
  assign n19653 = n19570 & n19571;
  assign n19654 = n19570 | n19571;
  assign n19655 = ~n19653 & n19654;
  assign n29973 = n19653 | n19655;
  assign n29974 = (n19653 & n29901) | (n19653 & n29973) | (n29901 & n29973);
  assign n34896 = (n19508 & n29864) | (n19508 & n29910) | (n29864 & n29910);
  assign n34897 = (n19353 & n19508) | (n19353 & n29910) | (n19508 & n29910);
  assign n34898 = (n19194 & n34896) | (n19194 & n34897) | (n34896 & n34897);
  assign n19658 = n19551 | n19555;
  assign n19659 = n19551 & n19555;
  assign n19660 = n19658 & ~n19659;
  assign n19661 = n34898 | n19660;
  assign n19662 = n34898 & n19660;
  assign n19663 = n19661 & ~n19662;
  assign n34899 = n19663 & n29941;
  assign n34900 = n19563 & n19663;
  assign n34901 = (n29878 & n34899) | (n29878 & n34900) | (n34899 & n34900);
  assign n29975 = n19556 & n19663;
  assign n34902 = (n19556 & n29941) | (n19556 & n29975) | (n29941 & n29975);
  assign n34903 = (n19556 & n19563) | (n19556 & n29975) | (n19563 & n29975);
  assign n34904 = (n29878 & n34902) | (n29878 & n34903) | (n34902 & n34903);
  assign n19667 = ~n34901 & n34904;
  assign n19668 = n29948 | n19667;
  assign n19669 = x122 & x151;
  assign n29977 = n34865 | n19544;
  assign n29978 = n29907 | n29977;
  assign n29979 = n34865 & n19544;
  assign n29980 = (n19544 & n29907) | (n19544 & n29979) | (n29907 & n29979);
  assign n19672 = n29978 & ~n29980;
  assign n19673 = n19545 & n19672;
  assign n34905 = n19673 | n29939;
  assign n34906 = n19673 | n29938;
  assign n34907 = (n29865 & n34905) | (n29865 & n34906) | (n34905 & n34906);
  assign n29981 = n34865 | n19542;
  assign n34908 = n29906 | n29981;
  assign n34909 = n19388 | n29981;
  assign n34910 = (n19350 & n34908) | (n19350 & n34909) | (n34908 & n34909);
  assign n19678 = x129 & x144;
  assign n19679 = x128 & x145;
  assign n19680 = n19678 & n19679;
  assign n19681 = n19678 | n19679;
  assign n19682 = ~n19680 & n19681;
  assign n19683 = x127 & x146;
  assign n19684 = n19682 & n19683;
  assign n19685 = n19682 | n19683;
  assign n19686 = ~n19684 & n19685;
  assign n34911 = n19517 | n19519;
  assign n34912 = (n19517 & n29912) | (n19517 & n34911) | (n29912 & n34911);
  assign n29986 = n19686 & ~n34912;
  assign n30067 = n19360 | n19517;
  assign n34913 = (n19517 & n19519) | (n19517 & n30067) | (n19519 & n30067);
  assign n29987 = n19686 & ~n34913;
  assign n34914 = (~n29867 & n29986) | (~n29867 & n29987) | (n29986 & n29987);
  assign n34915 = (n29986 & n29987) | (n29986 & ~n34836) | (n29987 & ~n34836);
  assign n34916 = (~n34764 & n34914) | (~n34764 & n34915) | (n34914 & n34915);
  assign n29989 = ~n19686 & n34912;
  assign n29990 = ~n19686 & n34913;
  assign n34917 = (n29867 & n29989) | (n29867 & n29990) | (n29989 & n29990);
  assign n34918 = (n29989 & n29990) | (n29989 & n34836) | (n29990 & n34836);
  assign n34919 = (n34764 & n34917) | (n34764 & n34918) | (n34917 & n34918);
  assign n19689 = n34916 | n34919;
  assign n29992 = n19524 | n19689;
  assign n29993 = n34887 | n29992;
  assign n29994 = n19524 | n34882;
  assign n29995 = n19524 | n34884;
  assign n34920 = (n29827 & n29994) | (n29827 & n29995) | (n29994 & n29995);
  assign n34921 = (n29994 & n29995) | (n29994 & n34811) | (n29995 & n34811);
  assign n34922 = (n29706 & n34920) | (n29706 & n34921) | (n34920 & n34921);
  assign n19692 = n19525 & n19689;
  assign n19693 = n34922 & n19692;
  assign n19694 = n29993 & ~n19693;
  assign n19695 = x126 & x147;
  assign n19696 = n19694 & n19695;
  assign n19697 = n19694 | n19695;
  assign n19698 = ~n19696 & n19697;
  assign n30047 = n19376 | n19534;
  assign n34923 = (n19534 & n19536) | (n19534 & n30047) | (n19536 & n30047);
  assign n30000 = n19698 | n34923;
  assign n29998 = n19534 | n19536;
  assign n30001 = n19698 | n29998;
  assign n30002 = (n34853 & n30000) | (n34853 & n30001) | (n30000 & n30001);
  assign n30003 = n19698 & n34923;
  assign n30004 = n19698 & n29998;
  assign n30005 = (n34853 & n30003) | (n34853 & n30004) | (n30003 & n30004);
  assign n19702 = n30002 & ~n30005;
  assign n19703 = x125 & x148;
  assign n19704 = n19702 & ~n19703;
  assign n19705 = ~n19702 & n19703;
  assign n19706 = n19704 | n19705;
  assign n19707 = x124 & x149;
  assign n19708 = n19706 | n19707;
  assign n19709 = n19706 & n19707;
  assign n19710 = n19708 & ~n19709;
  assign n19711 = n19543 & n19710;
  assign n19712 = n34910 & n19711;
  assign n19713 = n19542 | n19710;
  assign n19714 = n29980 | n19713;
  assign n19715 = ~n19712 & n19714;
  assign n19716 = x123 & x150;
  assign n19717 = n19715 & n19716;
  assign n19718 = n19715 | n19716;
  assign n19719 = ~n19717 & n19718;
  assign n19720 = n34907 | n19719;
  assign n19721 = n34907 & n19719;
  assign n19722 = n19720 & ~n19721;
  assign n19723 = n19554 & n19555;
  assign n30006 = n19663 | n19723;
  assign n30008 = n19722 | n30006;
  assign n30009 = n19722 | n19723;
  assign n30010 = (n29942 & n30008) | (n29942 & n30009) | (n30008 & n30009);
  assign n30011 = n19722 & n30006;
  assign n30012 = n19722 & n19723;
  assign n30013 = (n29942 & n30011) | (n29942 & n30012) | (n30011 & n30012);
  assign n19727 = n30010 & ~n30013;
  assign n19728 = n19669 & n19727;
  assign n19729 = n19669 | n19727;
  assign n19730 = ~n19728 & n19729;
  assign n19731 = n19668 | n19730;
  assign n19732 = n19668 & n19730;
  assign n19733 = n19731 & ~n19732;
  assign n19734 = x121 & x152;
  assign n19735 = x120 & x153;
  assign n19736 = n19734 & n19735;
  assign n19737 = n19734 | n19735;
  assign n19738 = ~n19736 & n19737;
  assign n19739 = n19733 & n19738;
  assign n19740 = n19733 | n19738;
  assign n19741 = ~n19739 & n19740;
  assign n19742 = n29974 | n19741;
  assign n19743 = n29974 & n19741;
  assign n19744 = n19742 & ~n19743;
  assign n19745 = x119 & x154;
  assign n19746 = n19744 | n19745;
  assign n19747 = n19744 & n19745;
  assign n19748 = n19746 & ~n19747;
  assign n30014 = n19581 & n19589;
  assign n30015 = (n19581 & n29951) | (n19581 & n30014) | (n29951 & n30014);
  assign n19750 = n29901 | n19655;
  assign n30016 = n19572 & ~n19655;
  assign n30017 = (n19572 & ~n29901) | (n19572 & n30016) | (~n29901 & n30016);
  assign n19752 = n19750 & n30017;
  assign n19753 = n30015 | n19752;
  assign n19754 = ~n19748 & n19753;
  assign n19755 = n19748 & ~n19753;
  assign n19756 = n19754 | n19755;
  assign n19757 = x118 & x155;
  assign n19758 = n19756 & n19757;
  assign n19759 = n19756 | n19757;
  assign n19760 = ~n19758 & n19759;
  assign n29971 = n19593 & n19600;
  assign n29972 = (n19593 & n29899) | (n19593 & n29971) | (n29899 & n29971);
  assign n30018 = n19581 | n19589;
  assign n30019 = n29951 | n30018;
  assign n19762 = n19582 & ~n30015;
  assign n19763 = n30019 & n19762;
  assign n19764 = n29972 | n19763;
  assign n19765 = ~n19760 & n19764;
  assign n19766 = n19760 & ~n19764;
  assign n19767 = n19765 | n19766;
  assign n29969 = n19593 | n19600;
  assign n29970 = n29899 | n29969;
  assign n19650 = n19594 & ~n29972;
  assign n19651 = n29970 & n19650;
  assign n30020 = n19651 & n19767;
  assign n30021 = (n19767 & n29958) | (n19767 & n30020) | (n29958 & n30020);
  assign n30022 = n19651 | n19767;
  assign n30023 = n29958 | n30022;
  assign n19770 = ~n30021 & n30023;
  assign n19771 = n19647 | n19770;
  assign n19772 = n19647 & n19770;
  assign n19773 = n19771 & ~n19772;
  assign n30024 = n19452 | n19609;
  assign n30025 = (n19609 & n29962) | (n19609 & n30024) | (n29962 & n30024);
  assign n19775 = n19608 & n30025;
  assign n19776 = n19773 & ~n19775;
  assign n19777 = ~n19773 & n19775;
  assign n19778 = n19776 | n19777;
  assign n19779 = x116 & x157;
  assign n19780 = n19778 | n19779;
  assign n19781 = n19778 & n19779;
  assign n19782 = n19780 & ~n19781;
  assign n19783 = ~n19646 & n19782;
  assign n19784 = n19646 & ~n19782;
  assign n19785 = n19783 | n19784;
  assign n19786 = ~n29893 & n19619;
  assign n19787 = n29893 & ~n19619;
  assign n19788 = n19786 | n19787;
  assign n19789 = n19479 & n19788;
  assign n19790 = n19626 | n19789;
  assign n19791 = n19479 | n19788;
  assign n19792 = n19790 & n19791;
  assign n19793 = n19785 & ~n19792;
  assign n19794 = ~n19785 & n19792;
  assign n19795 = n19793 | n19794;
  assign n19796 = x114 & x159;
  assign n19797 = n19795 | n19796;
  assign n19798 = n19795 & n19796;
  assign n19799 = n19797 & ~n19798;
  assign n19800 = n19474 | n19632;
  assign n19801 = n19631 & n19800;
  assign n19802 = n19799 & ~n19801;
  assign n19803 = ~n19799 & n19801;
  assign n19804 = n19802 | n19803;
  assign n19805 = x113 & x160;
  assign n19806 = n19804 | n19805;
  assign n19807 = n19804 & n19805;
  assign n19808 = n19806 & ~n19807;
  assign n19809 = ~n19638 & n19808;
  assign n19810 = n19638 & ~n19808;
  assign n19811 = n19809 | n19810;
  assign n19812 = x112 & x161;
  assign n19813 = n19811 & n19812;
  assign n19814 = n19811 | n19812;
  assign n19815 = ~n19813 & n19814;
  assign n30026 = n19780 & n19781;
  assign n30027 = (n19780 & n29968) | (n19780 & n30026) | (n29968 & n30026);
  assign n19818 = x116 & x158;
  assign n19819 = n30027 & n19818;
  assign n19820 = n30027 | n19818;
  assign n19821 = ~n19819 & n19820;
  assign n19822 = x118 & x156;
  assign n19828 = n19733 & n19734;
  assign n19829 = n19733 | n19734;
  assign n19830 = ~n19828 & n19829;
  assign n30032 = n19828 | n19830;
  assign n30033 = (n19828 & n29974) | (n19828 & n30032) | (n29974 & n30032);
  assign n30034 = n19728 | n19730;
  assign n30035 = (n19668 & n19728) | (n19668 & n30034) | (n19728 & n30034);
  assign n30036 = n19673 | n19715;
  assign n30037 = n29940 | n30036;
  assign n30038 = n19673 | n29910;
  assign n34924 = n19508 | n19545;
  assign n34925 = (n19508 & n19672) | (n19508 & n34924) | (n19672 & n34924);
  assign n30040 = (n29865 & n30038) | (n29865 & n34925) | (n30038 & n34925);
  assign n19836 = n19545 | n19672;
  assign n19837 = n19715 & n19836;
  assign n34926 = n19716 & ~n19837;
  assign n34927 = (n19716 & ~n30040) | (n19716 & n34926) | (~n30040 & n34926);
  assign n19840 = n30037 & n34927;
  assign n30041 = n19542 & n19706;
  assign n34928 = (n19706 & n29979) | (n19706 & n30041) | (n29979 & n30041);
  assign n34929 = (n19544 & n19706) | (n19544 & n30041) | (n19706 & n30041);
  assign n34930 = (n29907 & n34928) | (n29907 & n34929) | (n34928 & n34929);
  assign n37308 = n19541 & n19707;
  assign n37309 = n19540 & n37308;
  assign n34932 = (n19706 & n19707) | (n19706 & n37309) | (n19707 & n37309);
  assign n34933 = (n19707 & n29979) | (n19707 & n34932) | (n29979 & n34932);
  assign n34934 = (n19544 & n19707) | (n19544 & n34932) | (n19707 & n34932);
  assign n34935 = (n29907 & n34933) | (n29907 & n34934) | (n34933 & n34934);
  assign n19846 = ~n34930 & n34935;
  assign n19849 = n19689 & ~n19695;
  assign n19850 = ~n19689 & n19695;
  assign n19851 = n19849 | n19850;
  assign n30049 = n19524 | n19851;
  assign n30050 = n34887 | n30049;
  assign n30051 = n19524 & n19851;
  assign n30052 = (n19851 & n34887) | (n19851 & n30051) | (n34887 & n30051);
  assign n30053 = n30050 & ~n30052;
  assign n30054 = n19535 & n30053;
  assign n30055 = n30047 & n30054;
  assign n30056 = (n34853 & n30054) | (n34853 & n30055) | (n30054 & n30055);
  assign n19857 = n30002 & ~n30056;
  assign n19858 = n19703 & n19857;
  assign n30058 = n19706 | n19858;
  assign n20049 = n19542 | n19858;
  assign n34936 = (n19706 & n19858) | (n19706 & n20049) | (n19858 & n20049);
  assign n34937 = (n29979 & n30058) | (n29979 & n34936) | (n30058 & n34936);
  assign n34938 = (n19544 & n30058) | (n19544 & n34936) | (n30058 & n34936);
  assign n34939 = (n29907 & n34937) | (n29907 & n34938) | (n34937 & n34938);
  assign n19869 = x130 & x144;
  assign n19870 = x129 & x145;
  assign n19871 = n19869 | n19870;
  assign n19872 = n19869 & n19870;
  assign n19873 = n19871 & ~n19872;
  assign n19874 = n19681 & n19873;
  assign n30078 = n19680 | n34913;
  assign n30081 = n19874 & n30078;
  assign n37310 = n19680 & n19681;
  assign n37311 = n19873 & n37310;
  assign n34941 = (n19874 & n34912) | (n19874 & n37311) | (n34912 & n37311);
  assign n34942 = (n29867 & n30081) | (n29867 & n34941) | (n30081 & n34941);
  assign n34943 = (n30081 & n34836) | (n30081 & n34941) | (n34836 & n34941);
  assign n34944 = (n34764 & n34942) | (n34764 & n34943) | (n34942 & n34943);
  assign n19876 = n19680 | n19873;
  assign n19863 = n19518 & n19682;
  assign n34945 = n19362 | n30067;
  assign n30069 = n19863 & n34945;
  assign n30083 = n19876 | n30069;
  assign n30070 = n19863 & n30067;
  assign n30084 = n19876 | n30070;
  assign n34946 = (n29867 & n30083) | (n29867 & n30084) | (n30083 & n30084);
  assign n34947 = (n30083 & n30084) | (n30083 & n34836) | (n30084 & n34836);
  assign n34948 = (n34764 & n34946) | (n34764 & n34947) | (n34946 & n34947);
  assign n19878 = ~n34944 & n34948;
  assign n19879 = x128 & x146;
  assign n19880 = n19878 & n19879;
  assign n19881 = n19878 | n19879;
  assign n19882 = ~n19880 & n19881;
  assign n30063 = n19682 | n34912;
  assign n30064 = n19682 | n34913;
  assign n34949 = (n29867 & n30063) | (n29867 & n30064) | (n30063 & n30064);
  assign n34950 = (n30063 & n30064) | (n30063 & n34836) | (n30064 & n34836);
  assign n34951 = (n34764 & n34949) | (n34764 & n34950) | (n34949 & n34950);
  assign n30072 = n19683 & ~n30069;
  assign n34952 = n19683 & ~n30067;
  assign n34953 = (n19683 & ~n19863) | (n19683 & n34952) | (~n19863 & n34952);
  assign n34954 = (~n29867 & n30072) | (~n29867 & n34953) | (n30072 & n34953);
  assign n34955 = (n30072 & ~n34836) | (n30072 & n34953) | (~n34836 & n34953);
  assign n34956 = (~n34764 & n34954) | (~n34764 & n34955) | (n34954 & n34955);
  assign n19866 = n34951 & n34956;
  assign n34957 = n19689 | n19866;
  assign n34958 = (n19525 & n19866) | (n19525 & n34957) | (n19866 & n34957);
  assign n30086 = n19882 & n34958;
  assign n30087 = n19866 & n19882;
  assign n30088 = (n34922 & n30086) | (n34922 & n30087) | (n30086 & n30087);
  assign n30089 = n19882 | n34958;
  assign n30090 = n19866 | n19882;
  assign n30091 = (n34922 & n30089) | (n34922 & n30090) | (n30089 & n30090);
  assign n19885 = ~n30088 & n30091;
  assign n19886 = x127 & x147;
  assign n19887 = n19885 & n19886;
  assign n19888 = n19885 | n19886;
  assign n19889 = ~n19887 & n19888;
  assign n30060 = n19696 | n30055;
  assign n30092 = n19889 & n30060;
  assign n30061 = n19696 | n30054;
  assign n30093 = n19889 & n30061;
  assign n30094 = (n34853 & n30092) | (n34853 & n30093) | (n30092 & n30093);
  assign n30095 = n19889 | n30060;
  assign n30096 = n19889 | n30061;
  assign n30097 = (n34853 & n30095) | (n34853 & n30096) | (n30095 & n30096);
  assign n19892 = ~n30094 & n30097;
  assign n19893 = x126 & x148;
  assign n19894 = n19892 & n19893;
  assign n19895 = n19892 | n19893;
  assign n19896 = ~n19894 & n19895;
  assign n19897 = x125 & x149;
  assign n19898 = n19896 & n19897;
  assign n19899 = n19896 | n19897;
  assign n19900 = ~n19898 & n19899;
  assign n19901 = n34939 | n19900;
  assign n19902 = n34939 & n19900;
  assign n19903 = n19901 & ~n19902;
  assign n30098 = ~n19846 & n19903;
  assign n34959 = ~n19837 & n30098;
  assign n34960 = (~n30040 & n30098) | (~n30040 & n34959) | (n30098 & n34959);
  assign n30100 = n19846 & ~n19903;
  assign n34961 = (n19837 & ~n19903) | (n19837 & n30100) | (~n19903 & n30100);
  assign n34962 = ~n19903 & n30100;
  assign n34963 = (n30040 & n34961) | (n30040 & n34962) | (n34961 & n34962);
  assign n19906 = n34960 | n34963;
  assign n19907 = x124 & x150;
  assign n19908 = x123 & x151;
  assign n19909 = n19907 & n19908;
  assign n19910 = n19907 | n19908;
  assign n19911 = ~n19909 & n19910;
  assign n19912 = n19906 & n19911;
  assign n19913 = n19906 | n19911;
  assign n19914 = ~n19912 & n19913;
  assign n34964 = n19840 | n19914;
  assign n34965 = n30013 | n34964;
  assign n34966 = n19840 & n19914;
  assign n34967 = (n19914 & n30013) | (n19914 & n34966) | (n30013 & n34966);
  assign n19917 = n34965 & ~n34967;
  assign n19918 = x122 & x152;
  assign n19919 = n19917 | n19918;
  assign n19920 = n19917 & n19918;
  assign n19921 = n19919 & ~n19920;
  assign n19922 = n30035 | n19921;
  assign n19923 = n30035 & n19921;
  assign n19924 = n19922 & ~n19923;
  assign n19925 = x121 & x153;
  assign n19926 = n19924 | n19925;
  assign n19927 = n19924 & n19925;
  assign n19928 = n19926 & ~n19927;
  assign n19929 = n30033 | n19928;
  assign n19930 = n30033 & n19928;
  assign n19931 = n19929 & ~n19930;
  assign n19932 = x120 & x154;
  assign n19933 = n19931 | n19932;
  assign n19934 = n19931 & n19932;
  assign n19935 = n19933 & ~n19934;
  assign n30102 = n19744 & n19752;
  assign n30103 = (n19744 & n30015) | (n19744 & n30102) | (n30015 & n30102);
  assign n19937 = n29974 | n19830;
  assign n30104 = n19735 & ~n19830;
  assign n30105 = (n19735 & ~n29974) | (n19735 & n30104) | (~n29974 & n30104);
  assign n19939 = n19937 & n30105;
  assign n19940 = n30103 | n19939;
  assign n19941 = ~n19935 & n19940;
  assign n19942 = n19935 & ~n19940;
  assign n19943 = n19941 | n19942;
  assign n19944 = x119 & x155;
  assign n19945 = n19943 & n19944;
  assign n19946 = n19943 | n19944;
  assign n19947 = ~n19945 & n19946;
  assign n30030 = n19756 & n19763;
  assign n30031 = (n19756 & n29972) | (n19756 & n30030) | (n29972 & n30030);
  assign n30106 = n19744 | n19752;
  assign n30107 = n30015 | n30106;
  assign n19949 = n19745 & ~n30103;
  assign n19950 = n30107 & n19949;
  assign n19951 = n30031 | n19950;
  assign n19952 = ~n19947 & n19951;
  assign n19953 = n19947 & ~n19951;
  assign n19954 = n19952 | n19953;
  assign n30028 = n19756 | n19763;
  assign n30029 = n29972 | n30028;
  assign n19825 = n19757 & ~n30031;
  assign n19826 = n30029 & n19825;
  assign n30108 = n19826 & n19954;
  assign n30109 = (n19954 & n30021) | (n19954 & n30108) | (n30021 & n30108);
  assign n30110 = n19826 | n19954;
  assign n30111 = n30021 | n30110;
  assign n19957 = ~n30109 & n30111;
  assign n19958 = n19822 | n19957;
  assign n19959 = n19822 & n19957;
  assign n19960 = n19958 & ~n19959;
  assign n30112 = n19608 | n19772;
  assign n30113 = (n19772 & n30025) | (n19772 & n30112) | (n30025 & n30112);
  assign n19962 = n19771 & n30113;
  assign n19963 = n19960 & ~n19962;
  assign n19964 = ~n19960 & n19962;
  assign n19965 = n19963 | n19964;
  assign n19966 = x117 & x157;
  assign n19967 = n19965 | n19966;
  assign n19968 = n19965 & n19966;
  assign n19969 = n19967 & ~n19968;
  assign n19970 = ~n19821 & n19969;
  assign n19971 = n19821 & ~n19969;
  assign n19972 = n19970 | n19971;
  assign n19973 = ~n29968 & n19782;
  assign n19974 = n29968 & ~n19782;
  assign n19975 = n19973 | n19974;
  assign n19978 = n19643 | n19975;
  assign n19976 = n19643 & n19975;
  assign n30114 = n19976 & n19978;
  assign n30115 = (n19792 & n19978) | (n19792 & n30114) | (n19978 & n30114);
  assign n19980 = n19972 & ~n30115;
  assign n19981 = ~n19972 & n30115;
  assign n19982 = n19980 | n19981;
  assign n19983 = x115 & x159;
  assign n19984 = n19982 | n19983;
  assign n19985 = n19982 & n19983;
  assign n19986 = n19984 & ~n19985;
  assign n30116 = n19797 & n19798;
  assign n30117 = (n19797 & n19801) | (n19797 & n30116) | (n19801 & n30116);
  assign n19989 = n19986 & ~n30117;
  assign n19990 = ~n19986 & n30117;
  assign n19991 = n19989 | n19990;
  assign n19992 = x114 & x160;
  assign n19993 = n19991 | n19992;
  assign n19994 = n19991 & n19992;
  assign n19995 = n19993 & ~n19994;
  assign n30118 = n19812 & n19995;
  assign n30119 = n19811 & n30118;
  assign n30120 = n19812 | n19995;
  assign n30121 = (n19811 & n19995) | (n19811 & n30120) | (n19995 & n30120);
  assign n19998 = ~n30119 & n30121;
  assign n19999 = n19638 | n19807;
  assign n20001 = x113 & x161;
  assign n34968 = n19805 & ~n20001;
  assign n34969 = (n19804 & ~n20001) | (n19804 & n34968) | (~n20001 & n34968);
  assign n30123 = n19999 & n34969;
  assign n34970 = ~n19805 & n20001;
  assign n34971 = ~n19804 & n34970;
  assign n30125 = (~n19999 & n20001) | (~n19999 & n34971) | (n20001 & n34971);
  assign n20004 = n30123 | n30125;
  assign n20005 = ~n19998 & n20004;
  assign n20006 = n19998 & ~n20004;
  assign n20007 = n20005 | n20006;
  assign n20008 = x112 & x162;
  assign n20009 = n20007 & n20008;
  assign n20010 = n20007 | n20008;
  assign n20011 = ~n20009 & n20010;
  assign n20012 = x114 & x161;
  assign n20000 = n19806 & n19999;
  assign n30126 = n19993 & n19994;
  assign n30127 = (n19993 & n20000) | (n19993 & n30126) | (n20000 & n30126);
  assign n20015 = x115 & x160;
  assign n30128 = n19984 & n19985;
  assign n30129 = (n19984 & n30117) | (n19984 & n30128) | (n30117 & n30128);
  assign n30130 = n19943 | n19950;
  assign n30131 = n30031 | n30130;
  assign n30132 = n19943 & n19950;
  assign n30133 = (n19943 & n30031) | (n19943 & n30132) | (n30031 & n30132);
  assign n20020 = n19944 & ~n30133;
  assign n20021 = n30131 & n20020;
  assign n30134 = n19931 & n19939;
  assign n30135 = (n19931 & n30103) | (n19931 & n30134) | (n30103 & n30134);
  assign n20024 = n30033 | n19924;
  assign n30136 = ~n19924 & n19925;
  assign n30137 = (n19925 & ~n30033) | (n19925 & n30136) | (~n30033 & n30136);
  assign n20027 = n20024 & n30137;
  assign n20028 = n30135 | n20027;
  assign n20029 = x122 & x153;
  assign n20030 = n30035 | n19917;
  assign n30138 = ~n19917 & n19918;
  assign n30139 = (n19918 & ~n30035) | (n19918 & n30138) | (~n30035 & n30138);
  assign n20033 = n20030 & n30139;
  assign n30140 = n19924 | n20033;
  assign n30141 = (n20033 & n30033) | (n20033 & n30140) | (n30033 & n30140);
  assign n20035 = x123 & x152;
  assign n20036 = n19906 & n19907;
  assign n20037 = n19906 | n19907;
  assign n20038 = ~n20036 & n20037;
  assign n34972 = n19840 & n20038;
  assign n34973 = (n20038 & n30013) | (n20038 & n34972) | (n30013 & n34972);
  assign n19841 = n30013 | n19840;
  assign n30142 = n19908 & n20038;
  assign n30143 = (n19841 & n19908) | (n19841 & n30142) | (n19908 & n30142);
  assign n20042 = ~n34973 & n30143;
  assign n30144 = n19917 | n20042;
  assign n30145 = (n20042 & n30035) | (n20042 & n30144) | (n30035 & n30144);
  assign n20044 = x124 & x151;
  assign n20046 = x125 & x150;
  assign n19838 = n30040 & n19837;
  assign n20051 = n19703 | n19857;
  assign n20052 = n19896 & n20051;
  assign n37312 = n19894 | n20049;
  assign n37313 = (n19894 & n20052) | (n19894 & n37312) | (n20052 & n37312);
  assign n37314 = n19894 | n20051;
  assign n37315 = (n19894 & n19896) | (n19894 & n37314) | (n19896 & n37314);
  assign n34979 = (n29980 & n37313) | (n29980 & n37315) | (n37313 & n37315);
  assign n29868 = (n34764 & n34836) | (n34764 & n29867) | (n34836 & n29867);
  assign n20060 = x131 & x144;
  assign n20061 = x130 & x145;
  assign n20062 = n20060 & n20061;
  assign n20063 = n20060 | n20061;
  assign n20064 = ~n20062 & n20063;
  assign n20065 = x129 & x146;
  assign n20066 = n20064 & n20065;
  assign n20067 = n20064 | n20065;
  assign n20068 = ~n20066 & n20067;
  assign n37318 = n19681 | n19872;
  assign n37319 = (n19872 & n19873) | (n19872 & n37318) | (n19873 & n37318);
  assign n37316 = n19872 | n37311;
  assign n37317 = (n34912 & n37319) | (n34912 & n37316) | (n37319 & n37316);
  assign n34983 = n20068 & ~n37317;
  assign n34982 = (n19872 & n30078) | (n19872 & n37319) | (n30078 & n37319);
  assign n34984 = n20068 & ~n34982;
  assign n34985 = (~n29868 & n34983) | (~n29868 & n34984) | (n34983 & n34984);
  assign n34986 = ~n20068 & n37317;
  assign n34987 = ~n20068 & n34982;
  assign n34988 = (n29868 & n34986) | (n29868 & n34987) | (n34986 & n34987);
  assign n20071 = n34985 | n34988;
  assign n37320 = n19880 | n20071;
  assign n37321 = n30086 | n37320;
  assign n30162 = n19866 | n19880;
  assign n34980 = (n19880 & n19882) | (n19880 & n30162) | (n19882 & n30162);
  assign n34990 = n20071 | n34980;
  assign n34991 = (n34922 & n37321) | (n34922 & n34990) | (n37321 & n34990);
  assign n20077 = x128 & x147;
  assign n30161 = n19880 | n34958;
  assign n20074 = n19881 & n20071;
  assign n37322 = ~n20074 & n20077;
  assign n37323 = (n20077 & ~n30161) | (n20077 & n37322) | (~n30161 & n37322);
  assign n30165 = n20074 & n30162;
  assign n34993 = n20077 & ~n30165;
  assign n34994 = (~n34922 & n37323) | (~n34922 & n34993) | (n37323 & n34993);
  assign n30168 = n34991 & n34994;
  assign n37324 = n20074 & ~n20077;
  assign n37325 = n30161 & n37324;
  assign n34996 = ~n20077 & n30165;
  assign n34997 = (n34922 & n37325) | (n34922 & n34996) | (n37325 & n34996);
  assign n30170 = (n34991 & n20077) | (n34991 & ~n34997) | (n20077 & ~n34997);
  assign n20080 = ~n30168 & n30170;
  assign n30171 = n19887 | n20080;
  assign n30172 = n30094 | n30171;
  assign n30173 = n19887 & n20080;
  assign n30174 = (n20080 & n30094) | (n20080 & n30173) | (n30094 & n30173);
  assign n20084 = n30172 & ~n30174;
  assign n20085 = x127 & x148;
  assign n20086 = n20084 & ~n20085;
  assign n20087 = ~n20084 & n20085;
  assign n20088 = n20086 | n20087;
  assign n20089 = x126 & x149;
  assign n20090 = n20088 & n20089;
  assign n20091 = n20088 | n20089;
  assign n20092 = ~n20090 & n20091;
  assign n20093 = n34979 | n20092;
  assign n20094 = n34979 & n20092;
  assign n20095 = n20093 & ~n20094;
  assign n20048 = n34939 | n19896;
  assign n37326 = n19897 & ~n20049;
  assign n37327 = (n19897 & ~n20052) | (n19897 & n37326) | (~n20052 & n37326);
  assign n37733 = ~n19703 & n19897;
  assign n37734 = ~n19857 & n37733;
  assign n37329 = (~n19896 & n19897) | (~n19896 & n37734) | (n19897 & n37734);
  assign n34976 = (~n29980 & n37327) | (~n29980 & n37329) | (n37327 & n37329);
  assign n20055 = n20048 & n34976;
  assign n30148 = n19846 & n19903;
  assign n30152 = n20055 | n30148;
  assign n34998 = n20095 & n30152;
  assign n30153 = n19903 | n20055;
  assign n34999 = n20095 & n30153;
  assign n35000 = (n19838 & n34998) | (n19838 & n34999) | (n34998 & n34999);
  assign n35001 = n20095 | n30152;
  assign n35002 = n20095 | n30153;
  assign n35003 = (n19838 & n35001) | (n19838 & n35002) | (n35001 & n35002);
  assign n20098 = ~n35000 & n35003;
  assign n20099 = n20046 & n20098;
  assign n20100 = n20046 | n20098;
  assign n20101 = ~n20099 & n20100;
  assign n30146 = n20036 | n20038;
  assign n35004 = n20101 | n30146;
  assign n35005 = n20036 | n20101;
  assign n35006 = (n19841 & n35004) | (n19841 & n35005) | (n35004 & n35005);
  assign n35007 = n20101 & n30146;
  assign n35008 = n20036 & n20101;
  assign n35009 = (n19841 & n35007) | (n19841 & n35008) | (n35007 & n35008);
  assign n20104 = n35006 & ~n35009;
  assign n20105 = n20044 & n20104;
  assign n20106 = n20044 | n20104;
  assign n20107 = ~n20105 & n20106;
  assign n20108 = n30145 & n20107;
  assign n20109 = n30145 | n20107;
  assign n20110 = ~n20108 & n20109;
  assign n20111 = n20035 & n20110;
  assign n20112 = n20035 | n20110;
  assign n20113 = ~n20111 & n20112;
  assign n20114 = n30141 & n20113;
  assign n20115 = n30141 | n20113;
  assign n20116 = ~n20114 & n20115;
  assign n20117 = n20029 | n20116;
  assign n20118 = n20029 & n20116;
  assign n20119 = n20117 & ~n20118;
  assign n20120 = ~n20028 & n20119;
  assign n20121 = n20028 & ~n20119;
  assign n20122 = n20120 | n20121;
  assign n20123 = x121 & x154;
  assign n20124 = x120 & x155;
  assign n20125 = n20123 & n20124;
  assign n20126 = n20123 | n20124;
  assign n20127 = ~n20125 & n20126;
  assign n20128 = n20122 & n20127;
  assign n20129 = n20122 | n20127;
  assign n20130 = ~n20128 & n20129;
  assign n30175 = n19931 | n19939;
  assign n30176 = n30103 | n30175;
  assign n20132 = n19932 & ~n30135;
  assign n20133 = n30176 & n20132;
  assign n20134 = n30133 | n20133;
  assign n20135 = n20130 | n20134;
  assign n20136 = n20130 & n20134;
  assign n20137 = n20135 & ~n20136;
  assign n30177 = n20021 | n20137;
  assign n30178 = n30109 | n30177;
  assign n30179 = n20021 & n20137;
  assign n30180 = (n20137 & n30109) | (n20137 & n30179) | (n30109 & n30179);
  assign n20140 = n30178 & ~n30180;
  assign n20141 = x119 & x156;
  assign n20142 = x118 & x157;
  assign n20143 = n20141 & n20142;
  assign n20144 = n20141 | n20142;
  assign n20145 = ~n20143 & n20144;
  assign n20146 = n20140 & n20145;
  assign n20147 = n20140 | n20145;
  assign n20148 = ~n20146 & n20147;
  assign n30181 = n19771 | n19959;
  assign n30182 = (n19959 & n30113) | (n19959 & n30181) | (n30113 & n30181);
  assign n20150 = n19958 & n30182;
  assign n20151 = n20148 | n20150;
  assign n20152 = n20148 & n20150;
  assign n20153 = n20151 & ~n20152;
  assign n20154 = x117 & x158;
  assign n20155 = ~n20153 & n20154;
  assign n20156 = n20153 & ~n20154;
  assign n20157 = n20155 | n20156;
  assign n30183 = n19967 & n19968;
  assign n30184 = (n19967 & n30027) | (n19967 & n30183) | (n30027 & n30183);
  assign n20160 = n20157 & ~n30184;
  assign n20161 = ~n20157 & n30184;
  assign n20162 = n20160 | n20161;
  assign n20163 = x116 & x159;
  assign n20164 = n20162 & ~n20163;
  assign n20165 = ~n20162 & n20163;
  assign n20166 = n20164 | n20165;
  assign n20167 = ~n30027 & n19969;
  assign n20168 = n30027 & ~n19969;
  assign n20169 = n20167 | n20168;
  assign n20172 = n19818 | n20169;
  assign n20170 = n19818 & n20169;
  assign n30185 = n20170 & n20172;
  assign n30186 = (n20172 & n30115) | (n20172 & n30185) | (n30115 & n30185);
  assign n20174 = n20166 & ~n30186;
  assign n20175 = ~n20166 & n30186;
  assign n20176 = n20174 | n20175;
  assign n20177 = n30129 & n20176;
  assign n20178 = n30129 | n20176;
  assign n20179 = ~n20177 & n20178;
  assign n20180 = n20015 & n20179;
  assign n20181 = n20015 | n20179;
  assign n20182 = ~n20180 & n20181;
  assign n20183 = n30127 & n20182;
  assign n20184 = n30127 | n20182;
  assign n20185 = ~n20183 & n20184;
  assign n20186 = n20012 | n20185;
  assign n20187 = n20012 & n20185;
  assign n20188 = n20186 & ~n20187;
  assign n30187 = n19812 & n20001;
  assign n30188 = n19811 & n30187;
  assign n20190 = n19995 & ~n20000;
  assign n20191 = ~n19995 & n20000;
  assign n20192 = n20190 | n20191;
  assign n20193 = n30188 | n20192;
  assign n30189 = n19812 | n20001;
  assign n30190 = (n19811 & n20001) | (n19811 & n30189) | (n20001 & n30189);
  assign n20195 = n20193 & n30190;
  assign n20196 = n20188 & n20195;
  assign n20197 = n20188 | n20195;
  assign n20198 = ~n20196 & n20197;
  assign n20199 = x113 & x162;
  assign n20200 = n20198 | n20199;
  assign n20201 = n20198 & n20199;
  assign n20202 = n20200 & ~n20201;
  assign n20203 = n20009 & ~n20202;
  assign n20204 = ~n20009 & n20202;
  assign n20205 = n20203 | n20204;
  assign n20206 = x112 & x163;
  assign n20207 = n20205 & n20206;
  assign n20208 = n20205 | n20206;
  assign n20209 = ~n20207 & n20208;
  assign n20210 = x114 & x162;
  assign n30191 = n20187 | n20195;
  assign n30192 = (n20187 & n20188) | (n20187 & n30191) | (n20188 & n30191);
  assign n20212 = x115 & x161;
  assign n20214 = x116 & x160;
  assign n20220 = n20140 & n20141;
  assign n20221 = n20140 | n20141;
  assign n20222 = ~n20220 & n20221;
  assign n30197 = n20220 | n20222;
  assign n30198 = (n20150 & n20220) | (n20150 & n30197) | (n20220 & n30197);
  assign n20225 = n20122 | n20123;
  assign n20226 = n20122 & n20123;
  assign n20227 = n20225 & ~n20226;
  assign n20228 = n20134 | n20227;
  assign n20229 = n20134 & n20227;
  assign n20230 = n20124 & ~n20229;
  assign n20231 = n20228 & n20230;
  assign n30199 = n20117 & n20118;
  assign n30200 = (n20028 & n20117) | (n20028 & n30199) | (n20117 & n30199);
  assign n30201 = n20111 | n20113;
  assign n30202 = (n20111 & n30141) | (n20111 & n30201) | (n30141 & n30201);
  assign n20236 = x124 & x152;
  assign n30147 = (n19841 & n20036) | (n19841 & n30146) | (n20036 & n30146);
  assign n30150 = n20049 & n20052;
  assign n30205 = n19894 & n20088;
  assign n35010 = (n20088 & n30150) | (n20088 & n30205) | (n30150 & n30205);
  assign n35011 = (n20052 & n20088) | (n20052 & n30205) | (n20088 & n30205);
  assign n35012 = (n29980 & n35010) | (n29980 & n35011) | (n35010 & n35011);
  assign n37330 = n19893 & n20089;
  assign n37331 = n19892 & n37330;
  assign n35014 = (n20088 & n20089) | (n20088 & n37331) | (n20089 & n37331);
  assign n35015 = (n20089 & n30150) | (n20089 & n35014) | (n30150 & n35014);
  assign n35016 = (n20052 & n20089) | (n20052 & n35014) | (n20089 & n35014);
  assign n35017 = (n29980 & n35015) | (n29980 & n35016) | (n35015 & n35016);
  assign n20242 = ~n35012 & n35017;
  assign n30211 = n20095 | n20242;
  assign n35018 = (n20242 & n30152) | (n20242 & n30211) | (n30152 & n30211);
  assign n35019 = (n20242 & n30153) | (n20242 & n30211) | (n30153 & n30211);
  assign n35020 = (n19838 & n35018) | (n19838 & n35019) | (n35018 & n35019);
  assign n30214 = n19887 | n30061;
  assign n20245 = n20071 & ~n20077;
  assign n20246 = ~n20071 & n20077;
  assign n20247 = n20245 | n20246;
  assign n30155 = n19880 | n30086;
  assign n35023 = n20247 | n30155;
  assign n35024 = n20247 | n34980;
  assign n35025 = (n34922 & n35023) | (n34922 & n35024) | (n35023 & n35024);
  assign n35026 = n20247 & n30155;
  assign n35027 = n20247 & n34980;
  assign n35028 = (n34922 & n35026) | (n34922 & n35027) | (n35026 & n35027);
  assign n30216 = n35025 & ~n35028;
  assign n30217 = n19888 & n30216;
  assign n35029 = n30214 & n30217;
  assign n35021 = n19696 | n19887;
  assign n35022 = n30055 | n35021;
  assign n35030 = n30217 & n35022;
  assign n35031 = (n34853 & n35029) | (n34853 & n35030) | (n35029 & n35030);
  assign n35032 = n20085 & ~n35031;
  assign n35033 = n30172 & n35032;
  assign n30219 = n20088 | n35033;
  assign n35034 = n19894 | n35033;
  assign n35035 = (n20088 & n35033) | (n20088 & n35034) | (n35033 & n35034);
  assign n35036 = (n30150 & n30219) | (n30150 & n35035) | (n30219 & n35035);
  assign n35037 = (n20052 & n30219) | (n20052 & n35035) | (n30219 & n35035);
  assign n35038 = (n29980 & n35036) | (n29980 & n35037) | (n35036 & n35037);
  assign n20263 = x132 & x144;
  assign n20264 = x131 & x145;
  assign n20265 = n20263 | n20264;
  assign n20266 = n20263 & n20264;
  assign n20267 = n20265 & ~n20266;
  assign n20268 = n20063 & n20267;
  assign n35039 = n20062 & n20063;
  assign n35040 = n20267 & n35039;
  assign n35041 = (n20268 & n37317) | (n20268 & n35040) | (n37317 & n35040);
  assign n37332 = (n20268 & n35040) | (n20268 & n37319) | (n35040 & n37319);
  assign n37333 = (n19872 & n20268) | (n19872 & n35040) | (n20268 & n35040);
  assign n37334 = (n30078 & n37332) | (n30078 & n37333) | (n37332 & n37333);
  assign n35043 = (n29868 & n35041) | (n29868 & n37334) | (n35041 & n37334);
  assign n20270 = n20062 | n20267;
  assign n30226 = n20064 | n20270;
  assign n35044 = (n20270 & n37317) | (n20270 & n30226) | (n37317 & n30226);
  assign n35045 = (n20270 & n30226) | (n20270 & n34982) | (n30226 & n34982);
  assign n35046 = (n29868 & n35044) | (n29868 & n35045) | (n35044 & n35045);
  assign n20272 = ~n35043 & n35046;
  assign n20273 = x130 & x146;
  assign n20274 = n20272 & n20273;
  assign n20275 = n20272 | n20273;
  assign n20276 = ~n20274 & n20275;
  assign n30164 = n20074 & n30161;
  assign n35047 = n20064 & n37317;
  assign n37335 = n20064 & n37319;
  assign n37336 = n19872 & n20064;
  assign n37337 = (n30078 & n37335) | (n30078 & n37336) | (n37335 & n37336);
  assign n35049 = (n29868 & n35047) | (n29868 & n37337) | (n35047 & n37337);
  assign n35050 = (n20065 & n20066) | (n20065 & n37317) | (n20066 & n37317);
  assign n37338 = (n20065 & n20066) | (n20065 & n37319) | (n20066 & n37319);
  assign n37735 = n19872 & n20065;
  assign n37736 = (n20064 & n20065) | (n20064 & n37735) | (n20065 & n37735);
  assign n37340 = (n30078 & n37338) | (n30078 & n37736) | (n37338 & n37736);
  assign n35052 = (n29868 & n35050) | (n29868 & n37340) | (n35050 & n37340);
  assign n20260 = ~n35049 & n35052;
  assign n30228 = n20260 & n20276;
  assign n35053 = (n20276 & n30164) | (n20276 & n30228) | (n30164 & n30228);
  assign n35054 = (n20276 & n30165) | (n20276 & n30228) | (n30165 & n30228);
  assign n35055 = (n34922 & n35053) | (n34922 & n35054) | (n35053 & n35054);
  assign n30230 = n20260 | n20276;
  assign n35056 = n30164 | n30230;
  assign n35057 = n30165 | n30230;
  assign n35058 = (n34922 & n35056) | (n34922 & n35057) | (n35056 & n35057);
  assign n20279 = ~n35055 & n35058;
  assign n20280 = x129 & x147;
  assign n20281 = n20279 & n20280;
  assign n20282 = n20279 | n20280;
  assign n20283 = ~n20281 & n20282;
  assign n35059 = n30168 | n30216;
  assign n35060 = (n19888 & n30168) | (n19888 & n35059) | (n30168 & n35059);
  assign n30232 = n20283 & n35060;
  assign n30233 = n20283 & n30168;
  assign n35061 = (n30214 & n30232) | (n30214 & n30233) | (n30232 & n30233);
  assign n35062 = (n30232 & n30233) | (n30232 & n35022) | (n30233 & n35022);
  assign n35063 = (n34853 & n35061) | (n34853 & n35062) | (n35061 & n35062);
  assign n30235 = n20283 | n35060;
  assign n30236 = n20283 | n30168;
  assign n35064 = (n30214 & n30235) | (n30214 & n30236) | (n30235 & n30236);
  assign n35065 = (n30235 & n30236) | (n30235 & n35022) | (n30236 & n35022);
  assign n35066 = (n34853 & n35064) | (n34853 & n35065) | (n35064 & n35065);
  assign n20286 = ~n35063 & n35066;
  assign n20287 = x128 & x148;
  assign n20288 = n20286 & n20287;
  assign n20289 = n20286 | n20287;
  assign n20290 = ~n20288 & n20289;
  assign n20291 = x127 & x149;
  assign n20292 = n20290 & n20291;
  assign n20293 = n20290 | n20291;
  assign n20294 = ~n20292 & n20293;
  assign n20295 = n35038 | n20294;
  assign n20296 = n35038 & n20294;
  assign n20297 = n20295 & ~n20296;
  assign n20298 = x126 & x150;
  assign n20299 = n20297 | n20298;
  assign n20300 = n20297 & n20298;
  assign n20301 = n20299 & ~n20300;
  assign n20302 = ~n35020 & n20301;
  assign n20303 = n35020 & ~n20301;
  assign n20304 = n20302 | n20303;
  assign n20305 = x125 & x151;
  assign n20306 = n20304 & n20305;
  assign n20307 = n20304 | n20305;
  assign n20308 = ~n20306 & n20307;
  assign n30203 = n20099 | n20101;
  assign n35067 = n20308 | n30203;
  assign n35068 = n20099 | n20308;
  assign n35069 = (n30147 & n35067) | (n30147 & n35068) | (n35067 & n35068);
  assign n35070 = n20308 & n30203;
  assign n35071 = n20099 & n20308;
  assign n35072 = (n30147 & n35070) | (n30147 & n35071) | (n35070 & n35071);
  assign n20311 = n35069 & ~n35072;
  assign n30238 = n20105 | n20311;
  assign n35073 = n20107 | n30238;
  assign n35074 = (n30145 & n30238) | (n30145 & n35073) | (n30238 & n35073);
  assign n30240 = n20105 & n20311;
  assign n35075 = (n20107 & n20311) | (n20107 & n30240) | (n20311 & n30240);
  assign n35076 = n20311 & n30240;
  assign n35077 = (n30145 & n35075) | (n30145 & n35076) | (n35075 & n35076);
  assign n20314 = n35074 & ~n35077;
  assign n20315 = n20236 & n20314;
  assign n20316 = n20236 | n20314;
  assign n20317 = ~n20315 & n20316;
  assign n20318 = n30202 & n20317;
  assign n20319 = n30202 | n20317;
  assign n20320 = ~n20318 & n20319;
  assign n20321 = x123 & x153;
  assign n20322 = n20320 | n20321;
  assign n20323 = n20320 & n20321;
  assign n20324 = n20322 & ~n20323;
  assign n20325 = ~n30200 & n20324;
  assign n20326 = n30200 & ~n20324;
  assign n20327 = n20325 | n20326;
  assign n20328 = x122 & x154;
  assign n20329 = x121 & x155;
  assign n20330 = n20328 & n20329;
  assign n20331 = n20328 | n20329;
  assign n20332 = ~n20330 & n20331;
  assign n20333 = n20327 & n20332;
  assign n20334 = n20327 | n20332;
  assign n20335 = ~n20333 & n20334;
  assign n30242 = n20225 & n20226;
  assign n30243 = (n20134 & n20225) | (n20134 & n30242) | (n20225 & n30242);
  assign n20338 = n20335 | n30243;
  assign n20339 = n20335 & n30243;
  assign n20340 = n20338 & ~n20339;
  assign n30244 = n20231 | n20340;
  assign n30245 = n30180 | n30244;
  assign n30246 = n20231 & n20340;
  assign n30247 = (n20340 & n30180) | (n20340 & n30246) | (n30180 & n30246);
  assign n20343 = n30245 & ~n30247;
  assign n20344 = x120 & x156;
  assign n20345 = x119 & x157;
  assign n20346 = n20344 & n20345;
  assign n20347 = n20344 | n20345;
  assign n20348 = ~n20346 & n20347;
  assign n20349 = n20343 & n20348;
  assign n20350 = n20343 | n20348;
  assign n20351 = ~n20349 & n20350;
  assign n20352 = n30198 | n20351;
  assign n20353 = n30198 & n20351;
  assign n20354 = n20352 & ~n20353;
  assign n20355 = x118 & x158;
  assign n20356 = n20354 | n20355;
  assign n20357 = n20354 & n20355;
  assign n20358 = n20356 & ~n20357;
  assign n20360 = n20150 | n20222;
  assign n30248 = n20142 & ~n20222;
  assign n30249 = (n20142 & ~n20150) | (n20142 & n30248) | (~n20150 & n30248);
  assign n20362 = n20360 & n30249;
  assign n30250 = n20153 | n20362;
  assign n30251 = (n20362 & n30184) | (n20362 & n30250) | (n30184 & n30250);
  assign n20364 = ~n20358 & n30251;
  assign n20365 = n20358 & ~n30251;
  assign n20366 = n20364 | n20365;
  assign n20367 = x117 & x159;
  assign n20368 = n20366 & n20367;
  assign n20369 = n20366 | n20367;
  assign n20370 = ~n20368 & n20369;
  assign n20371 = n20153 | n30184;
  assign n30252 = (n20154 & n20155) | (n20154 & ~n30184) | (n20155 & ~n30184);
  assign n20373 = n20371 & n30252;
  assign n30253 = n20162 | n20373;
  assign n30254 = (n20373 & n30186) | (n20373 & n30253) | (n30186 & n30253);
  assign n20375 = ~n20370 & n30254;
  assign n20376 = n20370 & ~n30254;
  assign n20377 = n20375 | n20376;
  assign n20215 = n20162 & n30186;
  assign n30193 = n20162 & n20163;
  assign n30194 = (n20163 & n30186) | (n20163 & n30193) | (n30186 & n30193);
  assign n20218 = ~n20215 & n30194;
  assign n30195 = n20176 | n20218;
  assign n30255 = n20377 & n30195;
  assign n30256 = n20218 & n20377;
  assign n30257 = (n30129 & n30255) | (n30129 & n30256) | (n30255 & n30256);
  assign n30258 = n20377 | n30195;
  assign n30259 = n20218 | n20377;
  assign n30260 = (n30129 & n30258) | (n30129 & n30259) | (n30258 & n30259);
  assign n20380 = ~n30257 & n30260;
  assign n20381 = ~n20214 & n20380;
  assign n20382 = n20214 & ~n20380;
  assign n20383 = n20381 | n20382;
  assign n30261 = n20180 & n20383;
  assign n30262 = (n20183 & n20383) | (n20183 & n30261) | (n20383 & n30261);
  assign n30263 = n20180 | n20383;
  assign n30264 = n20183 | n30263;
  assign n20386 = ~n30262 & n30264;
  assign n20387 = n20212 & n20386;
  assign n20388 = n20212 | n20386;
  assign n20389 = ~n20387 & n20388;
  assign n20390 = n30192 & n20389;
  assign n20391 = n30192 | n20389;
  assign n20392 = ~n20390 & n20391;
  assign n20393 = n20210 | n20392;
  assign n20394 = n20210 & n20392;
  assign n20395 = n20393 & ~n20394;
  assign n20396 = x113 & x163;
  assign n35078 = n20008 | n20199;
  assign n35079 = (n20007 & n20199) | (n20007 & n35078) | (n20199 & n35078);
  assign n30266 = (n20009 & n20198) | (n20009 & n35079) | (n20198 & n35079);
  assign n20398 = n20200 & n30266;
  assign n20399 = n20396 | n20398;
  assign n20400 = n20396 & n20398;
  assign n20401 = n20399 & ~n20400;
  assign n20402 = n20395 & ~n20401;
  assign n20403 = ~n20395 & n20401;
  assign n20404 = n20402 | n20403;
  assign n20405 = ~n20207 & n20404;
  assign n20406 = n20207 & ~n20404;
  assign n20407 = n20405 | n20406;
  assign n20408 = x112 & x164;
  assign n20409 = n20407 & n20408;
  assign n20410 = n20407 | n20408;
  assign n20411 = ~n20409 & n20410;
  assign n20412 = n20394 | n20398;
  assign n20414 = x114 & x163;
  assign n35080 = n20210 & n20414;
  assign n35081 = (n20392 & n20414) | (n20392 & n35080) | (n20414 & n35080);
  assign n30268 = n20412 & n35081;
  assign n35082 = n20210 | n20414;
  assign n35083 = n20392 | n35082;
  assign n30270 = (n20412 & n20414) | (n20412 & n35083) | (n20414 & n35083);
  assign n20417 = ~n30268 & n30270;
  assign n20418 = x115 & x162;
  assign n20419 = n20387 | n20390;
  assign n20420 = x116 & x161;
  assign n20423 = x117 & x160;
  assign n20429 = n20343 & n20344;
  assign n20430 = n20343 | n20344;
  assign n20431 = ~n20429 & n20430;
  assign n30277 = n20429 | n20431;
  assign n30278 = (n20429 & n30198) | (n20429 & n30277) | (n30198 & n30277);
  assign n20434 = n20327 | n20328;
  assign n20435 = n20327 & n20328;
  assign n20436 = n20434 & ~n20435;
  assign n20437 = n30243 & n20436;
  assign n20438 = n30243 | n20436;
  assign n20439 = n20329 & n20438;
  assign n20440 = ~n20437 & n20439;
  assign n20446 = n20100 & n20304;
  assign n30283 = n20099 & n20446;
  assign n30154 = (n19838 & n30152) | (n19838 & n30153) | (n30152 & n30153);
  assign n30288 = n20297 & n30211;
  assign n30289 = n20242 & n20297;
  assign n30290 = (n30154 & n30288) | (n30154 & n30289) | (n30288 & n30289);
  assign n37341 = (n20298 & n20300) | (n20298 & n30211) | (n20300 & n30211);
  assign n37342 = n20242 & n20298;
  assign n37343 = (n20297 & n20298) | (n20297 & n37342) | (n20298 & n37342);
  assign n35086 = (n30154 & n37341) | (n30154 & n37343) | (n37341 & n37343);
  assign n20454 = ~n30290 & n35086;
  assign n20456 = n35038 | n20290;
  assign n35087 = ~n20085 & n35031;
  assign n35088 = (n20085 & n30172) | (n20085 & ~n35087) | (n30172 & ~n35087);
  assign n20460 = n20290 & n35088;
  assign n20457 = n19894 | n35033;
  assign n30294 = n20457 & n20460;
  assign n35089 = (n20460 & n30150) | (n20460 & n30294) | (n30150 & n30294);
  assign n35090 = (n20052 & n20460) | (n20052 & n30294) | (n20460 & n30294);
  assign n35091 = (n29980 & n35089) | (n29980 & n35090) | (n35089 & n35090);
  assign n20462 = n20291 & ~n35091;
  assign n20463 = n20456 & n20462;
  assign n37344 = n20297 | n20463;
  assign n37345 = (n20463 & n30211) | (n20463 & n37344) | (n30211 & n37344);
  assign n35093 = n20463 | n30289;
  assign n35094 = (n30154 & n37345) | (n30154 & n35093) | (n37345 & n35093);
  assign n30215 = (n34853 & n35022) | (n34853 & n30214) | (n35022 & n30214);
  assign n20467 = n19870 | n20264;
  assign n20468 = n19869 & n20467;
  assign n35095 = n19874 | n20468;
  assign n37346 = n20468 | n37311;
  assign n37347 = (n34912 & n35095) | (n34912 & n37346) | (n35095 & n37346);
  assign n20472 = x133 & x144;
  assign n20473 = x132 & x145;
  assign n20474 = n20472 & n20473;
  assign n20475 = n20472 | n20473;
  assign n20476 = ~n20474 & n20475;
  assign n20477 = x131 & x146;
  assign n20478 = n20476 & n20477;
  assign n20479 = n20476 | n20477;
  assign n20480 = ~n20478 & n20479;
  assign n35097 = n20063 | n20266;
  assign n35098 = (n20266 & n20267) | (n20266 & n35097) | (n20267 & n35097);
  assign n30304 = n20480 & ~n35098;
  assign n30305 = ~n20266 & n20480;
  assign n35099 = (~n37347 & n30304) | (~n37347 & n30305) | (n30304 & n30305);
  assign n35096 = (n20468 & n30078) | (n20468 & n35095) | (n30078 & n35095);
  assign n35100 = (n30304 & n30305) | (n30304 & ~n35096) | (n30305 & ~n35096);
  assign n35101 = (~n29868 & n35099) | (~n29868 & n35100) | (n35099 & n35100);
  assign n30307 = ~n20480 & n35098;
  assign n30308 = n20266 & ~n20480;
  assign n35102 = (n37347 & n30307) | (n37347 & n30308) | (n30307 & n30308);
  assign n35103 = (n30307 & n30308) | (n30307 & n35096) | (n30308 & n35096);
  assign n35104 = (n29868 & n35102) | (n29868 & n35103) | (n35102 & n35103);
  assign n20483 = n35101 | n35104;
  assign n30313 = n20260 | n20274;
  assign n35105 = (n20274 & n20276) | (n20274 & n30313) | (n20276 & n30313);
  assign n30310 = n20483 | n35105;
  assign n35106 = n20274 | n20483;
  assign n35107 = n20276 | n35106;
  assign n35108 = (n30164 & n30310) | (n30164 & n35107) | (n30310 & n35107);
  assign n35109 = (n30165 & n30310) | (n30165 & n35107) | (n30310 & n35107);
  assign n35110 = (n34922 & n35108) | (n34922 & n35109) | (n35108 & n35109);
  assign n20486 = n20275 & n20483;
  assign n30315 = n20486 & n30313;
  assign n35111 = (n20486 & n30164) | (n20486 & n30315) | (n30164 & n30315);
  assign n35112 = (n20486 & n30165) | (n20486 & n30315) | (n30165 & n30315);
  assign n35113 = (n34922 & n35111) | (n34922 & n35112) | (n35111 & n35112);
  assign n20488 = n35110 & ~n35113;
  assign n20489 = x130 & x147;
  assign n20490 = n20488 & n20489;
  assign n20491 = n20488 | n20489;
  assign n20492 = ~n20490 & n20491;
  assign n37348 = n20281 | n20492;
  assign n37349 = n30232 | n37348;
  assign n30321 = n20281 | n30168;
  assign n35114 = (n20281 & n20283) | (n20281 & n30321) | (n20283 & n30321);
  assign n35116 = n20492 | n35114;
  assign n35117 = (n30215 & n37349) | (n30215 & n35116) | (n37349 & n35116);
  assign n20505 = x129 & x148;
  assign n30320 = n20281 | n35060;
  assign n20496 = n20483 & ~n20489;
  assign n20497 = ~n20483 & n20489;
  assign n20498 = n20496 | n20497;
  assign n30326 = n20498 & n35105;
  assign n30297 = n20274 | n20276;
  assign n30327 = n20498 & n30297;
  assign n35121 = (n30164 & n30326) | (n30164 & n30327) | (n30326 & n30327);
  assign n35122 = (n30165 & n30326) | (n30165 & n30327) | (n30326 & n30327);
  assign n35123 = (n34922 & n35121) | (n34922 & n35122) | (n35121 & n35122);
  assign n30329 = n20280 & ~n35123;
  assign n30330 = (n20279 & ~n35123) | (n20279 & n30329) | (~n35123 & n30329);
  assign n30323 = n20498 | n35105;
  assign n30324 = n20498 | n30297;
  assign n35118 = (n30164 & n30323) | (n30164 & n30324) | (n30323 & n30324);
  assign n35119 = (n30165 & n30323) | (n30165 & n30324) | (n30323 & n30324);
  assign n35120 = (n34922 & n35118) | (n34922 & n35119) | (n35118 & n35119);
  assign n37737 = n20505 & ~n35120;
  assign n37738 = (n20505 & ~n30330) | (n20505 & n37737) | (~n30330 & n37737);
  assign n37351 = (n20505 & ~n30320) | (n20505 & n37738) | (~n30320 & n37738);
  assign n20502 = n35120 & n30330;
  assign n30332 = n20502 & n30321;
  assign n35125 = n20505 & ~n30332;
  assign n35126 = (~n30215 & n37351) | (~n30215 & n35125) | (n37351 & n35125);
  assign n30335 = n35117 & n35126;
  assign n37739 = ~n20505 & n35120;
  assign n37740 = n30330 & n37739;
  assign n37353 = n30320 & n37740;
  assign n35128 = ~n20505 & n30332;
  assign n35129 = (n30215 & n37353) | (n30215 & n35128) | (n37353 & n35128);
  assign n30337 = (n35117 & n20505) | (n35117 & ~n35129) | (n20505 & ~n35129);
  assign n20508 = ~n30335 & n30337;
  assign n20509 = x128 & x149;
  assign n20510 = n20508 & n20509;
  assign n20511 = n20508 | n20509;
  assign n20512 = ~n20510 & n20511;
  assign n30338 = ~n20288 & n20512;
  assign n30339 = ~n35091 & n30338;
  assign n30340 = n20288 & ~n20512;
  assign n30341 = (~n20512 & n35091) | (~n20512 & n30340) | (n35091 & n30340);
  assign n20515 = n30339 | n30341;
  assign n20516 = x127 & x150;
  assign n20517 = n20515 & n20516;
  assign n20518 = n20515 | n20516;
  assign n20519 = ~n20517 & n20518;
  assign n20520 = x126 & x151;
  assign n20521 = ~n20519 & n20520;
  assign n20522 = n20519 & ~n20520;
  assign n20523 = n20521 | n20522;
  assign n20524 = n35094 | n20523;
  assign n20525 = n35094 & n20523;
  assign n20526 = n20524 & ~n20525;
  assign n30342 = ~n20454 & n20526;
  assign n35130 = ~n30283 & n30342;
  assign n35131 = ~n20446 & n30342;
  assign n35132 = (~n30147 & n35130) | (~n30147 & n35131) | (n35130 & n35131);
  assign n30344 = n20454 & ~n20526;
  assign n35133 = (~n20526 & n30283) | (~n20526 & n30344) | (n30283 & n30344);
  assign n35134 = (n20446 & ~n20526) | (n20446 & n30344) | (~n20526 & n30344);
  assign n35135 = (n30147 & n35133) | (n30147 & n35134) | (n35133 & n35134);
  assign n20529 = n35132 | n35135;
  assign n20530 = x125 & x152;
  assign n20531 = n20529 & n20530;
  assign n20532 = n20529 | n20530;
  assign n20533 = ~n20531 & n20532;
  assign n20443 = n20099 | n20304;
  assign n30281 = n20101 | n20443;
  assign n30282 = (n20443 & n30147) | (n20443 & n30281) | (n30147 & n30281);
  assign n30284 = (n20446 & n30147) | (n20446 & n30283) | (n30147 & n30283);
  assign n20448 = n30282 & ~n30284;
  assign n20449 = n20305 & n20448;
  assign n30286 = n20311 | n20449;
  assign n35136 = n20533 | n30286;
  assign n30285 = n20449 | n30240;
  assign n35137 = n20533 | n30285;
  assign n35138 = (n20108 & n35136) | (n20108 & n35137) | (n35136 & n35137);
  assign n35139 = n20533 & n30286;
  assign n35140 = n20533 & n30285;
  assign n35141 = (n20108 & n35139) | (n20108 & n35140) | (n35139 & n35140);
  assign n20536 = n35138 & ~n35141;
  assign n35143 = n20315 | n20536;
  assign n37354 = n20317 | n35143;
  assign n35144 = (n30202 & n37354) | (n30202 & n35143) | (n37354 & n35143);
  assign n35146 = n20315 & n20536;
  assign n37355 = (n20317 & n20536) | (n20317 & n35146) | (n20536 & n35146);
  assign n35147 = (n30202 & n37355) | (n30202 & n35146) | (n37355 & n35146);
  assign n20539 = n35144 & ~n35147;
  assign n20540 = x124 & x153;
  assign n20541 = x123 & x154;
  assign n20542 = n20540 & n20541;
  assign n20543 = n20540 | n20541;
  assign n20544 = ~n20542 & n20543;
  assign n20545 = n20539 & n20544;
  assign n20546 = n20539 | n20544;
  assign n20547 = ~n20545 & n20546;
  assign n30346 = n20322 & n20323;
  assign n30347 = (n20322 & n30200) | (n20322 & n30346) | (n30200 & n30346);
  assign n20550 = n20547 | n30347;
  assign n20551 = n20547 & n30347;
  assign n20552 = n20550 & ~n20551;
  assign n20553 = x122 & x155;
  assign n20554 = n20552 | n20553;
  assign n20555 = n20552 & n20553;
  assign n20556 = n20554 & ~n20555;
  assign n30348 = n20434 & n20435;
  assign n30349 = (n20434 & n30243) | (n20434 & n30348) | (n30243 & n30348);
  assign n20559 = n20556 | n30349;
  assign n20560 = n20556 & n30349;
  assign n20561 = n20559 & ~n20560;
  assign n30350 = n20440 | n20561;
  assign n30351 = n30247 | n30350;
  assign n30352 = n20440 & n20561;
  assign n30353 = (n20561 & n30247) | (n20561 & n30352) | (n30247 & n30352);
  assign n20564 = n30351 & ~n30353;
  assign n20565 = x121 & x156;
  assign n20566 = x120 & x157;
  assign n20567 = n20565 & n20566;
  assign n20568 = n20565 | n20566;
  assign n20569 = ~n20567 & n20568;
  assign n20570 = n20564 & n20569;
  assign n20571 = n20564 | n20569;
  assign n20572 = ~n20570 & n20571;
  assign n20573 = n30278 | n20572;
  assign n20574 = n30278 & n20572;
  assign n20575 = n20573 & ~n20574;
  assign n20576 = x119 & x158;
  assign n20577 = n20575 | n20576;
  assign n20578 = n20575 & n20576;
  assign n20579 = n20577 & ~n20578;
  assign n30354 = n20354 & n30250;
  assign n30355 = n20354 & n20362;
  assign n30356 = (n30184 & n30354) | (n30184 & n30355) | (n30354 & n30355);
  assign n20581 = n30198 | n20431;
  assign n30357 = n20345 & ~n20431;
  assign n30358 = (n20345 & ~n30198) | (n20345 & n30357) | (~n30198 & n30357);
  assign n20583 = n20581 & n30358;
  assign n20584 = n30356 | n20583;
  assign n20585 = ~n20579 & n20584;
  assign n20586 = n20579 & ~n20584;
  assign n20587 = n20585 | n20586;
  assign n20588 = x118 & x159;
  assign n20589 = n20587 & n20588;
  assign n20590 = n20587 | n20588;
  assign n20591 = ~n20589 & n20590;
  assign n30274 = n20366 & n30253;
  assign n30275 = n20366 & n20373;
  assign n30276 = (n30186 & n30274) | (n30186 & n30275) | (n30274 & n30275);
  assign n30359 = n20354 | n30250;
  assign n30360 = n20354 | n20362;
  assign n30361 = (n30184 & n30359) | (n30184 & n30360) | (n30359 & n30360);
  assign n20593 = n20355 & ~n30356;
  assign n20594 = n30361 & n20593;
  assign n20595 = n30276 | n20594;
  assign n20596 = ~n20591 & n20595;
  assign n20597 = n20591 & ~n20595;
  assign n20598 = n20596 | n20597;
  assign n30271 = n20366 | n30253;
  assign n30272 = n20366 | n20373;
  assign n30273 = (n30186 & n30271) | (n30186 & n30272) | (n30271 & n30272);
  assign n20426 = n20367 & ~n30276;
  assign n20427 = n30273 & n20426;
  assign n30362 = n20427 & n20598;
  assign n30363 = (n20598 & n30257) | (n20598 & n30362) | (n30257 & n30362);
  assign n30364 = n20427 | n20598;
  assign n30365 = n30257 | n30364;
  assign n20601 = ~n30363 & n30365;
  assign n20602 = ~n20423 & n20601;
  assign n20603 = n20423 & ~n20601;
  assign n20604 = n20602 | n20603;
  assign n20421 = n20214 & n20380;
  assign n30366 = n20421 & n20604;
  assign n30367 = (n20604 & n30262) | (n20604 & n30366) | (n30262 & n30366);
  assign n30368 = n20421 | n20604;
  assign n30369 = n30262 | n30368;
  assign n20607 = ~n30367 & n30369;
  assign n20608 = n20420 & n20607;
  assign n20609 = n20420 | n20607;
  assign n20610 = ~n20608 & n20609;
  assign n20611 = n20419 & n20610;
  assign n20612 = n20419 | n20610;
  assign n20613 = ~n20611 & n20612;
  assign n20614 = n20418 | n20613;
  assign n20615 = n20418 & n20613;
  assign n20616 = n20614 & ~n20615;
  assign n20617 = ~n20417 & n20616;
  assign n20618 = n20417 & ~n20616;
  assign n20619 = n20617 | n20618;
  assign n30370 = n20206 & n20396;
  assign n30371 = n20205 & n30370;
  assign n20621 = n20395 & ~n20398;
  assign n20622 = ~n20395 & n20398;
  assign n20623 = n20621 | n20622;
  assign n20624 = n30371 | n20623;
  assign n30372 = n20206 | n20396;
  assign n30373 = (n20205 & n20396) | (n20205 & n30372) | (n20396 & n30372);
  assign n20626 = n20624 & n30373;
  assign n20627 = n20619 & ~n20626;
  assign n20628 = ~n20619 & n20626;
  assign n20629 = n20627 | n20628;
  assign n20630 = x113 & x164;
  assign n20631 = n20629 & ~n20630;
  assign n20632 = ~n20629 & n20630;
  assign n20633 = n20631 | n20632;
  assign n20634 = ~n20409 & n20633;
  assign n20635 = n20409 & ~n20633;
  assign n20636 = n20634 | n20635;
  assign n20637 = x112 & x165;
  assign n20638 = n20636 & n20637;
  assign n20639 = n20636 | n20637;
  assign n20640 = ~n20638 & n20639;
  assign n20641 = x116 & x162;
  assign n30374 = n20608 | n20610;
  assign n30375 = (n20419 & n20608) | (n20419 & n30374) | (n20608 & n30374);
  assign n20643 = x117 & x161;
  assign n20646 = x118 & x160;
  assign n20652 = n20564 & n20565;
  assign n20653 = n20564 | n20565;
  assign n20654 = ~n20652 & n20653;
  assign n30380 = n20652 | n20654;
  assign n30381 = (n20652 & n30278) | (n20652 & n30380) | (n30278 & n30380);
  assign n20657 = n20552 & n30349;
  assign n30382 = (n20553 & n20555) | (n20553 & n30349) | (n20555 & n30349);
  assign n20660 = ~n20657 & n30382;
  assign n37356 = n20311 | n20529;
  assign n37357 = n20449 | n37356;
  assign n35149 = n20529 | n30285;
  assign n35150 = (n20108 & n37357) | (n20108 & n35149) | (n37357 & n35149);
  assign n20665 = n20305 | n20448;
  assign n20666 = n20529 & n20665;
  assign n20663 = n20105 | n20449;
  assign n30383 = n20663 & n20666;
  assign n30384 = (n20108 & n20666) | (n20108 & n30383) | (n20666 & n30383);
  assign n20668 = n20530 & ~n30384;
  assign n20669 = n35150 & n20668;
  assign n30279 = n20315 | n20317;
  assign n30385 = n20536 | n20669;
  assign n35151 = (n20669 & n30279) | (n20669 & n30385) | (n30279 & n30385);
  assign n35152 = (n20315 & n20669) | (n20315 & n30385) | (n20669 & n30385);
  assign n35153 = (n30202 & n35151) | (n30202 & n35152) | (n35151 & n35152);
  assign n30402 = n20288 & n20508;
  assign n30403 = (n20508 & n35091) | (n20508 & n30402) | (n35091 & n30402);
  assign n37358 = n20287 & n20509;
  assign n37359 = n20286 & n37358;
  assign n35161 = (n20508 & n20509) | (n20508 & n37359) | (n20509 & n37359);
  assign n30407 = (n20509 & n35091) | (n20509 & n35161) | (n35091 & n35161);
  assign n20688 = ~n30403 & n30407;
  assign n20676 = n20242 | n20463;
  assign n30395 = n20095 | n20676;
  assign n30397 = ~n20291 & n35091;
  assign n30398 = (n20291 & n20456) | (n20291 & ~n30397) | (n20456 & ~n30397);
  assign n20680 = n20515 & n30398;
  assign n30408 = n20680 | n20688;
  assign n35162 = (n20688 & n30395) | (n20688 & n30408) | (n30395 & n30408);
  assign n35163 = (n20676 & n20688) | (n20676 & n30408) | (n20688 & n30408);
  assign n35164 = (n30154 & n35162) | (n30154 & n35163) | (n35162 & n35163);
  assign n20697 = x134 & x144;
  assign n20698 = x133 & x145;
  assign n20699 = n20697 | n20698;
  assign n20700 = n20697 & n20698;
  assign n20701 = n20699 & ~n20700;
  assign n20702 = n20474 | n20701;
  assign n30413 = n20476 & n35098;
  assign n30425 = n20702 | n30413;
  assign n30414 = n20266 & n20476;
  assign n30426 = n20702 | n30414;
  assign n35166 = (n37347 & n30425) | (n37347 & n30426) | (n30425 & n30426);
  assign n35167 = (n30425 & n30426) | (n30425 & n35096) | (n30426 & n35096);
  assign n35168 = (n29868 & n35166) | (n29868 & n35167) | (n35166 & n35167);
  assign n20706 = n20475 & n20701;
  assign n20704 = n20266 | n20474;
  assign n30428 = n20268 | n20704;
  assign n30430 = n20706 & n30428;
  assign n30431 = n20704 & n20706;
  assign n35169 = (n37347 & n30430) | (n37347 & n30431) | (n30430 & n30431);
  assign n35170 = (n30430 & n30431) | (n30430 & n35096) | (n30431 & n35096);
  assign n35171 = (n29868 & n35169) | (n29868 & n35170) | (n35169 & n35170);
  assign n20708 = n35168 & ~n35171;
  assign n20709 = x132 & x146;
  assign n20710 = n20708 & n20709;
  assign n20711 = n20708 | n20709;
  assign n20712 = ~n20710 & n20711;
  assign n35172 = (n37347 & n30413) | (n37347 & n30414) | (n30413 & n30414);
  assign n35173 = (n30413 & n30414) | (n30413 & n35096) | (n30414 & n35096);
  assign n35174 = (n29868 & n35172) | (n29868 & n35173) | (n35172 & n35173);
  assign n35175 = (n20477 & n20478) | (n20477 & n35098) | (n20478 & n35098);
  assign n35176 = n20266 & n20477;
  assign n35177 = (n20476 & n20477) | (n20476 & n35176) | (n20477 & n35176);
  assign n35178 = (n37347 & n35175) | (n37347 & n35177) | (n35175 & n35177);
  assign n35179 = (n35096 & n35175) | (n35096 & n35177) | (n35175 & n35177);
  assign n35180 = (n29868 & n35178) | (n29868 & n35179) | (n35178 & n35179);
  assign n20695 = ~n35174 & n35180;
  assign n35183 = n20483 | n20695;
  assign n35184 = (n20275 & n20695) | (n20275 & n35183) | (n20695 & n35183);
  assign n30434 = n20712 & n35184;
  assign n35181 = n20695 & n20712;
  assign n35182 = (n20712 & n30315) | (n20712 & n35181) | (n30315 & n35181);
  assign n35185 = (n30164 & n30434) | (n30164 & n35182) | (n30434 & n35182);
  assign n35186 = (n30165 & n30434) | (n30165 & n35182) | (n30434 & n35182);
  assign n35187 = (n34922 & n35185) | (n34922 & n35186) | (n35185 & n35186);
  assign n30437 = n20712 | n35184;
  assign n35188 = n20695 | n20712;
  assign n35189 = n30315 | n35188;
  assign n35190 = (n30164 & n30437) | (n30164 & n35189) | (n30437 & n35189);
  assign n35191 = (n30165 & n30437) | (n30165 & n35189) | (n30437 & n35189);
  assign n35192 = (n34922 & n35190) | (n34922 & n35191) | (n35190 & n35191);
  assign n20715 = ~n35187 & n35192;
  assign n20716 = x131 & x147;
  assign n20717 = n20715 & n20716;
  assign n20718 = n20715 | n20716;
  assign n20719 = ~n20717 & n20718;
  assign n30331 = n20502 & n30320;
  assign n30439 = n20490 & n20719;
  assign n35193 = (n20719 & n30331) | (n20719 & n30439) | (n30331 & n30439);
  assign n35194 = (n20719 & n30332) | (n20719 & n30439) | (n30332 & n30439);
  assign n35195 = (n30215 & n35193) | (n30215 & n35194) | (n35193 & n35194);
  assign n30441 = n20490 | n20719;
  assign n35196 = n30331 | n30441;
  assign n35197 = n30332 | n30441;
  assign n35198 = (n30215 & n35196) | (n30215 & n35197) | (n35196 & n35197);
  assign n20722 = ~n35195 & n35198;
  assign n20723 = x130 & x148;
  assign n20724 = n20722 & n20723;
  assign n20725 = n20722 | n20723;
  assign n20726 = ~n20724 & n20725;
  assign n20727 = x129 & x149;
  assign n20728 = n20726 & n20727;
  assign n20729 = n20726 | n20727;
  assign n20730 = ~n20728 & n20729;
  assign n30411 = n20508 | n30335;
  assign n35199 = n20730 | n30411;
  assign n30528 = n20288 | n30335;
  assign n35165 = (n20508 & n30335) | (n20508 & n30528) | (n30335 & n30528);
  assign n35200 = n20730 | n35165;
  assign n35201 = (n35091 & n35199) | (n35091 & n35200) | (n35199 & n35200);
  assign n35202 = n20730 & n30411;
  assign n35203 = n20730 & n35165;
  assign n35204 = (n35091 & n35202) | (n35091 & n35203) | (n35202 & n35203);
  assign n20733 = n35201 & ~n35204;
  assign n20734 = x128 & x150;
  assign n20735 = n20733 | n20734;
  assign n20736 = n20733 & n20734;
  assign n20737 = n20735 & ~n20736;
  assign n20738 = ~n35164 & n20737;
  assign n20739 = n35164 & ~n20737;
  assign n20740 = n20738 | n20739;
  assign n20741 = x127 & x151;
  assign n20742 = n20740 & n20741;
  assign n20743 = n20740 | n20741;
  assign n20744 = ~n20742 & n20743;
  assign n30393 = n20463 | n20515;
  assign n35154 = n30288 | n30393;
  assign n35155 = n30289 | n30393;
  assign n35156 = (n30154 & n35154) | (n30154 & n35155) | (n35154 & n35155);
  assign n35157 = n20680 & n30395;
  assign n35158 = n20676 & n20680;
  assign n35159 = (n30154 & n35157) | (n30154 & n35158) | (n35157 & n35158);
  assign n20682 = n35156 & ~n35159;
  assign n20683 = n20516 & n20682;
  assign n30387 = n20463 | n20519;
  assign n30388 = n30290 | n30387;
  assign n30389 = n20463 & n20519;
  assign n30390 = (n20519 & n30290) | (n20519 & n30389) | (n30290 & n30389);
  assign n20673 = n30388 & ~n30390;
  assign n30391 = n20454 & n20673;
  assign n30399 = n20683 | n30391;
  assign n35205 = n20744 | n30399;
  assign n30400 = n20673 | n20683;
  assign n35206 = n20744 | n30400;
  assign n35207 = (n30284 & n35205) | (n30284 & n35206) | (n35205 & n35206);
  assign n35208 = n20744 & n30399;
  assign n35209 = n20744 & n30400;
  assign n35210 = (n30284 & n35208) | (n30284 & n35209) | (n35208 & n35209);
  assign n20747 = n35207 & ~n35210;
  assign n20748 = x126 & x152;
  assign n20749 = n20747 | n20748;
  assign n20750 = n20747 & n20748;
  assign n20751 = n20749 & ~n20750;
  assign n30443 = n20454 | n20673;
  assign n35211 = n30283 | n30443;
  assign n35212 = n20446 | n30443;
  assign n35213 = (n30147 & n35211) | (n30147 & n35212) | (n35211 & n35212);
  assign n30446 = n20520 & ~n20673;
  assign n35214 = ~n20454 & n20520;
  assign n35215 = (n20520 & ~n20673) | (n20520 & n35214) | (~n20673 & n35214);
  assign n35216 = (~n30283 & n30446) | (~n30283 & n35215) | (n30446 & n35215);
  assign n35217 = (~n20446 & n30446) | (~n20446 & n35215) | (n30446 & n35215);
  assign n35218 = (~n30147 & n35216) | (~n30147 & n35217) | (n35216 & n35217);
  assign n20754 = n35213 & n35218;
  assign n35219 = ~n20751 & n20754;
  assign n35220 = (~n20751 & n30384) | (~n20751 & n35219) | (n30384 & n35219);
  assign n35221 = n20751 & ~n20754;
  assign n35222 = ~n30384 & n35221;
  assign n20758 = n35220 | n35222;
  assign n20759 = x125 & x153;
  assign n20760 = n20758 & n20759;
  assign n20761 = n20758 | n20759;
  assign n20762 = ~n20760 & n20761;
  assign n20763 = n35153 | n20762;
  assign n20764 = n35153 & n20762;
  assign n20765 = n20763 & ~n20764;
  assign n20766 = x124 & x154;
  assign n20767 = n20765 | n20766;
  assign n20768 = n20765 & n20766;
  assign n20769 = n20767 & ~n20768;
  assign n20770 = n20539 | n20540;
  assign n20771 = n20539 & n20540;
  assign n30448 = n20770 & n20771;
  assign n30449 = (n20770 & n30347) | (n20770 & n30448) | (n30347 & n30448);
  assign n20774 = n20769 | n30449;
  assign n20775 = n20769 & n30449;
  assign n20776 = n20774 & ~n20775;
  assign n20777 = x123 & x155;
  assign n20778 = n20776 | n20777;
  assign n20779 = n20776 & n20777;
  assign n20780 = n20778 & ~n20779;
  assign n20781 = n20770 & ~n20771;
  assign n20782 = n30347 & n20781;
  assign n35223 = n20541 & n20781;
  assign n35224 = (n20541 & n30347) | (n20541 & n35223) | (n30347 & n35223);
  assign n20785 = ~n20782 & n35224;
  assign n30450 = n20552 | n20785;
  assign n30451 = (n20785 & n30349) | (n20785 & n30450) | (n30349 & n30450);
  assign n20787 = n20780 | n30451;
  assign n20788 = n20780 & n30451;
  assign n20789 = n20787 & ~n20788;
  assign n30452 = n20660 | n20789;
  assign n30453 = n30353 | n30452;
  assign n30454 = n20660 & n20789;
  assign n30455 = (n20789 & n30353) | (n20789 & n30454) | (n30353 & n30454);
  assign n20792 = n30453 & ~n30455;
  assign n20793 = x122 & x156;
  assign n20794 = x121 & x157;
  assign n20795 = n20793 & n20794;
  assign n20796 = n20793 | n20794;
  assign n20797 = ~n20795 & n20796;
  assign n20798 = n20792 & n20797;
  assign n20799 = n20792 | n20797;
  assign n20800 = ~n20798 & n20799;
  assign n20801 = n30381 | n20800;
  assign n20802 = n30381 & n20800;
  assign n20803 = n20801 & ~n20802;
  assign n20804 = x120 & x158;
  assign n20805 = n20803 | n20804;
  assign n20806 = n20803 & n20804;
  assign n20807 = n20805 & ~n20806;
  assign n30456 = n20575 & n20583;
  assign n30457 = (n20575 & n30356) | (n20575 & n30456) | (n30356 & n30456);
  assign n20809 = n30278 | n20654;
  assign n30458 = n20566 & ~n20654;
  assign n30459 = (n20566 & ~n30278) | (n20566 & n30458) | (~n30278 & n30458);
  assign n20811 = n20809 & n30459;
  assign n20812 = n30457 | n20811;
  assign n20813 = ~n20807 & n20812;
  assign n20814 = n20807 & ~n20812;
  assign n20815 = n20813 | n20814;
  assign n20816 = x119 & x159;
  assign n20817 = n20815 & n20816;
  assign n20818 = n20815 | n20816;
  assign n20819 = ~n20817 & n20818;
  assign n30378 = n20587 & n20594;
  assign n30379 = (n20587 & n30276) | (n20587 & n30378) | (n30276 & n30378);
  assign n30460 = n20575 | n20583;
  assign n30461 = n30356 | n30460;
  assign n20821 = n20576 & ~n30457;
  assign n20822 = n30461 & n20821;
  assign n20823 = n30379 | n20822;
  assign n20824 = ~n20819 & n20823;
  assign n20825 = n20819 & ~n20823;
  assign n20826 = n20824 | n20825;
  assign n30376 = n20587 | n20594;
  assign n30377 = n30276 | n30376;
  assign n20649 = n20588 & ~n30379;
  assign n20650 = n30377 & n20649;
  assign n30462 = n20650 & n20826;
  assign n30463 = (n20826 & n30363) | (n20826 & n30462) | (n30363 & n30462);
  assign n30464 = n20650 | n20826;
  assign n30465 = n30363 | n30464;
  assign n20829 = ~n30463 & n30465;
  assign n20830 = ~n20646 & n20829;
  assign n20831 = n20646 & ~n20829;
  assign n20832 = n20830 | n20831;
  assign n20644 = n20423 & n20601;
  assign n30466 = n20644 & n20832;
  assign n30467 = (n20832 & n30367) | (n20832 & n30466) | (n30367 & n30466);
  assign n30468 = n20644 | n20832;
  assign n30469 = n30367 | n30468;
  assign n20835 = ~n30467 & n30469;
  assign n20836 = n20643 & n20835;
  assign n20837 = n20643 | n20835;
  assign n20838 = ~n20836 & n20837;
  assign n20839 = n30375 & n20838;
  assign n20840 = n30375 | n20838;
  assign n20841 = ~n20839 & n20840;
  assign n20842 = n20641 | n20841;
  assign n20843 = n20641 & n20841;
  assign n20844 = n20842 & ~n20843;
  assign n20413 = n20393 & n20412;
  assign n20845 = n20413 | n20615;
  assign n20846 = n20614 & n20845;
  assign n20847 = n20844 & ~n20846;
  assign n20848 = ~n20844 & n20846;
  assign n20849 = n20847 | n20848;
  assign n20850 = x115 & x163;
  assign n20851 = n20849 | n20850;
  assign n20852 = n20849 & n20850;
  assign n20853 = n20851 & ~n20852;
  assign n20854 = ~n20413 & n20616;
  assign n20855 = n20413 & ~n20616;
  assign n20856 = n20854 | n20855;
  assign n20857 = n20414 & n20856;
  assign n20858 = n20626 | n20857;
  assign n20859 = n20414 | n20856;
  assign n20860 = n20858 & n20859;
  assign n20861 = n20853 & ~n20860;
  assign n20862 = ~n20853 & n20860;
  assign n20863 = n20861 | n20862;
  assign n20864 = x114 & x164;
  assign n20865 = n20863 & ~n20864;
  assign n20866 = ~n20863 & n20864;
  assign n20867 = n20865 | n20866;
  assign n30470 = n20408 & n20630;
  assign n30471 = n20407 & n30470;
  assign n20869 = n20629 | n30471;
  assign n20872 = x113 & x165;
  assign n30472 = n20408 | n20630;
  assign n35225 = n20872 & n30472;
  assign n35226 = n20630 & n20872;
  assign n35227 = (n20407 & n35225) | (n20407 & n35226) | (n35225 & n35226);
  assign n30475 = n20869 & n35227;
  assign n35228 = n20872 | n30472;
  assign n35229 = n20630 | n20872;
  assign n35230 = (n20407 & n35228) | (n20407 & n35229) | (n35228 & n35229);
  assign n30477 = (n20869 & n20872) | (n20869 & n35230) | (n20872 & n35230);
  assign n20875 = ~n30475 & n30477;
  assign n20876 = n20867 & ~n20875;
  assign n20877 = ~n20867 & n20875;
  assign n20878 = n20876 | n20877;
  assign n20879 = ~n20638 & n20878;
  assign n20880 = n20638 & ~n20878;
  assign n20881 = n20879 | n20880;
  assign n20882 = x112 & x166;
  assign n20883 = n20881 & n20882;
  assign n20884 = n20881 | n20882;
  assign n20885 = ~n20883 & n20884;
  assign n30478 = n20842 & n20843;
  assign n30479 = (n20842 & n20846) | (n20842 & n30478) | (n20846 & n30478);
  assign n20888 = x116 & x163;
  assign n20889 = n30479 & n20888;
  assign n20890 = n30479 | n20888;
  assign n20891 = ~n20889 & n20890;
  assign n20892 = x117 & x162;
  assign n30480 = n20836 | n20838;
  assign n30481 = (n20836 & n30375) | (n20836 & n30480) | (n30375 & n30480);
  assign n20894 = x118 & x161;
  assign n20897 = x119 & x160;
  assign n20903 = n20792 & n20793;
  assign n20904 = n20792 | n20793;
  assign n20905 = ~n20903 & n20904;
  assign n30486 = n20903 | n20905;
  assign n30487 = (n20903 & n30381) | (n20903 & n30486) | (n30381 & n30486);
  assign n35231 = n20776 & n30450;
  assign n35232 = n20776 & n20785;
  assign n35233 = (n30349 & n35231) | (n30349 & n35232) | (n35231 & n35232);
  assign n30488 = (n20777 & n20779) | (n20777 & n30451) | (n20779 & n30451);
  assign n20911 = ~n35233 & n30488;
  assign n35234 = n20765 & n30448;
  assign n35235 = n20765 & n20770;
  assign n35236 = (n30347 & n35234) | (n30347 & n35235) | (n35234 & n35235);
  assign n35237 = (n20766 & n20768) | (n20766 & n30448) | (n20768 & n30448);
  assign n35238 = (n20766 & n20768) | (n20766 & n20770) | (n20768 & n20770);
  assign n35239 = (n30347 & n35237) | (n30347 & n35238) | (n35237 & n35238);
  assign n20916 = ~n35236 & n35239;
  assign n30490 = n20776 | n20916;
  assign n30491 = (n20916 & n30451) | (n20916 & n30490) | (n30451 & n30490);
  assign n20918 = n20315 | n20669;
  assign n30492 = n20317 | n20918;
  assign n30493 = (n20918 & n30202) | (n20918 & n30492) | (n30202 & n30492);
  assign n30494 = ~n20530 & n30384;
  assign n30495 = (n20530 & n35150) | (n20530 & ~n30494) | (n35150 & ~n30494);
  assign n20922 = n20758 & n30495;
  assign n20923 = n30493 & n20922;
  assign n30280 = (n20315 & n30202) | (n20315 & n30279) | (n30202 & n30279);
  assign n30496 = n20758 | n30385;
  assign n30497 = n20669 | n20758;
  assign n30498 = (n30280 & n30496) | (n30280 & n30497) | (n30496 & n30497);
  assign n20925 = ~n20923 & n30498;
  assign n20926 = n20759 & n20925;
  assign n30499 = n20765 | n20926;
  assign n30500 = (n20926 & n30449) | (n20926 & n30499) | (n30449 & n30499);
  assign n30501 = n20747 & n20754;
  assign n30502 = (n20747 & n30384) | (n20747 & n30501) | (n30384 & n30501);
  assign n35240 = n20748 & n20754;
  assign n35241 = (n20747 & n20748) | (n20747 & n35240) | (n20748 & n35240);
  assign n30506 = (n20748 & n30384) | (n20748 & n35241) | (n30384 & n35241);
  assign n20931 = ~n30502 & n30506;
  assign n30507 = n20922 | n20931;
  assign n30508 = (n20931 & n30493) | (n20931 & n30507) | (n30493 & n30507);
  assign n30509 = n20740 | n30400;
  assign n35242 = n20683 | n20740;
  assign n35243 = n30391 | n35242;
  assign n30511 = (n30284 & n30509) | (n30284 & n35243) | (n30509 & n35243);
  assign n20935 = n20516 | n20682;
  assign n20936 = n20740 & n20935;
  assign n30512 = n20454 | n20683;
  assign n30514 = n20936 & n30512;
  assign n30515 = (n20936 & n30284) | (n20936 & n30514) | (n30284 & n30514);
  assign n20938 = n30511 & ~n30515;
  assign n20939 = n20741 & n20938;
  assign n30516 = n20939 | n30501;
  assign n30517 = n20747 | n20939;
  assign n30518 = (n30384 & n30516) | (n30384 & n30517) | (n30516 & n30517);
  assign n30520 = n20688 & n20733;
  assign n35244 = (n20680 & n20733) | (n20680 & n30520) | (n20733 & n30520);
  assign n35245 = (n30395 & n30520) | (n30395 & n35244) | (n30520 & n35244);
  assign n35246 = (n20676 & n30520) | (n20676 & n35244) | (n30520 & n35244);
  assign n35247 = (n30154 & n35245) | (n30154 & n35246) | (n35245 & n35246);
  assign n30523 = n20688 | n20733;
  assign n35248 = n20680 | n30523;
  assign n35249 = (n30395 & n30523) | (n30395 & n35248) | (n30523 & n35248);
  assign n35250 = (n20676 & n30523) | (n20676 & n35248) | (n30523 & n35248);
  assign n35251 = (n30154 & n35249) | (n30154 & n35250) | (n35249 & n35250);
  assign n20943 = n20734 & n35251;
  assign n20944 = ~n35247 & n20943;
  assign n20946 = n30335 | n20726;
  assign n30525 = n20946 | n30402;
  assign n35252 = n20726 | n30411;
  assign n30527 = (n35091 & n30525) | (n35091 & n35252) | (n30525 & n35252);
  assign n20949 = n30337 & n20726;
  assign n35253 = n30337 & n30528;
  assign n35254 = n20726 & n35253;
  assign n30531 = (n20949 & n35091) | (n20949 & n35254) | (n35091 & n35254);
  assign n20951 = n30527 & ~n30531;
  assign n20952 = n20727 & n20951;
  assign n20957 = x135 & x144;
  assign n20958 = x134 & x145;
  assign n20959 = n20957 & n20958;
  assign n20960 = n20957 | n20958;
  assign n20961 = ~n20959 & n20960;
  assign n20962 = x133 & x146;
  assign n20963 = n20961 & n20962;
  assign n20964 = n20961 | n20962;
  assign n20965 = ~n20963 & n20964;
  assign n37360 = n20475 | n20700;
  assign n37361 = (n20700 & n20701) | (n20700 & n37360) | (n20701 & n37360);
  assign n35256 = (n20700 & n30428) | (n20700 & n37361) | (n30428 & n37361);
  assign n30535 = n20965 & ~n35256;
  assign n35257 = n20700 | n20704;
  assign n35258 = (n20700 & n20706) | (n20700 & n35257) | (n20706 & n35257);
  assign n30536 = n20965 & ~n35258;
  assign n35259 = (~n37347 & n30535) | (~n37347 & n30536) | (n30535 & n30536);
  assign n35260 = (n30535 & n30536) | (n30535 & ~n35096) | (n30536 & ~n35096);
  assign n35261 = (~n29868 & n35259) | (~n29868 & n35260) | (n35259 & n35260);
  assign n30538 = ~n20965 & n35256;
  assign n30539 = ~n20965 & n35258;
  assign n35262 = (n37347 & n30538) | (n37347 & n30539) | (n30538 & n30539);
  assign n35263 = (n30538 & n30539) | (n30538 & n35096) | (n30539 & n35096);
  assign n35264 = (n29868 & n35262) | (n29868 & n35263) | (n35262 & n35263);
  assign n20968 = n35261 | n35264;
  assign n30541 = n20710 | n20968;
  assign n30542 = n35187 | n30541;
  assign n20975 = x132 & x147;
  assign n20972 = n20711 & n20968;
  assign n20970 = n20695 | n20710;
  assign n30544 = n20486 | n20970;
  assign n30547 = n20972 & n30544;
  assign n35265 = n20970 & n20972;
  assign n35266 = (n20972 & n30315) | (n20972 & n35265) | (n30315 & n35265);
  assign n35267 = (n30164 & n30547) | (n30164 & n35266) | (n30547 & n35266);
  assign n35268 = (n30165 & n30547) | (n30165 & n35266) | (n30547 & n35266);
  assign n35269 = (n34922 & n35267) | (n34922 & n35268) | (n35267 & n35268);
  assign n30549 = n20975 & ~n35269;
  assign n30550 = n30542 & n30549;
  assign n30551 = ~n20975 & n35269;
  assign n30552 = (n20975 & n30542) | (n20975 & ~n30551) | (n30542 & ~n30551);
  assign n20978 = ~n30550 & n30552;
  assign n30559 = n20490 | n20717;
  assign n35270 = (n20717 & n20719) | (n20717 & n30559) | (n20719 & n30559);
  assign n30556 = n20978 | n35270;
  assign n30554 = n20717 | n20719;
  assign n30557 = n20978 | n30554;
  assign n35271 = (n30331 & n30556) | (n30331 & n30557) | (n30556 & n30557);
  assign n35272 = (n30332 & n30556) | (n30332 & n30557) | (n30556 & n30557);
  assign n35273 = (n30215 & n35271) | (n30215 & n35272) | (n35271 & n35272);
  assign n20982 = n20968 & ~n20975;
  assign n20983 = ~n20968 & n20975;
  assign n20984 = n20982 | n20983;
  assign n30561 = n20710 | n20984;
  assign n30562 = n35187 | n30561;
  assign n30563 = n20710 & n20984;
  assign n30564 = (n20984 & n35187) | (n20984 & n30563) | (n35187 & n30563);
  assign n30565 = n30562 & ~n30564;
  assign n30566 = n20718 & n30565;
  assign n30567 = n30559 & n30566;
  assign n35274 = (n30331 & n30566) | (n30331 & n30567) | (n30566 & n30567);
  assign n35275 = (n30332 & n30566) | (n30332 & n30567) | (n30566 & n30567);
  assign n35276 = (n30215 & n35274) | (n30215 & n35275) | (n35274 & n35275);
  assign n20990 = n35273 & ~n35276;
  assign n20991 = x131 & x148;
  assign n20992 = n20990 & n20991;
  assign n20993 = n20990 | n20991;
  assign n20994 = ~n20992 & n20993;
  assign n20995 = x130 & x149;
  assign n20996 = n20994 & n20995;
  assign n20997 = n20994 | n20995;
  assign n20998 = ~n20996 & n20997;
  assign n30569 = ~n20724 & n20998;
  assign n30570 = ~n30531 & n30569;
  assign n30571 = n20724 & ~n20998;
  assign n30572 = (~n20998 & n30531) | (~n20998 & n30571) | (n30531 & n30571);
  assign n21001 = n30570 | n30572;
  assign n21002 = x129 & x150;
  assign n21003 = n21001 & n21002;
  assign n21004 = n21001 | n21002;
  assign n21005 = ~n21003 & n21004;
  assign n30573 = n20952 | n21005;
  assign n30574 = n35247 | n30573;
  assign n30575 = n20952 & n21005;
  assign n30576 = (n21005 & n35247) | (n21005 & n30575) | (n35247 & n30575);
  assign n21008 = n30574 & ~n30576;
  assign n21009 = x128 & x151;
  assign n21010 = n21008 | n21009;
  assign n21011 = n21008 & n21009;
  assign n21012 = n21010 & ~n21011;
  assign n30577 = ~n20944 & n21012;
  assign n30578 = ~n30515 & n30577;
  assign n30579 = n20944 & ~n21012;
  assign n30580 = (~n21012 & n30515) | (~n21012 & n30579) | (n30515 & n30579);
  assign n21015 = n30578 | n30580;
  assign n21016 = x127 & x152;
  assign n21017 = n21015 & n21016;
  assign n21018 = n21015 | n21016;
  assign n21019 = ~n21017 & n21018;
  assign n21020 = ~n30518 & n21019;
  assign n21021 = n30518 & ~n21019;
  assign n21022 = n21020 | n21021;
  assign n21023 = x126 & x153;
  assign n21024 = n21022 | n21023;
  assign n21025 = n21022 & n21023;
  assign n21026 = n21024 & ~n21025;
  assign n21027 = ~n30508 & n21026;
  assign n21028 = n30508 & ~n21026;
  assign n21029 = n21027 | n21028;
  assign n21030 = x125 & x154;
  assign n21031 = n21029 & n21030;
  assign n21032 = n21029 | n21030;
  assign n21033 = ~n21031 & n21032;
  assign n21034 = n30500 | n21033;
  assign n21035 = n30500 & n21033;
  assign n21036 = n21034 & ~n21035;
  assign n21037 = x124 & x155;
  assign n21038 = n21036 | n21037;
  assign n21039 = n21036 & n21037;
  assign n21040 = n21038 & ~n21039;
  assign n21041 = n30491 | n21040;
  assign n21042 = n30491 & n21040;
  assign n21043 = n21041 & ~n21042;
  assign n30581 = n20911 | n21043;
  assign n30582 = n30455 | n30581;
  assign n30583 = n20911 & n21043;
  assign n30584 = (n21043 & n30455) | (n21043 & n30583) | (n30455 & n30583);
  assign n21046 = n30582 & ~n30584;
  assign n21047 = x123 & x156;
  assign n21048 = x122 & x157;
  assign n21049 = n21047 & n21048;
  assign n21050 = n21047 | n21048;
  assign n21051 = ~n21049 & n21050;
  assign n21052 = n21046 & n21051;
  assign n21053 = n21046 | n21051;
  assign n21054 = ~n21052 & n21053;
  assign n21055 = n30487 | n21054;
  assign n21056 = n30487 & n21054;
  assign n21057 = n21055 & ~n21056;
  assign n21058 = x121 & x158;
  assign n21059 = n21057 | n21058;
  assign n21060 = n21057 & n21058;
  assign n21061 = n21059 & ~n21060;
  assign n30585 = n20803 & n20811;
  assign n30586 = (n20803 & n30457) | (n20803 & n30585) | (n30457 & n30585);
  assign n21063 = n30381 | n20905;
  assign n30587 = n20794 & ~n20905;
  assign n30588 = (n20794 & ~n30381) | (n20794 & n30587) | (~n30381 & n30587);
  assign n21065 = n21063 & n30588;
  assign n21066 = n30586 | n21065;
  assign n21067 = ~n21061 & n21066;
  assign n21068 = n21061 & ~n21066;
  assign n21069 = n21067 | n21068;
  assign n21070 = x120 & x159;
  assign n21071 = n21069 & n21070;
  assign n21072 = n21069 | n21070;
  assign n21073 = ~n21071 & n21072;
  assign n30484 = n20815 & n20822;
  assign n30485 = (n20815 & n30379) | (n20815 & n30484) | (n30379 & n30484);
  assign n30589 = n20803 | n20811;
  assign n30590 = n30457 | n30589;
  assign n21075 = n20804 & ~n30586;
  assign n21076 = n30590 & n21075;
  assign n21077 = n30485 | n21076;
  assign n21078 = ~n21073 & n21077;
  assign n21079 = n21073 & ~n21077;
  assign n21080 = n21078 | n21079;
  assign n30482 = n20815 | n20822;
  assign n30483 = n30379 | n30482;
  assign n20900 = n20816 & ~n30485;
  assign n20901 = n30483 & n20900;
  assign n30591 = n20901 & n21080;
  assign n30592 = (n21080 & n30463) | (n21080 & n30591) | (n30463 & n30591);
  assign n30593 = n20901 | n21080;
  assign n30594 = n30463 | n30593;
  assign n21083 = ~n30592 & n30594;
  assign n21084 = ~n20897 & n21083;
  assign n21085 = n20897 & ~n21083;
  assign n21086 = n21084 | n21085;
  assign n20895 = n20646 & n20829;
  assign n30595 = n20895 & n21086;
  assign n30596 = (n21086 & n30467) | (n21086 & n30595) | (n30467 & n30595);
  assign n30597 = n20895 | n21086;
  assign n30598 = n30467 | n30597;
  assign n21089 = ~n30596 & n30598;
  assign n21090 = n20894 & n21089;
  assign n21091 = n20894 | n21089;
  assign n21092 = ~n21090 & n21091;
  assign n21093 = n30481 & n21092;
  assign n21094 = n30481 | n21092;
  assign n21095 = ~n21093 & n21094;
  assign n21096 = n20892 | n21095;
  assign n21097 = n20892 & n21095;
  assign n21098 = n21096 & ~n21097;
  assign n21099 = ~n20891 & n21098;
  assign n21100 = n20891 & ~n21098;
  assign n21101 = n21099 | n21100;
  assign n30599 = n20851 & n20852;
  assign n30600 = (n20851 & n20860) | (n20851 & n30599) | (n20860 & n30599);
  assign n21104 = n21101 & ~n30600;
  assign n21105 = ~n21101 & n30600;
  assign n21106 = n21104 | n21105;
  assign n21107 = x115 & x164;
  assign n21108 = n21106 | n21107;
  assign n21109 = n21106 & n21107;
  assign n21110 = n21108 & ~n21109;
  assign n35277 = n20864 & n30472;
  assign n35278 = n20630 & n20864;
  assign n35279 = (n20407 & n35277) | (n20407 & n35278) | (n35277 & n35278);
  assign n30604 = n20869 & n35279;
  assign n35280 = n20864 | n30472;
  assign n35281 = n20630 | n20864;
  assign n35282 = (n20407 & n35280) | (n20407 & n35281) | (n35280 & n35281);
  assign n30602 = (n20864 & n20869) | (n20864 & n35282) | (n20869 & n35282);
  assign n30605 = n30602 | n30604;
  assign n30606 = (n20863 & n30604) | (n20863 & n30605) | (n30604 & n30605);
  assign n21115 = n21110 & ~n30606;
  assign n21116 = ~n21110 & n30606;
  assign n21117 = n21115 | n21116;
  assign n21118 = x114 & x165;
  assign n21119 = n21117 & n21118;
  assign n21120 = n21117 | n21118;
  assign n21121 = ~n21119 & n21120;
  assign n30473 = (n20407 & n20630) | (n20407 & n30472) | (n20630 & n30472);
  assign n20871 = n20869 & n30473;
  assign n21123 = ~n20867 & n20871;
  assign n30607 = n20637 & n20872;
  assign n30608 = n20636 & n30607;
  assign n21125 = n21123 | n30608;
  assign n30609 = n20637 | n20872;
  assign n30610 = (n20636 & n20872) | (n20636 & n30609) | (n20872 & n30609);
  assign n21122 = n20867 & ~n20871;
  assign n30611 = n21122 & n30610;
  assign n30612 = (n21125 & n30610) | (n21125 & n30611) | (n30610 & n30611);
  assign n21129 = n21121 & ~n30612;
  assign n21130 = ~n21121 & n30612;
  assign n21131 = n21129 | n21130;
  assign n21132 = x113 & x166;
  assign n21133 = n21131 | n21132;
  assign n21134 = n21131 & n21132;
  assign n21135 = n21133 & ~n21134;
  assign n21136 = ~n20883 & n21135;
  assign n21137 = n20883 & ~n21135;
  assign n21138 = n21136 | n21137;
  assign n21139 = x112 & x167;
  assign n21140 = n21138 & n21139;
  assign n21141 = n21138 | n21139;
  assign n21142 = ~n21140 & n21141;
  assign n30613 = n21096 & n21097;
  assign n30614 = (n21096 & n30479) | (n21096 & n30613) | (n30479 & n30613);
  assign n21145 = x117 & x163;
  assign n21146 = n30614 & n21145;
  assign n21147 = n30614 | n21145;
  assign n21148 = ~n21146 & n21147;
  assign n30615 = n21069 & n21076;
  assign n30616 = (n21069 & n30485) | (n21069 & n30615) | (n30485 & n30615);
  assign n30617 = n21057 & n21065;
  assign n30618 = (n21057 & n30586) | (n21057 & n30617) | (n30586 & n30617);
  assign n30619 = n21057 | n21065;
  assign n30620 = n30586 | n30619;
  assign n21152 = n21058 & n30620;
  assign n21153 = ~n30618 & n21152;
  assign n21154 = n30616 | n21153;
  assign n21156 = n21046 | n21047;
  assign n21155 = n21046 & n21047;
  assign n30623 = n21155 & n21156;
  assign n30624 = (n21156 & n30487) | (n21156 & n30623) | (n30487 & n30623);
  assign n30625 = n21036 & n30490;
  assign n30626 = n20916 & n21036;
  assign n30627 = (n30451 & n30625) | (n30451 & n30626) | (n30625 & n30626);
  assign n30628 = n21036 | n30490;
  assign n30629 = n20916 | n21036;
  assign n30630 = (n30451 & n30628) | (n30451 & n30629) | (n30628 & n30629);
  assign n21167 = n21037 & n30630;
  assign n21168 = ~n30627 & n21167;
  assign n21169 = n30584 | n21168;
  assign n21170 = n20926 | n21029;
  assign n30631 = n20765 | n21170;
  assign n30632 = (n21170 & n30449) | (n21170 & n30631) | (n30449 & n30631);
  assign n21173 = n20759 | n20925;
  assign n21174 = n21029 & n21173;
  assign n30633 = n20926 & n21174;
  assign n30634 = (n21174 & n30449) | (n21174 & n30633) | (n30449 & n30633);
  assign n21176 = n30632 & ~n30634;
  assign n21177 = n21030 & n21176;
  assign n21178 = n30627 | n21177;
  assign n35283 = n21022 & n30507;
  assign n35284 = n20931 & n21022;
  assign n35285 = (n30493 & n35283) | (n30493 & n35284) | (n35283 & n35284);
  assign n35286 = (n21023 & n21025) | (n21023 & n30507) | (n21025 & n30507);
  assign n37362 = n20931 & n21023;
  assign n37363 = (n21022 & n21023) | (n21022 & n37362) | (n21023 & n37362);
  assign n35288 = (n30493 & n35286) | (n30493 & n37363) | (n35286 & n37363);
  assign n21182 = ~n35285 & n35288;
  assign n21185 = n20741 | n20938;
  assign n21186 = n21015 & n21185;
  assign n35289 = n20741 | n20754;
  assign n35290 = (n20754 & n20938) | (n20754 & n35289) | (n20938 & n35289);
  assign n30638 = n21186 & n35290;
  assign n30639 = (n21186 & n30384) | (n21186 & n30638) | (n30384 & n30638);
  assign n30645 = n20944 & n21008;
  assign n35291 = (n21008 & n30514) | (n21008 & n30645) | (n30514 & n30645);
  assign n35292 = (n20936 & n21008) | (n20936 & n30645) | (n21008 & n30645);
  assign n35293 = (n30284 & n35291) | (n30284 & n35292) | (n35291 & n35292);
  assign n30647 = n20944 | n21008;
  assign n30649 = n21009 & n30647;
  assign n35294 = (n21009 & n30514) | (n21009 & n30649) | (n30514 & n30649);
  assign n35295 = (n20936 & n21009) | (n20936 & n30649) | (n21009 & n30649);
  assign n35296 = (n30284 & n35294) | (n30284 & n35295) | (n35294 & n35295);
  assign n21196 = ~n35293 & n35296;
  assign n21198 = n20952 | n21001;
  assign n21199 = n35247 | n21198;
  assign n30396 = (n20676 & n30154) | (n20676 & n30395) | (n30154 & n30395);
  assign n21202 = n20727 | n20951;
  assign n21203 = n21001 & n21202;
  assign n21200 = n20688 | n20952;
  assign n30651 = n20680 | n21200;
  assign n35297 = n21203 & n30651;
  assign n35298 = n21200 & n21203;
  assign n35299 = (n30396 & n35297) | (n30396 & n35298) | (n35297 & n35298);
  assign n21205 = n21199 & ~n35299;
  assign n21206 = n21002 & n21205;
  assign n30653 = n21206 | n30645;
  assign n30654 = n21008 | n21206;
  assign n35300 = (n30514 & n30653) | (n30514 & n30654) | (n30653 & n30654);
  assign n35301 = (n20936 & n30653) | (n20936 & n30654) | (n30653 & n30654);
  assign n35302 = (n30284 & n35300) | (n30284 & n35301) | (n35300 & n35301);
  assign n21208 = x129 & x151;
  assign n30652 = (n21200 & n30396) | (n21200 & n30651) | (n30396 & n30651);
  assign n21215 = x132 & x148;
  assign n30333 = (n30215 & n30331) | (n30215 & n30332) | (n30331 & n30332);
  assign n21217 = x133 & x147;
  assign n21224 = x136 & x144;
  assign n21225 = x135 & x145;
  assign n21226 = n21224 | n21225;
  assign n21227 = n21224 & n21225;
  assign n21228 = n21226 & ~n21227;
  assign n21229 = n20960 & n21228;
  assign n37364 = n20959 & n20960;
  assign n37365 = n21228 & n37364;
  assign n37366 = (n21229 & n37361) | (n21229 & n37365) | (n37361 & n37365);
  assign n37367 = (n20700 & n21229) | (n20700 & n37365) | (n21229 & n37365);
  assign n37368 = (n30428 & n37366) | (n30428 & n37367) | (n37366 & n37367);
  assign n35305 = (n21229 & n35258) | (n21229 & n37365) | (n35258 & n37365);
  assign n35306 = (n37347 & n37368) | (n37347 & n35305) | (n37368 & n35305);
  assign n35307 = (n35096 & n37368) | (n35096 & n35305) | (n37368 & n35305);
  assign n35308 = (n29868 & n35306) | (n29868 & n35307) | (n35306 & n35307);
  assign n21231 = n20959 | n21228;
  assign n35309 = n20961 | n21231;
  assign n35310 = (n21231 & n35256) | (n21231 & n35309) | (n35256 & n35309);
  assign n35311 = (n21231 & n35258) | (n21231 & n35309) | (n35258 & n35309);
  assign n35312 = (n37347 & n35310) | (n37347 & n35311) | (n35310 & n35311);
  assign n35313 = (n35096 & n35310) | (n35096 & n35311) | (n35310 & n35311);
  assign n35314 = (n29868 & n35312) | (n29868 & n35313) | (n35312 & n35313);
  assign n21233 = ~n35308 & n35314;
  assign n21234 = x134 & x146;
  assign n21235 = n21233 & n21234;
  assign n21236 = n21233 | n21234;
  assign n21237 = ~n21235 & n21236;
  assign n37369 = n20961 & n37361;
  assign n37370 = n20700 & n20961;
  assign n37371 = (n30428 & n37369) | (n30428 & n37370) | (n37369 & n37370);
  assign n30671 = n20961 & n35258;
  assign n35315 = (n37347 & n37371) | (n37347 & n30671) | (n37371 & n30671);
  assign n35316 = (n37371 & n30671) | (n37371 & n35096) | (n30671 & n35096);
  assign n35317 = (n29868 & n35315) | (n29868 & n35316) | (n35315 & n35316);
  assign n37372 = (n20962 & n20963) | (n20962 & n37361) | (n20963 & n37361);
  assign n37741 = n20700 & n20962;
  assign n37742 = (n20961 & n20962) | (n20961 & n37741) | (n20962 & n37741);
  assign n37374 = (n30428 & n37372) | (n30428 & n37742) | (n37372 & n37742);
  assign n35319 = (n20962 & n20963) | (n20962 & n35258) | (n20963 & n35258);
  assign n35320 = (n37347 & n37374) | (n37347 & n35319) | (n37374 & n35319);
  assign n35321 = (n35096 & n37374) | (n35096 & n35319) | (n37374 & n35319);
  assign n35322 = (n29868 & n35320) | (n29868 & n35321) | (n35320 & n35321);
  assign n21221 = ~n35317 & n35322;
  assign n30688 = n21221 & n21237;
  assign n30689 = (n21237 & n35269) | (n21237 & n30688) | (n35269 & n30688);
  assign n30690 = n21221 | n21237;
  assign n30691 = n35269 | n30690;
  assign n21240 = ~n30689 & n30691;
  assign n21241 = n21217 & n21240;
  assign n21242 = n21217 | n21240;
  assign n21243 = ~n21241 & n21242;
  assign n30667 = n30550 | n30567;
  assign n30692 = n21243 & n30667;
  assign n30668 = n30550 | n30566;
  assign n30693 = n21243 & n30668;
  assign n30694 = (n30333 & n30692) | (n30333 & n30693) | (n30692 & n30693);
  assign n30695 = n21243 | n30667;
  assign n30696 = n21243 | n30668;
  assign n30697 = (n30333 & n30695) | (n30333 & n30696) | (n30695 & n30696);
  assign n21246 = ~n30694 & n30697;
  assign n21247 = n21215 & n21246;
  assign n21248 = n21215 | n21246;
  assign n21249 = ~n21247 & n21248;
  assign n21250 = x131 & x149;
  assign n21251 = n21249 & n21250;
  assign n21252 = n21249 | n21250;
  assign n21253 = ~n21251 & n21252;
  assign n21476 = n20724 | n20992;
  assign n35323 = (n20992 & n20994) | (n20992 & n21476) | (n20994 & n21476);
  assign n30698 = n21253 | n35323;
  assign n30665 = n20992 | n20994;
  assign n30699 = n21253 | n30665;
  assign n30700 = (n30531 & n30698) | (n30531 & n30699) | (n30698 & n30699);
  assign n30701 = n21253 & n35323;
  assign n30702 = n21253 & n30665;
  assign n30703 = (n30531 & n30701) | (n30531 & n30702) | (n30701 & n30702);
  assign n21256 = n30700 & ~n30703;
  assign n21257 = x130 & x150;
  assign n21258 = n21256 | n21257;
  assign n21259 = n21256 & n21257;
  assign n21260 = n21258 & ~n21259;
  assign n30656 = n20724 & n20994;
  assign n35324 = (n20994 & n30656) | (n20994 & n35254) | (n30656 & n35254);
  assign n35325 = (n20949 & n20994) | (n20949 & n30656) | (n20994 & n30656);
  assign n35326 = (n35091 & n35324) | (n35091 & n35325) | (n35324 & n35325);
  assign n37375 = n20723 & n20995;
  assign n37376 = n20722 & n37375;
  assign n35328 = (n20994 & n20995) | (n20994 & n37376) | (n20995 & n37376);
  assign n35329 = (n20995 & n35254) | (n20995 & n35328) | (n35254 & n35328);
  assign n35330 = (n20949 & n20995) | (n20949 & n35328) | (n20995 & n35328);
  assign n35331 = (n35091 & n35329) | (n35091 & n35330) | (n35329 & n35330);
  assign n21212 = ~n35326 & n35331;
  assign n30662 = n21203 | n21212;
  assign n30704 = n21260 & n30662;
  assign n30705 = n21212 & n21260;
  assign n30706 = (n30652 & n30704) | (n30652 & n30705) | (n30704 & n30705);
  assign n30707 = n21260 | n30662;
  assign n30708 = n21212 | n21260;
  assign n30709 = (n30652 & n30707) | (n30652 & n30708) | (n30707 & n30708);
  assign n21263 = ~n30706 & n30709;
  assign n21264 = n21208 & n21263;
  assign n21265 = n21208 | n21263;
  assign n21266 = ~n21264 & n21265;
  assign n21267 = x128 & x152;
  assign n21268 = n21266 & ~n21267;
  assign n21269 = ~n21266 & n21267;
  assign n21270 = n21268 | n21269;
  assign n21271 = n35302 | n21270;
  assign n21272 = n35302 & n21270;
  assign n21273 = n21271 & ~n21272;
  assign n30710 = ~n21196 & n21273;
  assign n30711 = ~n30639 & n30710;
  assign n30712 = n21196 & ~n21273;
  assign n30713 = (~n21273 & n30639) | (~n21273 & n30712) | (n30639 & n30712);
  assign n21276 = n30711 | n30713;
  assign n21277 = x127 & x153;
  assign n21278 = n21276 & n21277;
  assign n21279 = n21276 | n21277;
  assign n21280 = ~n21278 & n21279;
  assign n21188 = n20939 | n21015;
  assign n30640 = n21188 | n30501;
  assign n30641 = n20747 | n21188;
  assign n30642 = (n30384 & n30640) | (n30384 & n30641) | (n30640 & n30641);
  assign n21190 = ~n30639 & n30642;
  assign n21191 = n21016 & n21190;
  assign n30643 = n21022 | n21191;
  assign n30714 = n21280 & ~n30643;
  assign n30715 = ~n21191 & n21280;
  assign n30716 = (~n30508 & n30714) | (~n30508 & n30715) | (n30714 & n30715);
  assign n30717 = ~n21280 & n30643;
  assign n30718 = n21191 & ~n21280;
  assign n30719 = (n30508 & n30717) | (n30508 & n30718) | (n30717 & n30718);
  assign n21283 = n30716 | n30719;
  assign n21284 = x126 & x154;
  assign n21285 = n21283 | n21284;
  assign n21286 = n21283 & n21284;
  assign n21287 = n21285 & ~n21286;
  assign n30720 = ~n21182 & n21287;
  assign n30721 = ~n30634 & n30720;
  assign n30722 = n21182 & ~n21287;
  assign n30723 = (~n21287 & n30634) | (~n21287 & n30722) | (n30634 & n30722);
  assign n21290 = n30721 | n30723;
  assign n21291 = x125 & x155;
  assign n21292 = n21290 & n21291;
  assign n21293 = n21290 | n21291;
  assign n21294 = ~n21292 & n21293;
  assign n21295 = x124 & x156;
  assign n21296 = n21294 & ~n21295;
  assign n21297 = ~n21294 & n21295;
  assign n21298 = n21296 | n21297;
  assign n21299 = n21178 | n21298;
  assign n21300 = n21178 & n21298;
  assign n21301 = n21299 & ~n21300;
  assign n21302 = ~n21169 & n21301;
  assign n21303 = n21169 & ~n21301;
  assign n21304 = n21302 | n21303;
  assign n21305 = x123 & x157;
  assign n21306 = n21304 & n21305;
  assign n21307 = n21304 | n21305;
  assign n21308 = ~n21306 & n21307;
  assign n21309 = n30624 & n21308;
  assign n21310 = n30624 | n21308;
  assign n21311 = ~n21309 & n21310;
  assign n21157 = ~n21155 & n21156;
  assign n21158 = n30487 | n21157;
  assign n30621 = n21048 & ~n21157;
  assign n30622 = (n21048 & ~n30487) | (n21048 & n30621) | (~n30487 & n30621);
  assign n21161 = n21158 & n30622;
  assign n30724 = n21161 & n21311;
  assign n30725 = (n21311 & n30618) | (n21311 & n30724) | (n30618 & n30724);
  assign n30726 = n21161 | n21311;
  assign n30727 = n30618 | n30726;
  assign n21314 = ~n30725 & n30727;
  assign n21315 = x122 & x158;
  assign n21316 = n21314 & n21315;
  assign n21317 = n21314 | n21315;
  assign n21318 = ~n21316 & n21317;
  assign n21319 = n21154 | n21318;
  assign n21320 = n21154 & n21318;
  assign n21321 = n21319 & ~n21320;
  assign n21322 = x121 & x159;
  assign n21323 = n21321 | n21322;
  assign n21324 = n21321 & n21322;
  assign n21325 = n21323 & ~n21324;
  assign n30728 = n21069 | n21076;
  assign n30729 = n30485 | n30728;
  assign n21327 = n21070 & ~n30616;
  assign n21328 = n30729 & n21327;
  assign n21329 = n30592 | n21328;
  assign n21330 = n21325 & ~n21329;
  assign n21331 = ~n21325 & n21329;
  assign n21332 = n21330 | n21331;
  assign n21333 = x120 & x160;
  assign n21334 = n21332 | n21333;
  assign n21335 = n21332 & n21333;
  assign n21336 = n21334 & ~n21335;
  assign n21339 = x119 & x161;
  assign n35332 = n20897 & ~n21339;
  assign n35333 = n21083 & n35332;
  assign n30731 = (~n21339 & n30596) | (~n21339 & n35333) | (n30596 & n35333);
  assign n35334 = ~n20897 & n21339;
  assign n35335 = (~n21083 & n21339) | (~n21083 & n35334) | (n21339 & n35334);
  assign n30733 = ~n30596 & n35335;
  assign n21342 = n30731 | n30733;
  assign n21343 = ~n21336 & n21342;
  assign n21344 = n21336 & ~n21342;
  assign n21345 = n21343 | n21344;
  assign n30734 = n21090 | n21092;
  assign n30735 = (n21090 & n30481) | (n21090 & n30734) | (n30481 & n30734);
  assign n21347 = n21345 & ~n30735;
  assign n21348 = ~n21345 & n30735;
  assign n21349 = n21347 | n21348;
  assign n21350 = x118 & x162;
  assign n21351 = n21349 | n21350;
  assign n21352 = n21349 & n21350;
  assign n21353 = n21351 & ~n21352;
  assign n21354 = ~n21148 & n21353;
  assign n21355 = n21148 & ~n21353;
  assign n21356 = n21354 | n21355;
  assign n21357 = ~n30479 & n21098;
  assign n21358 = n30479 & ~n21098;
  assign n21359 = n21357 | n21358;
  assign n21362 = n20888 | n21359;
  assign n21360 = n20888 & n21359;
  assign n30736 = n21360 & n21362;
  assign n30737 = (n21362 & n30600) | (n21362 & n30736) | (n30600 & n30736);
  assign n21364 = n21356 & ~n30737;
  assign n21365 = ~n21356 & n30737;
  assign n21366 = n21364 | n21365;
  assign n21367 = x116 & x164;
  assign n21368 = n21366 | n21367;
  assign n21369 = n21366 & n21367;
  assign n21370 = n21368 & ~n21369;
  assign n21371 = n21109 | n30606;
  assign n21372 = n21108 & n21371;
  assign n21373 = n21370 & ~n21372;
  assign n21374 = ~n21370 & n21372;
  assign n21375 = n21373 | n21374;
  assign n21376 = x115 & x165;
  assign n21377 = n21375 | n21376;
  assign n21378 = n21375 & n21376;
  assign n21379 = n21377 & ~n21378;
  assign n21380 = n21119 | n30612;
  assign n21381 = n21120 & n21380;
  assign n21382 = n21379 & ~n21381;
  assign n21383 = ~n21379 & n21381;
  assign n21384 = n21382 | n21383;
  assign n21385 = x114 & x166;
  assign n21386 = n21384 | n21385;
  assign n21387 = n21384 & n21385;
  assign n21388 = n21386 & ~n21387;
  assign n35336 = n20882 | n21132;
  assign n35337 = (n20881 & n21132) | (n20881 & n35336) | (n21132 & n35336);
  assign n30739 = (n20883 & n21131) | (n20883 & n35337) | (n21131 & n35337);
  assign n21390 = n21133 & n30739;
  assign n21391 = n21388 & ~n21390;
  assign n21392 = ~n21388 & n21390;
  assign n21393 = n21391 | n21392;
  assign n21394 = x113 & x167;
  assign n21395 = n21393 | n21394;
  assign n21396 = n21393 & n21394;
  assign n21397 = n21395 & ~n21396;
  assign n21398 = ~n21140 & n21397;
  assign n21399 = n21140 & ~n21397;
  assign n21400 = n21398 | n21399;
  assign n21401 = x112 & x168;
  assign n21402 = n21400 & n21401;
  assign n21403 = n21400 | n21401;
  assign n21404 = ~n21402 & n21403;
  assign n21405 = x115 & x166;
  assign n30740 = n21377 & n21378;
  assign n30741 = (n21377 & n21381) | (n21377 & n30740) | (n21381 & n30740);
  assign n21408 = x116 & x165;
  assign n30742 = n21368 & n21369;
  assign n30743 = (n21368 & n21372) | (n21368 & n30742) | (n21372 & n30742);
  assign n21337 = n20897 & n21083;
  assign n21338 = n30596 | n21337;
  assign n21411 = n21336 & ~n21338;
  assign n21412 = ~n21336 & n21338;
  assign n21413 = n21411 | n21412;
  assign n21416 = n21339 | n21413;
  assign n21414 = n21339 & n21413;
  assign n30744 = n21414 & n21416;
  assign n30745 = (n21416 & n30735) | (n21416 & n30744) | (n30735 & n30744);
  assign n37377 = n20897 | n21333;
  assign n37378 = (n21083 & n21333) | (n21083 & n37377) | (n21333 & n37377);
  assign n35339 = (n21332 & n21337) | (n21332 & n37378) | (n21337 & n37378);
  assign n35340 = n21334 & n35339;
  assign n35341 = (n21334 & n30596) | (n21334 & n35340) | (n30596 & n35340);
  assign n21420 = x121 & x160;
  assign n21421 = x120 & x161;
  assign n21422 = n21420 & n21421;
  assign n21423 = n21420 | n21421;
  assign n21424 = ~n21422 & n21423;
  assign n30748 = n21323 & n21324;
  assign n30749 = (n21323 & n21329) | (n21323 & n30748) | (n21329 & n30748);
  assign n30863 = n21304 | n30623;
  assign n30864 = n21156 | n21304;
  assign n30865 = (n30487 & n30863) | (n30487 & n30864) | (n30863 & n30864);
  assign n21163 = n30487 | n21155;
  assign n37379 = ~n21047 & n21305;
  assign n37380 = ~n21046 & n37379;
  assign n35343 = (~n21304 & n21305) | (~n21304 & n37380) | (n21305 & n37380);
  assign n30867 = (~n21163 & n21305) | (~n21163 & n35343) | (n21305 & n35343);
  assign n21607 = n30865 & n30867;
  assign n21608 = n30725 | n21607;
  assign n21427 = n21178 | n21294;
  assign n21428 = n21178 & n21294;
  assign n21429 = n21427 & ~n21428;
  assign n30750 = n21168 & n21429;
  assign n30751 = (n21429 & n30584) | (n21429 & n30750) | (n30584 & n30750);
  assign n21431 = n21177 | n21290;
  assign n21432 = n30627 | n21431;
  assign n35344 = n20916 | n21030;
  assign n35345 = (n20916 & n21176) | (n20916 & n35344) | (n21176 & n35344);
  assign n21435 = n21030 | n21176;
  assign n21436 = n21290 & n21435;
  assign n30752 = n35345 & n21436;
  assign n35346 = n21291 & ~n21436;
  assign n35347 = n21291 & ~n35233;
  assign n35348 = (~n30752 & n35346) | (~n30752 & n35347) | (n35346 & n35347);
  assign n21439 = n21432 & n35348;
  assign n21440 = n30751 | n21439;
  assign n21441 = x125 & x156;
  assign n21447 = n21191 | n21276;
  assign n30760 = n21022 | n21447;
  assign n30761 = (n21447 & n30508) | (n21447 & n30760) | (n30508 & n30760);
  assign n21449 = n20931 | n21191;
  assign n30762 = n20922 | n21449;
  assign n30763 = (n21449 & n30493) | (n21449 & n30762) | (n30493 & n30762);
  assign n21451 = n21016 | n21190;
  assign n21452 = n21276 & n21451;
  assign n21453 = n30763 & n21452;
  assign n21454 = n30761 & ~n21453;
  assign n21455 = n21277 & n21454;
  assign n30754 = n21182 & n21283;
  assign n30764 = n21455 | n30754;
  assign n30765 = n21283 | n21455;
  assign n30766 = (n30634 & n30764) | (n30634 & n30765) | (n30764 & n30765);
  assign n21461 = n21206 | n21263;
  assign n30775 = n21461 | n30645;
  assign n30776 = n21008 | n21461;
  assign n30777 = (n30515 & n30775) | (n30515 & n30776) | (n30775 & n30776);
  assign n21463 = n20944 | n21206;
  assign n21465 = n21002 | n21205;
  assign n21466 = n21263 & n21465;
  assign n30778 = n21463 & n21466;
  assign n35349 = n21208 & ~n30778;
  assign n35350 = n21208 & ~n21466;
  assign n35351 = (~n30515 & n35349) | (~n30515 & n35350) | (n35349 & n35350);
  assign n21469 = n30777 & n35351;
  assign n30767 = n21266 | n30654;
  assign n30768 = n21266 | n30653;
  assign n30769 = (n30515 & n30767) | (n30515 & n30768) | (n30767 & n30768);
  assign n30770 = n21266 & n30654;
  assign n30771 = n21266 & n30653;
  assign n30772 = (n30515 & n30770) | (n30515 & n30771) | (n30770 & n30771);
  assign n21459 = n30769 & ~n30772;
  assign n30773 = n21196 & n21459;
  assign n30780 = n21469 | n30773;
  assign n30781 = n21459 | n21469;
  assign n30782 = (n30639 & n30780) | (n30639 & n30781) | (n30780 & n30781);
  assign n30779 = (n21466 & n30515) | (n21466 & n30778) | (n30515 & n30778);
  assign n30784 = n21212 & n21256;
  assign n35352 = (n21203 & n21256) | (n21203 & n30784) | (n21256 & n30784);
  assign n35353 = (n30651 & n30784) | (n30651 & n35352) | (n30784 & n35352);
  assign n35354 = (n21200 & n30784) | (n21200 & n35352) | (n30784 & n35352);
  assign n35355 = (n30396 & n35353) | (n30396 & n35354) | (n35353 & n35354);
  assign n30787 = n21212 | n21256;
  assign n35356 = n21203 | n30787;
  assign n35357 = (n30651 & n30787) | (n30651 & n35356) | (n30787 & n35356);
  assign n35358 = (n21200 & n30787) | (n21200 & n35356) | (n30787 & n35356);
  assign n35359 = (n30396 & n35357) | (n30396 & n35358) | (n35357 & n35358);
  assign n21473 = n21257 & n35359;
  assign n21474 = ~n35355 & n21473;
  assign n21478 = n20993 & n21249;
  assign n35360 = n20993 & n21476;
  assign n35361 = n21249 & n35360;
  assign n35362 = (n21478 & n35254) | (n21478 & n35361) | (n35254 & n35361);
  assign n35363 = (n20949 & n21478) | (n20949 & n35361) | (n21478 & n35361);
  assign n35364 = (n35091 & n35362) | (n35091 & n35363) | (n35362 & n35363);
  assign n30791 = n21249 | n35323;
  assign n30792 = n21249 | n30665;
  assign n35365 = (n30791 & n30792) | (n30791 & n35254) | (n30792 & n35254);
  assign n35366 = (n20949 & n30791) | (n20949 & n30792) | (n30791 & n30792);
  assign n35367 = (n35091 & n35365) | (n35091 & n35366) | (n35365 & n35366);
  assign n21481 = ~n35364 & n35367;
  assign n21482 = n21250 & n21481;
  assign n21490 = x137 & x144;
  assign n21491 = x136 & x145;
  assign n21492 = n21490 & n21491;
  assign n21493 = n21490 | n21491;
  assign n21494 = ~n21492 & n21493;
  assign n21495 = x135 & x146;
  assign n21496 = n21494 & n21495;
  assign n21497 = n21494 | n21495;
  assign n21498 = ~n21496 & n21497;
  assign n37381 = n20960 | n21227;
  assign n37382 = (n21227 & n21228) | (n21227 & n37381) | (n21228 & n37381);
  assign n21485 = n20698 | n21225;
  assign n21486 = n20697 & n21485;
  assign n35375 = n20704 | n21486;
  assign n35376 = (n20706 & n21486) | (n20706 & n35375) | (n21486 & n35375);
  assign n35377 = (n21227 & n37382) | (n21227 & n35376) | (n37382 & n35376);
  assign n30807 = n21498 & ~n35377;
  assign n35368 = n20706 | n21486;
  assign n35369 = (n21486 & n30428) | (n21486 & n35368) | (n30428 & n35368);
  assign n35372 = n21498 & ~n37382;
  assign n35373 = ~n21227 & n21498;
  assign n35374 = (~n35369 & n35372) | (~n35369 & n35373) | (n35372 & n35373);
  assign n35378 = (~n37347 & n30807) | (~n37347 & n35374) | (n30807 & n35374);
  assign n35379 = (n30807 & ~n35096) | (n30807 & n35374) | (~n35096 & n35374);
  assign n35380 = (~n29868 & n35378) | (~n29868 & n35379) | (n35378 & n35379);
  assign n30810 = ~n21498 & n35377;
  assign n35381 = ~n21498 & n37382;
  assign n35382 = n21227 & ~n21498;
  assign n35383 = (n35369 & n35381) | (n35369 & n35382) | (n35381 & n35382);
  assign n35384 = (n37347 & n30810) | (n37347 & n35383) | (n30810 & n35383);
  assign n35385 = (n30810 & n35096) | (n30810 & n35383) | (n35096 & n35383);
  assign n35386 = (n29868 & n35384) | (n29868 & n35385) | (n35384 & n35385);
  assign n21501 = n35380 | n35386;
  assign n21503 = n21221 | n21235;
  assign n35387 = (n21235 & n21237) | (n21235 & n21503) | (n21237 & n21503);
  assign n30812 = n21501 | n35387;
  assign n35388 = n21235 | n21501;
  assign n35389 = n21237 | n35388;
  assign n30814 = (n35269 & n30812) | (n35269 & n35389) | (n30812 & n35389);
  assign n21505 = n21236 & n21501;
  assign n30815 = n21503 & n21505;
  assign n30816 = (n21505 & n35269) | (n21505 & n30815) | (n35269 & n30815);
  assign n21507 = n30814 & ~n30816;
  assign n21508 = x134 & x147;
  assign n21509 = n21507 & n21508;
  assign n21510 = n21507 | n21508;
  assign n21511 = ~n21509 & n21510;
  assign n30817 = n21241 | n21511;
  assign n35390 = n30692 | n30817;
  assign n35391 = n30693 | n30817;
  assign n35392 = (n30333 & n35390) | (n30333 & n35391) | (n35390 & n35391);
  assign n21525 = x133 & x148;
  assign n21514 = n30550 | n21241;
  assign n30819 = n21514 | n30567;
  assign n21516 = n21501 & ~n21508;
  assign n21517 = ~n21501 & n21508;
  assign n21518 = n21516 | n21517;
  assign n30822 = n21518 | n35387;
  assign n30795 = n21235 | n21237;
  assign n30823 = n21518 | n30795;
  assign n30824 = (n35269 & n30822) | (n35269 & n30823) | (n30822 & n30823);
  assign n37383 = n21217 & ~n21518;
  assign n37384 = (n21217 & ~n30795) | (n21217 & n37383) | (~n30795 & n37383);
  assign n37385 = (n21217 & ~n35387) | (n21217 & n37383) | (~n35387 & n37383);
  assign n35395 = (~n35269 & n37384) | (~n35269 & n37385) | (n37384 & n37385);
  assign n35396 = n30824 & n35395;
  assign n30825 = n21518 & n35387;
  assign n30826 = n21518 & n30795;
  assign n30827 = (n35269 & n30825) | (n35269 & n30826) | (n30825 & n30826);
  assign n35397 = n30824 & ~n30827;
  assign n35398 = (n21240 & n35396) | (n21240 & n35397) | (n35396 & n35397);
  assign n37386 = n21525 & ~n35398;
  assign n37387 = (n21525 & ~n30819) | (n21525 & n37386) | (~n30819 & n37386);
  assign n35399 = n30566 & n35398;
  assign n35400 = (n21514 & n35398) | (n21514 & n35399) | (n35398 & n35399);
  assign n35402 = n21525 & ~n35400;
  assign n35403 = (~n30333 & n37387) | (~n30333 & n35402) | (n37387 & n35402);
  assign n30834 = n35392 & n35403;
  assign n37388 = ~n21525 & n35398;
  assign n37389 = n30819 & n37388;
  assign n35405 = ~n21525 & n35400;
  assign n35406 = (n30333 & n37389) | (n30333 & n35405) | (n37389 & n35405);
  assign n30836 = (n21525 & n35392) | (n21525 & ~n35406) | (n35392 & ~n35406);
  assign n21528 = ~n30834 & n30836;
  assign n21529 = x132 & x149;
  assign n21530 = n21528 & n21529;
  assign n21531 = n21528 | n21529;
  assign n21532 = ~n21530 & n21531;
  assign n30837 = n21247 | n35361;
  assign n35409 = ~n21532 & n30837;
  assign n35407 = n20993 | n21247;
  assign n35408 = (n21247 & n21249) | (n21247 & n35407) | (n21249 & n35407);
  assign n35410 = ~n21532 & n35408;
  assign n35411 = (n30531 & n35409) | (n30531 & n35410) | (n35409 & n35410);
  assign n35412 = n21532 & ~n30837;
  assign n35413 = n21532 & ~n35408;
  assign n35414 = (~n30531 & n35412) | (~n30531 & n35413) | (n35412 & n35413);
  assign n21536 = n35411 | n35414;
  assign n21537 = x131 & x150;
  assign n21538 = n21536 & n21537;
  assign n21539 = n21536 | n21537;
  assign n21540 = ~n21538 & n21539;
  assign n30840 = n21482 | n21540;
  assign n30841 = n35355 | n30840;
  assign n30842 = n21482 & n21540;
  assign n30843 = (n21540 & n35355) | (n21540 & n30842) | (n35355 & n30842);
  assign n21543 = n30841 & ~n30843;
  assign n21544 = x130 & x151;
  assign n21545 = n21543 | n21544;
  assign n21546 = n21543 & n21544;
  assign n21547 = n21545 & ~n21546;
  assign n30844 = ~n21474 & n21547;
  assign n30845 = ~n30779 & n30844;
  assign n30846 = n21474 & ~n21547;
  assign n30847 = (~n21547 & n30779) | (~n21547 & n30846) | (n30779 & n30846);
  assign n21550 = n30845 | n30847;
  assign n21551 = x129 & x152;
  assign n21552 = n21550 & n21551;
  assign n21553 = n21550 | n21551;
  assign n21554 = ~n21552 & n21553;
  assign n21555 = n30782 | n21554;
  assign n21556 = n30782 & n21554;
  assign n21557 = n21555 & ~n21556;
  assign n21558 = x128 & x153;
  assign n21559 = n21557 | n21558;
  assign n21560 = n21557 & n21558;
  assign n21561 = n21559 & ~n21560;
  assign n30848 = n21196 | n21459;
  assign n30849 = n30639 | n30848;
  assign n35415 = ~n21196 & n21267;
  assign n35416 = (n21267 & ~n21459) | (n21267 & n35415) | (~n21459 & n35415);
  assign n30851 = n21267 & ~n21459;
  assign n30852 = (~n30639 & n35416) | (~n30639 & n30851) | (n35416 & n30851);
  assign n21564 = n30849 & n30852;
  assign n30853 = n21452 | n21564;
  assign n30854 = (n21564 & n30763) | (n21564 & n30853) | (n30763 & n30853);
  assign n21566 = ~n21561 & n30854;
  assign n21567 = n21561 & ~n30854;
  assign n21568 = n21566 | n21567;
  assign n21569 = x127 & x154;
  assign n21570 = n21568 & n21569;
  assign n21571 = n21568 | n21569;
  assign n21572 = ~n21570 & n21571;
  assign n21573 = x126 & x155;
  assign n21574 = n21572 & ~n21573;
  assign n21575 = ~n21572 & n21573;
  assign n21576 = n21574 | n21575;
  assign n21577 = n30766 | n21576;
  assign n21578 = n30766 & n21576;
  assign n21579 = n21577 & ~n21578;
  assign n30753 = (n35233 & n21436) | (n35233 & n30752) | (n21436 & n30752);
  assign n30755 = (n21283 & n30634) | (n21283 & n30754) | (n30634 & n30754);
  assign n35417 = n21182 & n21284;
  assign n35418 = (n21283 & n21284) | (n21283 & n35417) | (n21284 & n35417);
  assign n30759 = (n21284 & n30634) | (n21284 & n35418) | (n30634 & n35418);
  assign n21445 = ~n30755 & n30759;
  assign n30855 = n21445 & n21579;
  assign n30856 = (n21579 & n30753) | (n21579 & n30855) | (n30753 & n30855);
  assign n30857 = n21445 | n21579;
  assign n30858 = n30753 | n30857;
  assign n21582 = ~n30856 & n30858;
  assign n21583 = n21441 & n21582;
  assign n21584 = n21441 | n21582;
  assign n21585 = ~n21583 & n21584;
  assign n21586 = ~n21440 & n21585;
  assign n21587 = n21440 & ~n21585;
  assign n21588 = n21586 | n21587;
  assign n21589 = x124 & x157;
  assign n21590 = n21588 | n21589;
  assign n21591 = n21588 & n21589;
  assign n21592 = n21590 & ~n21591;
  assign n30859 = n21168 | n21429;
  assign n30860 = n30584 | n30859;
  assign n21596 = n21295 & ~n30751;
  assign n21597 = n30860 & n21596;
  assign n21593 = n21156 & n21304;
  assign n30861 = n21593 | n21597;
  assign n30862 = (n21163 & n21597) | (n21163 & n30861) | (n21597 & n30861);
  assign n21599 = n21592 | n30862;
  assign n21600 = n21592 & n30862;
  assign n21601 = n21599 & ~n21600;
  assign n21602 = x123 & x158;
  assign n21603 = n21601 | n21602;
  assign n21604 = n21601 & n21602;
  assign n30868 = n21603 & ~n21604;
  assign n30869 = n21608 & n30868;
  assign n21611 = n21588 | n30862;
  assign n21612 = n21588 & n30862;
  assign n21613 = n21611 & ~n21612;
  assign n21614 = n21589 & n21602;
  assign n21615 = n21589 | n21602;
  assign n21616 = ~n21614 & n21615;
  assign n21617 = n21613 & ~n21616;
  assign n21618 = ~n21613 & n21616;
  assign n21619 = n21617 | n21618;
  assign n21620 = n21608 | n21619;
  assign n21621 = ~n30869 & n21620;
  assign n21622 = x122 & x159;
  assign n21623 = n21621 & n21622;
  assign n21624 = n21621 | n21622;
  assign n21625 = ~n21623 & n21624;
  assign n30870 = n21316 | n21318;
  assign n30871 = (n21154 & n21316) | (n21154 & n30870) | (n21316 & n30870);
  assign n21627 = n21625 | n30871;
  assign n21628 = n21625 & n30871;
  assign n21629 = n21627 & ~n21628;
  assign n21630 = n30749 & n21629;
  assign n21631 = n30749 | n21629;
  assign n21632 = ~n21630 & n21631;
  assign n21633 = n21424 & n21632;
  assign n21634 = n21424 | n21632;
  assign n21635 = ~n21633 & n21634;
  assign n21636 = n35341 & n21635;
  assign n21637 = n35341 | n21635;
  assign n21638 = ~n21636 & n21637;
  assign n21639 = x119 & x162;
  assign n21640 = n21638 | n21639;
  assign n21641 = n21638 & n21639;
  assign n21642 = n21640 & ~n21641;
  assign n21643 = n30745 & n21642;
  assign n21644 = n30745 | n21642;
  assign n21645 = ~n21643 & n21644;
  assign n21646 = x118 & x163;
  assign n21647 = ~n21645 & n21646;
  assign n21648 = n21645 & ~n21646;
  assign n21649 = n21647 | n21648;
  assign n30872 = n21351 & n21352;
  assign n30873 = (n21351 & n30614) | (n21351 & n30872) | (n30614 & n30872);
  assign n21652 = n21649 & ~n30873;
  assign n21653 = ~n21649 & n30873;
  assign n21654 = n21652 | n21653;
  assign n21655 = x117 & x164;
  assign n21656 = n21654 & ~n21655;
  assign n21657 = ~n21654 & n21655;
  assign n21658 = n21656 | n21657;
  assign n21659 = ~n30614 & n21353;
  assign n21660 = n30614 & ~n21353;
  assign n21661 = n21659 | n21660;
  assign n21664 = n21145 | n21661;
  assign n21662 = n21145 & n21661;
  assign n30874 = n21662 & n21664;
  assign n30875 = (n21664 & n30737) | (n21664 & n30874) | (n30737 & n30874);
  assign n21666 = n21658 & ~n30875;
  assign n21667 = ~n21658 & n30875;
  assign n21668 = n21666 | n21667;
  assign n21669 = n30743 & n21668;
  assign n21670 = n30743 | n21668;
  assign n21671 = ~n21669 & n21670;
  assign n21672 = n21408 & n21671;
  assign n21673 = n21408 | n21671;
  assign n21674 = ~n21672 & n21673;
  assign n21675 = n30741 & n21674;
  assign n21676 = n30741 | n21674;
  assign n21677 = ~n21675 & n21676;
  assign n21678 = n21405 | n21677;
  assign n21679 = n21405 & n21677;
  assign n21680 = n21678 & ~n21679;
  assign n21681 = n21387 | n21390;
  assign n21682 = n21386 & n21681;
  assign n21683 = n21680 & ~n21682;
  assign n21684 = ~n21680 & n21682;
  assign n21685 = n21683 | n21684;
  assign n21686 = x114 & x167;
  assign n21687 = n21685 | n21686;
  assign n21688 = n21685 & n21686;
  assign n21689 = n21687 & ~n21688;
  assign n21690 = n21140 | n21396;
  assign n21691 = n21395 & n21690;
  assign n21692 = n21689 & ~n21691;
  assign n21693 = ~n21689 & n21691;
  assign n21694 = n21692 | n21693;
  assign n21695 = x113 & x168;
  assign n21696 = n21694 | n21695;
  assign n21697 = n21694 & n21695;
  assign n21698 = n21696 & ~n21697;
  assign n21699 = ~n21402 & n21698;
  assign n21700 = n21402 & ~n21698;
  assign n21701 = n21699 | n21700;
  assign n21702 = x112 & x169;
  assign n21703 = n21701 & n21702;
  assign n21704 = n21701 | n21702;
  assign n21705 = ~n21703 & n21704;
  assign n21706 = x113 & x169;
  assign n21707 = n21402 | n21697;
  assign n21708 = n21696 & n21707;
  assign n21709 = x116 & x166;
  assign n21717 = n21420 & n21632;
  assign n21718 = n21420 | n21632;
  assign n21719 = ~n21717 & n21718;
  assign n21720 = n35341 & n21719;
  assign n30879 = n21421 & n21719;
  assign n30880 = (n35341 & n21421) | (n35341 & n30879) | (n21421 & n30879);
  assign n21723 = ~n21720 & n30880;
  assign n30881 = n21638 | n21723;
  assign n30882 = (n21723 & n30745) | (n21723 & n30881) | (n30745 & n30881);
  assign n30883 = n21717 | n21719;
  assign n30884 = (n35341 & n21717) | (n35341 & n30883) | (n21717 & n30883);
  assign n21726 = n21621 | n30871;
  assign n30885 = n21153 | n21316;
  assign n30886 = n30616 | n30885;
  assign n21728 = n21317 & n21620;
  assign n21729 = ~n30869 & n21728;
  assign n21730 = n30886 & n21729;
  assign n21731 = n21622 & ~n21730;
  assign n21732 = n21726 & n21731;
  assign n30887 = n21629 | n21732;
  assign n30888 = (n21732 & n30749) | (n21732 & n30887) | (n30749 & n30887);
  assign n30889 = n21601 & n21607;
  assign n30890 = (n21601 & n30725) | (n21601 & n30889) | (n30725 & n30889);
  assign n30891 = n21601 | n21607;
  assign n30892 = n30725 | n30891;
  assign n21736 = n21602 & n30892;
  assign n21737 = ~n30890 & n21736;
  assign n21739 = n21589 & n21613;
  assign n21740 = n30890 | n21739;
  assign n21741 = n21439 | n21582;
  assign n21742 = n30751 | n21741;
  assign n21743 = n21168 | n21439;
  assign n21744 = n30584 | n21743;
  assign n21745 = n21432 & ~n30753;
  assign n21746 = n21291 | n21745;
  assign n21747 = n21582 & n21746;
  assign n30893 = n21441 & ~n21747;
  assign n30894 = (n21441 & ~n21744) | (n21441 & n30893) | (~n21744 & n30893);
  assign n21750 = n21742 & n30894;
  assign n30895 = n21588 | n21750;
  assign n30896 = (n21750 & n30862) | (n21750 & n30895) | (n30862 & n30895);
  assign n21752 = n30766 | n21572;
  assign n21753 = n30766 & n21572;
  assign n21754 = n21752 & ~n21753;
  assign n30897 = n21445 & n21754;
  assign n30898 = (n21754 & n30753) | (n21754 & n30897) | (n30753 & n30897);
  assign n35419 = n21445 & n21573;
  assign n35420 = (n21573 & n21754) | (n21573 & n35419) | (n21754 & n35419);
  assign n30902 = (n21573 & n30753) | (n21573 & n35420) | (n30753 & n35420);
  assign n21758 = ~n30898 & n30902;
  assign n30903 = n21747 | n21758;
  assign n30904 = (n21744 & n21758) | (n21744 & n30903) | (n21758 & n30903);
  assign n21760 = n21455 | n21568;
  assign n30905 = n21760 | n30754;
  assign n30906 = n21283 | n21760;
  assign n30907 = (n30634 & n30905) | (n30634 & n30906) | (n30905 & n30906);
  assign n21764 = n21277 | n21454;
  assign n21765 = n21568 & n21764;
  assign n35421 = n21182 | n21277;
  assign n35422 = (n21182 & n21454) | (n21182 & n35421) | (n21454 & n35421);
  assign n30908 = n35422 & n21765;
  assign n30909 = (n21765 & n30634) | (n21765 & n30908) | (n30634 & n30908);
  assign n21767 = n21569 & ~n30909;
  assign n21768 = n30907 & n21767;
  assign n30910 = n21768 | n30897;
  assign n30911 = n21754 | n21768;
  assign n30912 = (n30753 & n30910) | (n30753 & n30911) | (n30910 & n30911);
  assign n30913 = n21557 & n30853;
  assign n30914 = n21557 & n21564;
  assign n30915 = (n30763 & n30913) | (n30763 & n30914) | (n30913 & n30914);
  assign n30916 = n21557 | n30853;
  assign n30917 = n21557 | n21564;
  assign n30918 = (n30763 & n30916) | (n30763 & n30917) | (n30916 & n30917);
  assign n21772 = n21558 & n30918;
  assign n21773 = ~n30915 & n21772;
  assign n21777 = n30777 & ~n30779;
  assign n21778 = n21208 | n21777;
  assign n21779 = n21550 & n21778;
  assign n21775 = n21196 | n21469;
  assign n30919 = n21775 & n21779;
  assign n30920 = (n21779 & n30639) | (n21779 & n30919) | (n30639 & n30919);
  assign n30921 = n21550 | n30781;
  assign n30922 = n21550 | n30780;
  assign n30923 = (n30639 & n30921) | (n30639 & n30922) | (n30921 & n30922);
  assign n21782 = ~n30920 & n30923;
  assign n21783 = n21551 & n21782;
  assign n30924 = n21474 & n21543;
  assign n35423 = (n21543 & n30778) | (n21543 & n30924) | (n30778 & n30924);
  assign n35424 = (n21466 & n21543) | (n21466 & n30924) | (n21543 & n30924);
  assign n35425 = (n30515 & n35423) | (n30515 & n35424) | (n35423 & n35424);
  assign n30926 = n21474 | n21543;
  assign n30928 = n21544 & n30926;
  assign n35426 = (n21544 & n30778) | (n21544 & n30928) | (n30778 & n30928);
  assign n35427 = (n21466 & n21544) | (n21466 & n30928) | (n21544 & n30928);
  assign n35428 = (n30515 & n35426) | (n30515 & n35427) | (n35426 & n35427);
  assign n21788 = ~n35425 & n35428;
  assign n21790 = x130 & x152;
  assign n30933 = n21212 | n21482;
  assign n35429 = n21203 | n30933;
  assign n35430 = (n30651 & n30933) | (n30651 & n35429) | (n30933 & n35429);
  assign n35431 = (n21200 & n30933) | (n21200 & n35429) | (n30933 & n35429);
  assign n35432 = (n30396 & n35430) | (n30396 & n35431) | (n35430 & n35431);
  assign n30839 = (n30531 & n30837) | (n30531 & n35408) | (n30837 & n35408);
  assign n35434 = n21227 | n21492;
  assign n37390 = n21492 | n37382;
  assign n37391 = (n35376 & n35434) | (n35376 & n37390) | (n35434 & n37390);
  assign n35433 = n21492 | n37382;
  assign n35435 = (n35369 & n35433) | (n35369 & n35434) | (n35433 & n35434);
  assign n35436 = (n37347 & n37391) | (n37347 & n35435) | (n37391 & n35435);
  assign n35437 = (n37391 & n35096) | (n37391 & n35435) | (n35096 & n35435);
  assign n35438 = (n29868 & n35436) | (n29868 & n35437) | (n35436 & n35437);
  assign n21812 = x138 & x144;
  assign n21813 = x137 & x145;
  assign n21814 = n21812 | n21813;
  assign n21815 = n21812 & n21813;
  assign n21816 = n21814 & ~n21815;
  assign n21817 = n21493 & n21816;
  assign n21818 = n35438 & n21817;
  assign n35440 = n21227 & n21494;
  assign n37392 = n21494 & n37382;
  assign n37393 = (n35376 & n35440) | (n35376 & n37392) | (n35440 & n37392);
  assign n35439 = n21494 & n37382;
  assign n35441 = (n35369 & n35439) | (n35369 & n35440) | (n35439 & n35440);
  assign n35442 = (n37347 & n37393) | (n37347 & n35441) | (n37393 & n35441);
  assign n35443 = (n37393 & n35096) | (n37393 & n35441) | (n35096 & n35441);
  assign n35444 = (n29868 & n35442) | (n29868 & n35443) | (n35442 & n35443);
  assign n21819 = n21492 | n21816;
  assign n21820 = n35444 | n21819;
  assign n21821 = ~n21818 & n21820;
  assign n21822 = x136 & x146;
  assign n21823 = n21821 & n21822;
  assign n21824 = n21821 | n21822;
  assign n21825 = ~n21823 & n21824;
  assign n35446 = n21227 | n21494;
  assign n37394 = n21494 | n37382;
  assign n37395 = (n35376 & n35446) | (n35376 & n37394) | (n35446 & n37394);
  assign n35445 = n21494 | n37382;
  assign n35447 = (n35369 & n35445) | (n35369 & n35446) | (n35445 & n35446);
  assign n35448 = (n37347 & n37395) | (n37347 & n35447) | (n37395 & n35447);
  assign n35449 = (n37395 & n35096) | (n37395 & n35447) | (n35096 & n35447);
  assign n35450 = (n29868 & n35448) | (n29868 & n35449) | (n35448 & n35449);
  assign n21808 = n21495 & n35450;
  assign n21809 = ~n35444 & n21808;
  assign n30949 = n21809 | n30815;
  assign n30955 = n21825 & n30949;
  assign n30950 = n21505 | n21809;
  assign n30956 = n21825 & n30950;
  assign n30957 = (n35269 & n30955) | (n35269 & n30956) | (n30955 & n30956);
  assign n30958 = n21825 | n30949;
  assign n30959 = n21825 | n30950;
  assign n30960 = (n35269 & n30958) | (n35269 & n30959) | (n30958 & n30959);
  assign n21828 = ~n30957 & n30960;
  assign n21829 = x135 & x147;
  assign n21830 = n21828 & n21829;
  assign n21831 = n21828 | n21829;
  assign n21832 = ~n21830 & n21831;
  assign n30831 = n35398 & n30819;
  assign n30961 = n21509 & n21832;
  assign n35451 = (n21832 & n30831) | (n21832 & n30961) | (n30831 & n30961);
  assign n35452 = (n21832 & n30961) | (n21832 & n35400) | (n30961 & n35400);
  assign n35453 = (n30333 & n35451) | (n30333 & n35452) | (n35451 & n35452);
  assign n30963 = n21509 | n21832;
  assign n35454 = n30831 | n30963;
  assign n35455 = n30963 | n35400;
  assign n35456 = (n30333 & n35454) | (n30333 & n35455) | (n35454 & n35455);
  assign n21835 = ~n35453 & n35456;
  assign n21836 = x134 & x148;
  assign n21837 = n21835 & n21836;
  assign n21838 = n21835 | n21836;
  assign n21839 = ~n21837 & n21838;
  assign n21840 = x133 & x149;
  assign n21841 = n21839 & n21840;
  assign n21842 = n21839 | n21840;
  assign n21843 = ~n21841 & n21842;
  assign n30941 = n21528 | n30834;
  assign n30965 = n21843 | n30941;
  assign n30966 = n21843 | n30834;
  assign n30967 = (n30839 & n30965) | (n30839 & n30966) | (n30965 & n30966);
  assign n30968 = n21843 & n30941;
  assign n30969 = n21843 & n30834;
  assign n30970 = (n30839 & n30968) | (n30839 & n30969) | (n30968 & n30969);
  assign n21846 = n30967 & ~n30970;
  assign n21847 = x132 & x150;
  assign n21848 = n21846 | n21847;
  assign n21849 = n21846 & n21847;
  assign n21850 = n21848 & ~n21849;
  assign n21793 = n21250 | n21481;
  assign n21794 = n21536 & n21793;
  assign n37396 = n21247 & n21528;
  assign n37397 = (n21528 & n35361) | (n21528 & n37396) | (n35361 & n37396);
  assign n35458 = n21528 & n35408;
  assign n35459 = (n30531 & n37397) | (n30531 & n35458) | (n37397 & n35458);
  assign n37398 = (n21247 & n21529) | (n21247 & n21530) | (n21529 & n21530);
  assign n37400 = (n35361 & n37398) | (n35361 & n21529) | (n37398 & n21529);
  assign n35461 = (n21529 & n21530) | (n21529 & n35408) | (n21530 & n35408);
  assign n35462 = (n30531 & n37400) | (n30531 & n35461) | (n37400 & n35461);
  assign n21802 = ~n35459 & n35462;
  assign n30939 = n21794 | n21802;
  assign n30971 = n21850 & ~n30939;
  assign n30972 = ~n21802 & n21850;
  assign n30973 = (~n35432 & n30971) | (~n35432 & n30972) | (n30971 & n30972);
  assign n30974 = ~n21850 & n30939;
  assign n30975 = n21802 & ~n21850;
  assign n30976 = (n35432 & n30974) | (n35432 & n30975) | (n30974 & n30975);
  assign n21853 = n30973 | n30976;
  assign n21854 = x131 & x151;
  assign n21855 = n21853 & n21854;
  assign n21856 = n21853 | n21854;
  assign n21857 = ~n21855 & n21856;
  assign n30930 = n21482 | n21536;
  assign n30931 = n35355 | n30930;
  assign n21795 = n35432 & n21794;
  assign n21796 = n30931 & ~n21795;
  assign n21797 = n21537 & n21796;
  assign n30936 = n21543 | n21797;
  assign n30977 = n21857 | n30936;
  assign n30935 = n21797 | n30924;
  assign n30978 = n21857 | n30935;
  assign n30979 = (n30779 & n30977) | (n30779 & n30978) | (n30977 & n30978);
  assign n30980 = n21857 & n30936;
  assign n30981 = n21857 & n30935;
  assign n30982 = (n30779 & n30980) | (n30779 & n30981) | (n30980 & n30981);
  assign n21860 = n30979 & ~n30982;
  assign n21861 = n21790 & n21860;
  assign n21862 = n21790 | n21860;
  assign n21863 = ~n21861 & n21862;
  assign n30983 = ~n21788 & n21863;
  assign n30984 = ~n30920 & n30983;
  assign n30985 = n21788 & ~n21863;
  assign n30986 = (~n21863 & n30920) | (~n21863 & n30985) | (n30920 & n30985);
  assign n21866 = n30984 | n30986;
  assign n21867 = x129 & x153;
  assign n21868 = n21866 & n21867;
  assign n21869 = n21866 | n21867;
  assign n21870 = ~n21868 & n21869;
  assign n30987 = ~n21783 & n21870;
  assign n30988 = ~n30915 & n30987;
  assign n30989 = n21783 & ~n21870;
  assign n30990 = (~n21870 & n30915) | (~n21870 & n30989) | (n30915 & n30989);
  assign n21873 = n30988 | n30990;
  assign n21874 = x128 & x154;
  assign n21875 = n21873 | n21874;
  assign n21876 = n21873 & n21874;
  assign n21877 = n21875 & ~n21876;
  assign n30991 = ~n21773 & n21877;
  assign n30992 = ~n30909 & n30991;
  assign n30993 = n21773 & ~n21877;
  assign n30994 = (~n21877 & n30909) | (~n21877 & n30993) | (n30909 & n30993);
  assign n21880 = n30992 | n30994;
  assign n21881 = x127 & x155;
  assign n21882 = n21880 & n21881;
  assign n21883 = n21880 | n21881;
  assign n21884 = ~n21882 & n21883;
  assign n21885 = x126 & x156;
  assign n21886 = n21884 & ~n21885;
  assign n21887 = ~n21884 & n21885;
  assign n21888 = n21886 | n21887;
  assign n21889 = n30912 | n21888;
  assign n21890 = n30912 & n21888;
  assign n21891 = n21889 & ~n21890;
  assign n21892 = ~n30904 & n21891;
  assign n21893 = n30904 & ~n21891;
  assign n21894 = n21892 | n21893;
  assign n21895 = x125 & x157;
  assign n21896 = n21894 & n21895;
  assign n21897 = n21894 | n21895;
  assign n21898 = ~n21896 & n21897;
  assign n21899 = n30896 | n21898;
  assign n21900 = n30896 & n21898;
  assign n21901 = n21899 & ~n21900;
  assign n21902 = x124 & x158;
  assign n21903 = n21901 | n21902;
  assign n21904 = n21901 & n21902;
  assign n21905 = n21903 & ~n21904;
  assign n21906 = n21740 | n21905;
  assign n21907 = n21740 & n21905;
  assign n21908 = n21906 & ~n21907;
  assign n30995 = n21737 | n21908;
  assign n30996 = n21730 | n30995;
  assign n30997 = n21737 & n21908;
  assign n30998 = (n21730 & n21908) | (n21730 & n30997) | (n21908 & n30997);
  assign n21911 = n30996 & ~n30998;
  assign n21912 = x123 & x159;
  assign n21913 = x122 & x160;
  assign n21914 = n21912 & n21913;
  assign n21915 = n21912 | n21913;
  assign n21916 = ~n21914 & n21915;
  assign n21917 = n21911 & n21916;
  assign n21918 = n21911 | n21916;
  assign n21919 = ~n21917 & n21918;
  assign n21920 = n30888 | n21919;
  assign n21921 = n30888 & n21919;
  assign n21922 = n21920 & ~n21921;
  assign n21923 = x121 & x161;
  assign n21924 = n21922 | n21923;
  assign n21925 = n21922 & n21923;
  assign n21926 = n21924 & ~n21925;
  assign n21927 = n30884 | n21926;
  assign n21928 = n30884 & n21926;
  assign n21929 = n21927 & ~n21928;
  assign n21930 = x120 & x162;
  assign n21931 = n21929 | n21930;
  assign n21932 = n21929 & n21930;
  assign n21933 = n21931 & ~n21932;
  assign n21934 = n30882 | n21933;
  assign n21935 = n30882 & n21933;
  assign n21936 = n21934 & ~n21935;
  assign n21937 = x119 & x163;
  assign n21938 = ~n21936 & n21937;
  assign n21939 = n21936 & ~n21937;
  assign n21940 = n21938 | n21939;
  assign n21942 = n30745 | n21638;
  assign n30999 = ~n21638 & n21639;
  assign n31000 = (n21639 & ~n30745) | (n21639 & n30999) | (~n30745 & n30999);
  assign n21944 = n21942 & n31000;
  assign n31001 = n21645 | n21944;
  assign n31002 = (n21944 & n30873) | (n21944 & n31001) | (n30873 & n31001);
  assign n21946 = n21940 & n31002;
  assign n21947 = n21940 | n31002;
  assign n21948 = ~n21946 & n21947;
  assign n21949 = x118 & x164;
  assign n21950 = ~n21948 & n21949;
  assign n21951 = n21948 & ~n21949;
  assign n21952 = n21950 | n21951;
  assign n21941 = n21645 & n30873;
  assign n21953 = n21645 | n30873;
  assign n21954 = ~n21941 & n21953;
  assign n21957 = n21646 | n21954;
  assign n21955 = n21646 & n21954;
  assign n31003 = n21955 & n21957;
  assign n31004 = (n21957 & n30875) | (n21957 & n31003) | (n30875 & n31003);
  assign n21959 = n21952 & ~n31004;
  assign n21960 = ~n21952 & n31004;
  assign n21961 = n21959 | n21960;
  assign n21711 = n21654 | n30875;
  assign n30876 = (n21655 & n21657) | (n21655 & ~n30875) | (n21657 & ~n30875);
  assign n21714 = n21711 & n30876;
  assign n30877 = n21668 | n21714;
  assign n31005 = n21961 | n30877;
  assign n31006 = n21714 | n21961;
  assign n31007 = (n30743 & n31005) | (n30743 & n31006) | (n31005 & n31006);
  assign n31008 = n21961 & n30877;
  assign n31009 = n21714 & n21961;
  assign n31010 = (n30743 & n31008) | (n30743 & n31009) | (n31008 & n31009);
  assign n21964 = n31007 & ~n31010;
  assign n21965 = x117 & x165;
  assign n21966 = n21964 & ~n21965;
  assign n21967 = ~n21964 & n21965;
  assign n21968 = n21966 | n21967;
  assign n31011 = n21672 & n21968;
  assign n31012 = (n21675 & n21968) | (n21675 & n31011) | (n21968 & n31011);
  assign n31013 = n21672 | n21968;
  assign n31014 = n21675 | n31013;
  assign n21971 = ~n31012 & n31014;
  assign n21972 = n21709 | n21971;
  assign n21973 = n21709 & n21971;
  assign n21974 = n21972 & ~n21973;
  assign n31015 = n21678 & n21679;
  assign n31016 = (n21678 & n21682) | (n21678 & n31015) | (n21682 & n31015);
  assign n21977 = n21974 & ~n31016;
  assign n21978 = ~n21974 & n31016;
  assign n21979 = n21977 | n21978;
  assign n21980 = x115 & x167;
  assign n21981 = n21979 | n21980;
  assign n21982 = n21979 & n21980;
  assign n21983 = n21981 & ~n21982;
  assign n31017 = n21687 & n21688;
  assign n31018 = (n21687 & n21691) | (n21687 & n31017) | (n21691 & n31017);
  assign n21986 = n21983 & ~n31018;
  assign n21987 = ~n21983 & n31018;
  assign n21988 = n21986 | n21987;
  assign n21989 = x114 & x168;
  assign n21990 = n21988 | n21989;
  assign n21991 = n21988 & n21989;
  assign n21992 = n21990 & ~n21991;
  assign n21993 = ~n21708 & n21992;
  assign n21994 = n21708 & ~n21992;
  assign n21995 = n21993 | n21994;
  assign n21996 = n21706 & ~n21995;
  assign n21997 = ~n21706 & n21995;
  assign n21998 = n21996 | n21997;
  assign n21999 = ~n21703 & n21998;
  assign n22000 = n21703 & ~n21998;
  assign n22001 = n21999 | n22000;
  assign n22002 = x112 & x170;
  assign n22003 = n22001 & n22002;
  assign n22004 = n22001 | n22002;
  assign n22005 = ~n22003 & n22004;
  assign n22006 = x113 & x170;
  assign n31019 = n21702 & n21706;
  assign n31020 = n21701 & n31019;
  assign n22008 = n21995 | n31020;
  assign n31021 = n21702 | n21706;
  assign n31022 = (n21701 & n21706) | (n21701 & n31021) | (n21706 & n31021);
  assign n22010 = n22008 & n31022;
  assign n22011 = x114 & x169;
  assign n31023 = n21990 & n21991;
  assign n31024 = (n21708 & n21990) | (n21708 & n31023) | (n21990 & n31023);
  assign n22014 = x117 & x166;
  assign n31025 = n21654 | n21955;
  assign n31026 = (n21955 & n30875) | (n21955 & n31025) | (n30875 & n31025);
  assign n22018 = n21948 & n31026;
  assign n31027 = n21948 & n21949;
  assign n31028 = (n21949 & n31026) | (n21949 & n31027) | (n31026 & n31027);
  assign n22021 = ~n22018 & n31028;
  assign n31029 = n21929 & n30881;
  assign n31030 = n21723 & n21929;
  assign n31031 = (n30745 & n31029) | (n30745 & n31030) | (n31029 & n31030);
  assign n35463 = n21922 | n35341;
  assign n35464 = n21717 | n21922;
  assign n35465 = (n30883 & n35463) | (n30883 & n35464) | (n35463 & n35464);
  assign n30747 = n30596 | n35339;
  assign n31032 = n21334 | n21717;
  assign n31033 = (n21717 & n30747) | (n21717 & n31032) | (n30747 & n31032);
  assign n22026 = n21718 & n21922;
  assign n31034 = n21923 & ~n22026;
  assign n31035 = (n21923 & ~n31033) | (n21923 & n31034) | (~n31033 & n31034);
  assign n22029 = n35465 & n31035;
  assign n22030 = n31031 | n22029;
  assign n22031 = n21911 & n21912;
  assign n22032 = n21911 | n21912;
  assign n22033 = ~n22031 & n22032;
  assign n31036 = n22031 | n22033;
  assign n31037 = (n22031 & n30888) | (n22031 & n31036) | (n30888 & n31036);
  assign n31038 = n21739 & n21901;
  assign n31039 = (n21901 & n30890) | (n21901 & n31038) | (n30890 & n31038);
  assign n31040 = n21739 | n21901;
  assign n31041 = n30890 | n31040;
  assign n22038 = n21902 & n31041;
  assign n22039 = ~n31039 & n22038;
  assign n22041 = n21750 | n21894;
  assign n31042 = n21588 | n22041;
  assign n31043 = (n22041 & n30862) | (n22041 & n31042) | (n30862 & n31042);
  assign n22043 = n21597 | n21750;
  assign n31044 = n21593 | n22043;
  assign n31045 = (n21163 & n22043) | (n21163 & n31044) | (n22043 & n31044);
  assign n21748 = n21744 & n21747;
  assign n22045 = n21742 & ~n21748;
  assign n22046 = n21441 | n22045;
  assign n22047 = n21894 & n22046;
  assign n22048 = n31045 & n22047;
  assign n22049 = n31043 & ~n22048;
  assign n22050 = n21895 & n22049;
  assign n22051 = n31039 | n22050;
  assign n22052 = x125 & x158;
  assign n22053 = n30912 | n21884;
  assign n22054 = n30912 & n21884;
  assign n22055 = n22053 & ~n22054;
  assign n22056 = n30904 & n22055;
  assign n31046 = n21885 & n22055;
  assign n31047 = (n21885 & n30904) | (n21885 & n31046) | (n30904 & n31046);
  assign n22059 = ~n22056 & n31047;
  assign n31048 = n22047 | n22059;
  assign n31049 = (n22059 & n31045) | (n22059 & n31048) | (n31045 & n31048);
  assign n22061 = n30912 | n21880;
  assign n22064 = n30907 & ~n30909;
  assign n22065 = n21569 | n22064;
  assign n22066 = n21880 & n22065;
  assign n22062 = n21445 | n21768;
  assign n31050 = n22062 & n22066;
  assign n31051 = (n22066 & n30753) | (n22066 & n31050) | (n30753 & n31050);
  assign n31052 = n21881 & ~n31051;
  assign n31053 = n22061 & n31052;
  assign n31054 = n22055 | n31053;
  assign n31055 = (n30904 & n31053) | (n30904 & n31054) | (n31053 & n31054);
  assign n22072 = n21783 | n21866;
  assign n22073 = n30915 | n22072;
  assign n31058 = n21783 | n30853;
  assign n31059 = n21564 | n21783;
  assign n31060 = (n30763 & n31058) | (n30763 & n31059) | (n31058 & n31059);
  assign n22075 = n21551 | n21782;
  assign n22076 = n21866 & n22075;
  assign n22077 = n31060 & n22076;
  assign n22078 = n22073 & ~n22077;
  assign n22079 = n21867 & n22078;
  assign n31056 = n21773 & n21873;
  assign n31061 = n22079 | n31056;
  assign n31062 = n21873 | n22079;
  assign n31063 = (n30909 & n31061) | (n30909 & n31062) | (n31061 & n31062);
  assign n22083 = n21537 | n21796;
  assign n22084 = n21853 & n22083;
  assign n31066 = n21474 | n21797;
  assign n31068 = n22084 & n31066;
  assign n31069 = (n22084 & n30779) | (n22084 & n31068) | (n30779 & n31068);
  assign n35466 = n21543 | n21853;
  assign n35467 = n21797 | n35466;
  assign n31071 = n21853 | n30935;
  assign n31072 = (n30779 & n35467) | (n30779 & n31071) | (n35467 & n31071);
  assign n22087 = ~n31069 & n31072;
  assign n22088 = n21854 & n22087;
  assign n31064 = n21788 & n21860;
  assign n31073 = n22088 | n31064;
  assign n31074 = n21860 | n22088;
  assign n31075 = (n30920 & n31073) | (n30920 & n31074) | (n31073 & n31074);
  assign n31076 = n21846 & n30939;
  assign n31077 = n21802 & n21846;
  assign n31078 = (n35432 & n31076) | (n35432 & n31077) | (n31076 & n31077);
  assign n37401 = (n21847 & n21849) | (n21847 & n30939) | (n21849 & n30939);
  assign n37402 = n21802 & n21847;
  assign n37403 = (n21846 & n21847) | (n21846 & n37402) | (n21847 & n37402);
  assign n35470 = (n35432 & n37401) | (n35432 & n37403) | (n37401 & n37403);
  assign n22093 = ~n31078 & n35470;
  assign n22095 = n30834 | n21839;
  assign n35471 = n21839 | n30941;
  assign n35472 = (n22095 & n30837) | (n22095 & n35471) | (n30837 & n35471);
  assign n35473 = (n22095 & n35408) | (n22095 & n35471) | (n35408 & n35471);
  assign n35474 = (n30531 & n35472) | (n30531 & n35473) | (n35472 & n35473);
  assign n22099 = n30836 & n21839;
  assign n22097 = n21247 | n30834;
  assign n31085 = n21478 | n22097;
  assign n35475 = n22099 & n31085;
  assign n31084 = n22097 | n35361;
  assign n35476 = n22099 & n31084;
  assign n35477 = (n30531 & n35475) | (n30531 & n35476) | (n35475 & n35476);
  assign n22101 = n35474 & ~n35477;
  assign n22102 = n21840 & n22101;
  assign n31086 = (n30531 & n31084) | (n30531 & n31085) | (n31084 & n31085);
  assign n22106 = x139 & x144;
  assign n22107 = x138 & x145;
  assign n22108 = n22106 & n22107;
  assign n22109 = n22106 | n22107;
  assign n22110 = ~n22108 & n22109;
  assign n22111 = x137 & x146;
  assign n22112 = n22110 & n22111;
  assign n22113 = n22110 | n22111;
  assign n22114 = ~n22112 & n22113;
  assign n35480 = n21493 | n21815;
  assign n35481 = (n21815 & n21816) | (n21815 & n35480) | (n21816 & n35480);
  assign n31092 = n22114 & ~n35481;
  assign n31093 = ~n21815 & n22114;
  assign n31094 = (~n35438 & n31092) | (~n35438 & n31093) | (n31092 & n31093);
  assign n31095 = ~n22114 & n35481;
  assign n31096 = n21815 & ~n22114;
  assign n31097 = (n35438 & n31095) | (n35438 & n31096) | (n31095 & n31096);
  assign n22117 = n31094 | n31097;
  assign n37404 = n21823 | n22117;
  assign n37405 = n30956 | n37404;
  assign n35478 = n21823 | n21825;
  assign n35479 = (n21823 & n30949) | (n21823 & n35478) | (n30949 & n35478);
  assign n35483 = n22117 | n35479;
  assign n35484 = (n35269 & n37405) | (n35269 & n35483) | (n37405 & n35483);
  assign n22124 = x136 & x147;
  assign n22119 = n21809 | n21823;
  assign n31098 = n22119 | n30815;
  assign n22133 = ~n22117 & n22124;
  assign n37743 = (~n21824 & n22124) | (~n21824 & n22133) | (n22124 & n22133);
  assign n37407 = (n22124 & ~n31098) | (n22124 & n37743) | (~n31098 & n37743);
  assign n31099 = n21505 | n22119;
  assign n37408 = (n22124 & ~n31099) | (n22124 & n37743) | (~n31099 & n37743);
  assign n35487 = (~n35269 & n37407) | (~n35269 & n37408) | (n37407 & n37408);
  assign n31105 = n35484 & n35487;
  assign n22132 = n22117 & ~n22124;
  assign n37744 = n21824 & n22132;
  assign n37410 = n31098 & n37744;
  assign n37411 = n31099 & n37744;
  assign n35490 = (n35269 & n37410) | (n35269 & n37411) | (n37410 & n37411);
  assign n31107 = (n35484 & n22124) | (n35484 & ~n35490) | (n22124 & ~n35490);
  assign n22127 = ~n31105 & n31107;
  assign n22130 = n21509 | n21830;
  assign n35491 = (n21830 & n21832) | (n21830 & n22130) | (n21832 & n22130);
  assign n31111 = n22127 | n35491;
  assign n35492 = n21830 | n22127;
  assign n35493 = n21832 | n35492;
  assign n35494 = (n30831 & n31111) | (n30831 & n35493) | (n31111 & n35493);
  assign n35495 = (n31111 & n35400) | (n31111 & n35493) | (n35400 & n35493);
  assign n35496 = (n30333 & n35494) | (n30333 & n35495) | (n35494 & n35495);
  assign n22134 = n22132 | n22133;
  assign n37412 = n21823 | n22134;
  assign n37413 = n30956 | n37412;
  assign n35498 = n22134 | n35479;
  assign n35499 = (n35269 & n37413) | (n35269 & n35498) | (n37413 & n35498);
  assign n37414 = n21823 & n22134;
  assign n37415 = (n22134 & n30956) | (n22134 & n37414) | (n30956 & n37414);
  assign n35501 = n22134 & n35479;
  assign n35502 = (n35269 & n37415) | (n35269 & n35501) | (n37415 & n35501);
  assign n31114 = n35499 & ~n35502;
  assign n31115 = n21831 & n31114;
  assign n31116 = n22130 & n31115;
  assign n35503 = (n30831 & n31115) | (n30831 & n31116) | (n31115 & n31116);
  assign n35504 = (n31115 & n31116) | (n31115 & n35400) | (n31116 & n35400);
  assign n35505 = (n30333 & n35503) | (n30333 & n35504) | (n35503 & n35504);
  assign n22140 = n35496 & ~n35505;
  assign n22141 = x135 & x148;
  assign n22142 = n22140 & n22141;
  assign n22143 = n22140 | n22141;
  assign n22144 = ~n22142 & n22143;
  assign n22145 = x134 & x149;
  assign n22146 = n22144 & n22145;
  assign n22147 = n22144 | n22145;
  assign n22148 = ~n22146 & n22147;
  assign n35506 = n21837 | n30836;
  assign n35507 = (n21837 & n21839) | (n21837 & n35506) | (n21839 & n35506);
  assign n31120 = ~n22148 & n35507;
  assign n31121 = n21837 & ~n22148;
  assign n31122 = (n31086 & n31120) | (n31086 & n31121) | (n31120 & n31121);
  assign n31123 = n22148 & ~n35507;
  assign n31124 = ~n21837 & n22148;
  assign n31125 = (~n31086 & n31123) | (~n31086 & n31124) | (n31123 & n31124);
  assign n22152 = n31122 | n31125;
  assign n22153 = x133 & x150;
  assign n22154 = n22152 & n22153;
  assign n22155 = n22152 | n22153;
  assign n22156 = ~n22154 & n22155;
  assign n31126 = n22102 | n22156;
  assign n31127 = n31078 | n31126;
  assign n31128 = n22102 & n22156;
  assign n31129 = (n22156 & n31078) | (n22156 & n31128) | (n31078 & n31128);
  assign n22159 = n31127 & ~n31129;
  assign n22160 = x132 & x151;
  assign n22161 = n22159 | n22160;
  assign n22162 = n22159 & n22160;
  assign n22163 = n22161 & ~n22162;
  assign n31130 = ~n22093 & n22163;
  assign n31131 = ~n31069 & n31130;
  assign n31132 = n22093 & ~n22163;
  assign n31133 = (~n22163 & n31069) | (~n22163 & n31132) | (n31069 & n31132);
  assign n22166 = n31131 | n31133;
  assign n22167 = x131 & x152;
  assign n22168 = n22166 & n22167;
  assign n22169 = n22166 | n22167;
  assign n22170 = ~n22168 & n22169;
  assign n22171 = n31075 | n22170;
  assign n22172 = n31075 & n22170;
  assign n22173 = n22171 & ~n22172;
  assign n22174 = x130 & x153;
  assign n22175 = n22173 | n22174;
  assign n22176 = n22173 & n22174;
  assign n22177 = n22175 & ~n22176;
  assign n31134 = n21788 | n21860;
  assign n31135 = n30920 | n31134;
  assign n35508 = ~n21788 & n21790;
  assign n35509 = (n21790 & ~n21860) | (n21790 & n35508) | (~n21860 & n35508);
  assign n31137 = n21790 & ~n21860;
  assign n31138 = (~n30920 & n35509) | (~n30920 & n31137) | (n35509 & n31137);
  assign n22180 = n31135 & n31138;
  assign n31139 = n22076 | n22180;
  assign n31140 = (n22180 & n31060) | (n22180 & n31139) | (n31060 & n31139);
  assign n22182 = ~n22177 & n31140;
  assign n22183 = n22177 & ~n31140;
  assign n22184 = n22182 | n22183;
  assign n22185 = x129 & x154;
  assign n22186 = n22184 & n22185;
  assign n22187 = n22184 | n22185;
  assign n22188 = ~n22186 & n22187;
  assign n22189 = n31063 | n22188;
  assign n22190 = n31063 & n22188;
  assign n22191 = n22189 & ~n22190;
  assign n22192 = x128 & x155;
  assign n22193 = n22191 | n22192;
  assign n22194 = n22191 & n22192;
  assign n22195 = n22193 & ~n22194;
  assign n31141 = n21773 | n21873;
  assign n31142 = n30909 | n31141;
  assign n31143 = n21874 & ~n31056;
  assign n31144 = ~n21873 & n21874;
  assign n31145 = (~n30909 & n31143) | (~n30909 & n31144) | (n31143 & n31144);
  assign n22198 = n31142 & n31145;
  assign n22199 = n31051 | n22198;
  assign n22200 = ~n22195 & n22199;
  assign n22201 = n22195 & ~n22199;
  assign n22202 = n22200 | n22201;
  assign n22203 = x127 & x156;
  assign n22204 = n22202 & n22203;
  assign n22205 = n22202 | n22203;
  assign n22206 = ~n22204 & n22205;
  assign n22207 = n31055 | n22206;
  assign n22208 = n31055 & n22206;
  assign n22209 = n22207 & ~n22208;
  assign n22210 = x126 & x157;
  assign n22211 = ~n22209 & n22210;
  assign n22212 = n22209 & ~n22210;
  assign n22213 = n22211 | n22212;
  assign n22214 = n31049 | n22213;
  assign n22215 = n31049 & n22213;
  assign n22216 = n22214 & ~n22215;
  assign n22217 = n22052 & n22216;
  assign n22218 = n22052 | n22216;
  assign n22219 = ~n22217 & n22218;
  assign n22220 = ~n22051 & n22219;
  assign n22221 = n22051 & ~n22219;
  assign n22222 = n22220 | n22221;
  assign n31146 = n22039 | n22222;
  assign n31147 = n30998 | n31146;
  assign n31148 = n22039 & n22222;
  assign n31149 = (n22222 & n30998) | (n22222 & n31148) | (n30998 & n31148);
  assign n22225 = n31147 & ~n31149;
  assign n22226 = x124 & x159;
  assign n22227 = x123 & x160;
  assign n22228 = n22226 & n22227;
  assign n22229 = n22226 | n22227;
  assign n22230 = ~n22228 & n22229;
  assign n22231 = n22225 & n22230;
  assign n22232 = n22225 | n22230;
  assign n22233 = ~n22231 & n22232;
  assign n22234 = n31037 | n22233;
  assign n22235 = n31037 & n22233;
  assign n22236 = n22234 & ~n22235;
  assign n22237 = x122 & x161;
  assign n22238 = n22236 | n22237;
  assign n22239 = n22236 & n22237;
  assign n22240 = n22238 & ~n22239;
  assign n22241 = n30888 | n22033;
  assign n31150 = n21913 & ~n22033;
  assign n31151 = (n21913 & ~n30888) | (n21913 & n31150) | (~n30888 & n31150);
  assign n22243 = n22241 & n31151;
  assign n31152 = n22026 | n22243;
  assign n31153 = (n22243 & n31033) | (n22243 & n31152) | (n31033 & n31152);
  assign n22245 = n22240 | n31153;
  assign n22246 = n22240 & n31153;
  assign n22247 = n22245 & ~n22246;
  assign n22248 = x121 & x162;
  assign n22249 = n22247 | n22248;
  assign n22250 = n22247 & n22248;
  assign n22251 = n22249 & ~n22250;
  assign n22252 = n22030 | n22251;
  assign n22253 = n22030 & n22251;
  assign n22254 = n22252 & ~n22253;
  assign n22255 = x120 & x163;
  assign n22256 = ~n22254 & n22255;
  assign n22257 = n22254 & ~n22255;
  assign n22258 = n22256 | n22257;
  assign n31154 = n21936 & n31001;
  assign n31155 = n21936 & n21944;
  assign n31156 = (n30873 & n31154) | (n30873 & n31155) | (n31154 & n31155);
  assign n31157 = n21929 | n30881;
  assign n31158 = n21723 | n21929;
  assign n31159 = (n30745 & n31157) | (n30745 & n31158) | (n31157 & n31158);
  assign n22261 = n21930 & ~n31031;
  assign n22262 = n31159 & n22261;
  assign n22263 = n31156 | n22262;
  assign n22264 = n22258 & n22263;
  assign n22265 = n22258 | n22263;
  assign n22266 = ~n22264 & n22265;
  assign n22267 = x119 & x164;
  assign n22268 = ~n22266 & n22267;
  assign n22269 = n22266 & ~n22267;
  assign n22270 = n22268 | n22269;
  assign n31160 = n21936 | n31001;
  assign n31161 = n21936 | n21944;
  assign n31162 = (n30873 & n31160) | (n30873 & n31161) | (n31160 & n31161);
  assign n22272 = n21937 & ~n31156;
  assign n22273 = n31162 & n22272;
  assign n31163 = n21948 | n22273;
  assign n31164 = (n22273 & n31026) | (n22273 & n31163) | (n31026 & n31163);
  assign n22275 = n22270 & n31164;
  assign n22276 = n22270 | n31164;
  assign n22277 = ~n22275 & n22276;
  assign n31165 = ~n22021 & n22277;
  assign n31166 = ~n31010 & n31165;
  assign n31167 = n22021 & ~n22277;
  assign n31168 = (~n22277 & n31010) | (~n22277 & n31167) | (n31010 & n31167);
  assign n22280 = n31166 | n31168;
  assign n22281 = x118 & x165;
  assign n22282 = n22280 & n22281;
  assign n22283 = n22280 | n22281;
  assign n22284 = ~n22282 & n22283;
  assign n22015 = n21964 & n21965;
  assign n31169 = n22015 & n22284;
  assign n31170 = (n22284 & n31012) | (n22284 & n31169) | (n31012 & n31169);
  assign n31171 = n22015 | n22284;
  assign n31172 = n31012 | n31171;
  assign n22287 = ~n31170 & n31172;
  assign n22288 = n22014 | n22287;
  assign n22289 = n22014 & n22287;
  assign n22290 = n22288 & ~n22289;
  assign n31173 = n21972 & n21973;
  assign n31174 = (n21972 & n31016) | (n21972 & n31173) | (n31016 & n31173);
  assign n22293 = n22290 & ~n31174;
  assign n22294 = ~n22290 & n31174;
  assign n22295 = n22293 | n22294;
  assign n22296 = x116 & x167;
  assign n22297 = n22295 | n22296;
  assign n22298 = n22295 & n22296;
  assign n22299 = n22297 & ~n22298;
  assign n31175 = n21981 & n21982;
  assign n31176 = (n21981 & n31018) | (n21981 & n31175) | (n31018 & n31175);
  assign n22302 = n22299 & ~n31176;
  assign n22303 = ~n22299 & n31176;
  assign n22304 = n22302 | n22303;
  assign n22305 = x115 & x168;
  assign n22306 = n22304 | n22305;
  assign n22307 = n22304 & n22305;
  assign n22308 = n22306 & ~n22307;
  assign n22309 = ~n31024 & n22308;
  assign n22310 = n31024 & ~n22308;
  assign n22311 = n22309 | n22310;
  assign n22312 = n22011 & n22311;
  assign n22313 = n22011 | n22311;
  assign n22314 = ~n22312 & n22313;
  assign n22315 = n22010 & n22314;
  assign n22316 = n22010 | n22314;
  assign n22317 = ~n22315 & n22316;
  assign n22318 = n22006 | n22317;
  assign n22319 = n22006 & n22317;
  assign n22320 = n22318 & ~n22319;
  assign n22321 = ~n22003 & n22320;
  assign n22322 = n22003 & ~n22320;
  assign n22323 = n22321 | n22322;
  assign n22324 = x112 & x171;
  assign n22325 = n22323 & n22324;
  assign n22326 = n22323 | n22324;
  assign n22327 = ~n22325 & n22326;
  assign n22328 = x113 & x171;
  assign n22329 = x118 & x166;
  assign n31177 = n22021 & n22277;
  assign n31178 = (n22277 & n31010) | (n22277 & n31177) | (n31010 & n31177);
  assign n31179 = n22266 & n31163;
  assign n31180 = n22266 & n22273;
  assign n31181 = (n31026 & n31179) | (n31026 & n31180) | (n31179 & n31180);
  assign n31182 = n22266 | n31163;
  assign n31183 = n22266 | n22273;
  assign n31184 = (n31026 & n31182) | (n31026 & n31183) | (n31182 & n31183);
  assign n22334 = n22267 & n31184;
  assign n22335 = ~n31181 & n22334;
  assign n22338 = n22236 & n31153;
  assign n31187 = (n22237 & n22239) | (n22237 & n31153) | (n22239 & n31153);
  assign n22341 = ~n22338 & n31187;
  assign n31185 = n22029 & n22247;
  assign n31188 = n22341 | n31185;
  assign n31189 = n22247 | n22341;
  assign n31190 = (n31031 & n31188) | (n31031 & n31189) | (n31188 & n31189);
  assign n22343 = n22225 & n22226;
  assign n22344 = n22225 | n22226;
  assign n22345 = ~n22343 & n22344;
  assign n31191 = n22343 | n22345;
  assign n31192 = (n22343 & n31037) | (n22343 & n31191) | (n31037 & n31191);
  assign n22348 = n22050 | n22216;
  assign n22349 = n31039 | n22348;
  assign n22350 = n21739 | n22050;
  assign n22351 = n30890 | n22350;
  assign n22352 = n21895 | n22049;
  assign n22353 = n22216 & n22352;
  assign n31193 = n22052 & ~n22353;
  assign n31194 = (n22052 & ~n22351) | (n22052 & n31193) | (~n22351 & n31193);
  assign n22356 = n22349 & n31194;
  assign n22357 = n31149 | n22356;
  assign n22358 = n31049 & n22209;
  assign n31195 = n22209 & n22210;
  assign n31196 = (n22210 & n31049) | (n22210 & n31195) | (n31049 & n31195);
  assign n22361 = ~n22358 & n31196;
  assign n31197 = n22353 | n22361;
  assign n31198 = (n22351 & n22361) | (n22351 & n31197) | (n22361 & n31197);
  assign n22364 = n30904 | n31053;
  assign n31202 = ~n21881 & n31051;
  assign n31203 = (n21881 & n22061) | (n21881 & ~n31202) | (n22061 & ~n31202);
  assign n22366 = n22202 & n31203;
  assign n22367 = n22364 & n22366;
  assign n31199 = n22202 | n31054;
  assign n31200 = n22202 | n31053;
  assign n31201 = (n30904 & n31199) | (n30904 & n31200) | (n31199 & n31200);
  assign n31204 = n22203 & n31201;
  assign n31205 = ~n22367 & n31204;
  assign n31206 = n22209 | n31205;
  assign n31207 = (n31049 & n31205) | (n31049 & n31206) | (n31205 & n31206);
  assign n31208 = n22191 & n22198;
  assign n31209 = (n22191 & n31051) | (n22191 & n31208) | (n31051 & n31208);
  assign n35510 = n22192 & n22198;
  assign n35511 = (n22191 & n22192) | (n22191 & n35510) | (n22192 & n35510);
  assign n31213 = (n22192 & n31051) | (n22192 & n35511) | (n31051 & n35511);
  assign n22374 = ~n31209 & n31213;
  assign n35512 = n22374 | n31203;
  assign n35513 = (n22202 & n22374) | (n22202 & n35512) | (n22374 & n35512);
  assign n31215 = (n22364 & n22374) | (n22364 & n35513) | (n22374 & n35513);
  assign n22378 = n21867 | n22078;
  assign n22379 = n22184 & n22378;
  assign n22376 = n21773 | n22079;
  assign n31216 = n22376 & n22379;
  assign n31217 = (n22379 & n30909) | (n22379 & n31216) | (n30909 & n31216);
  assign n31218 = n22184 | n31062;
  assign n31219 = n22184 | n31061;
  assign n31220 = (n30909 & n31218) | (n30909 & n31219) | (n31218 & n31219);
  assign n22382 = ~n31217 & n31220;
  assign n22383 = n22185 & n22382;
  assign n31221 = n22383 | n31208;
  assign n31222 = n22191 | n22383;
  assign n31223 = (n31051 & n31221) | (n31051 & n31222) | (n31221 & n31222);
  assign n31224 = n22173 & n31139;
  assign n31225 = n22173 & n22180;
  assign n31226 = (n31060 & n31224) | (n31060 & n31225) | (n31224 & n31225);
  assign n31227 = n22173 | n31139;
  assign n31228 = n22173 | n22180;
  assign n31229 = (n31060 & n31227) | (n31060 & n31228) | (n31227 & n31228);
  assign n22387 = n22174 & n31229;
  assign n22388 = ~n31226 & n22387;
  assign n31230 = n22166 | n31074;
  assign n31231 = n22166 | n31073;
  assign n31232 = (n30920 & n31230) | (n30920 & n31231) | (n31230 & n31231);
  assign n22392 = n21854 | n22087;
  assign n22393 = n22166 & n22392;
  assign n35514 = n21788 | n21854;
  assign n35515 = (n21788 & n22087) | (n21788 & n35514) | (n22087 & n35514);
  assign n31235 = n22393 & n35515;
  assign n31236 = (n22393 & n30920) | (n22393 & n31235) | (n30920 & n31235);
  assign n22395 = n31232 & ~n31236;
  assign n22396 = n22167 & n22395;
  assign n31237 = n22093 & n22159;
  assign n35516 = (n22159 & n31068) | (n22159 & n31237) | (n31068 & n31237);
  assign n35517 = (n22084 & n22159) | (n22084 & n31237) | (n22159 & n31237);
  assign n35518 = (n30779 & n35516) | (n30779 & n35517) | (n35516 & n35517);
  assign n35519 = n22093 & n22160;
  assign n35520 = (n22159 & n22160) | (n22159 & n35519) | (n22160 & n35519);
  assign n35521 = (n22160 & n31068) | (n22160 & n35520) | (n31068 & n35520);
  assign n35522 = (n22084 & n22160) | (n22084 & n35520) | (n22160 & n35520);
  assign n35523 = (n30779 & n35521) | (n30779 & n35522) | (n35521 & n35522);
  assign n22401 = ~n35518 & n35523;
  assign n22405 = n21802 | n22102;
  assign n31243 = n21794 | n22405;
  assign n31244 = (n22405 & n35432) | (n22405 & n31243) | (n35432 & n31243);
  assign n31248 = n22144 & n35507;
  assign n31249 = n21837 & n22144;
  assign n35524 = (n31085 & n31248) | (n31085 & n31249) | (n31248 & n31249);
  assign n35525 = (n31084 & n31248) | (n31084 & n31249) | (n31248 & n31249);
  assign n35526 = (n30531 & n35524) | (n30531 & n35525) | (n35524 & n35525);
  assign n22426 = x140 & x144;
  assign n22427 = x139 & x145;
  assign n22428 = n22426 | n22427;
  assign n22429 = n22426 & n22427;
  assign n22430 = n22428 & ~n22429;
  assign n22431 = n22109 & n22430;
  assign n31271 = n22108 | n35481;
  assign n31274 = n22431 & n31271;
  assign n31272 = n21815 | n22108;
  assign n31275 = n22431 & n31272;
  assign n31276 = (n35438 & n31274) | (n35438 & n31275) | (n31274 & n31275);
  assign n22433 = n22108 | n22430;
  assign n31259 = n22110 & n35481;
  assign n31277 = n22433 | n31259;
  assign n31260 = n21815 & n22110;
  assign n31278 = n22433 | n31260;
  assign n31279 = (n35438 & n31277) | (n35438 & n31278) | (n31277 & n31278);
  assign n22435 = ~n31276 & n31279;
  assign n22436 = x138 & x146;
  assign n22437 = n22435 & n22436;
  assign n22438 = n22435 | n22436;
  assign n22439 = ~n22437 & n22438;
  assign n31261 = (n35438 & n31259) | (n35438 & n31260) | (n31259 & n31260);
  assign n35527 = (n22111 & n22112) | (n22111 & n35481) | (n22112 & n35481);
  assign n35528 = n21815 & n22111;
  assign n35529 = (n22110 & n22111) | (n22110 & n35528) | (n22111 & n35528);
  assign n31267 = (n35438 & n35527) | (n35438 & n35529) | (n35527 & n35529);
  assign n22423 = ~n31261 & n31267;
  assign n37416 = n22117 | n22423;
  assign n37417 = (n21824 & n22423) | (n21824 & n37416) | (n22423 & n37416);
  assign n37418 = n22439 & n37417;
  assign n37419 = n22423 & n22439;
  assign n37420 = (n31099 & n37418) | (n31099 & n37419) | (n37418 & n37419);
  assign n37421 = (n31098 & n37418) | (n31098 & n37419) | (n37418 & n37419);
  assign n35535 = (n35269 & n37420) | (n35269 & n37421) | (n37420 & n37421);
  assign n37422 = n22439 | n37417;
  assign n37423 = n22423 | n22439;
  assign n37424 = (n31099 & n37422) | (n31099 & n37423) | (n37422 & n37423);
  assign n37425 = (n31098 & n37422) | (n31098 & n37423) | (n37422 & n37423);
  assign n35538 = (n35269 & n37424) | (n35269 & n37425) | (n37424 & n37425);
  assign n22442 = ~n35535 & n35538;
  assign n22443 = x137 & x147;
  assign n22444 = n22442 & n22443;
  assign n22445 = n22442 | n22443;
  assign n22446 = ~n22444 & n22445;
  assign n35541 = n31105 | n31114;
  assign n35542 = (n21831 & n31105) | (n21831 & n35541) | (n31105 & n35541);
  assign n31281 = n22446 & n35542;
  assign n35539 = n22446 & n31105;
  assign n35540 = (n22446 & n31116) | (n22446 & n35539) | (n31116 & n35539);
  assign n35543 = (n30831 & n31281) | (n30831 & n35540) | (n31281 & n35540);
  assign n35544 = (n31281 & n35400) | (n31281 & n35540) | (n35400 & n35540);
  assign n35545 = (n30333 & n35543) | (n30333 & n35544) | (n35543 & n35544);
  assign n31284 = n22446 | n35542;
  assign n35546 = n22446 | n31105;
  assign n35547 = n31116 | n35546;
  assign n35548 = (n30831 & n31284) | (n30831 & n35547) | (n31284 & n35547);
  assign n35549 = (n31284 & n35400) | (n31284 & n35547) | (n35400 & n35547);
  assign n35550 = (n30333 & n35548) | (n30333 & n35549) | (n35548 & n35549);
  assign n22449 = ~n35545 & n35550;
  assign n22450 = x136 & x148;
  assign n22451 = n22449 & n22450;
  assign n22452 = n22449 | n22450;
  assign n22453 = ~n22451 & n22452;
  assign n22454 = x135 & x149;
  assign n22455 = n22453 & n22454;
  assign n22456 = n22453 | n22454;
  assign n22457 = ~n22455 & n22456;
  assign n31286 = ~n22142 & n22457;
  assign n31287 = ~n35526 & n31286;
  assign n31288 = n22142 & ~n22457;
  assign n31289 = (~n22457 & n35526) | (~n22457 & n31288) | (n35526 & n31288);
  assign n22460 = n31287 | n31289;
  assign n22461 = x134 & x150;
  assign n22462 = n22460 | n22461;
  assign n22463 = n22460 & n22461;
  assign n22464 = n22462 & ~n22463;
  assign n22407 = n21840 | n22101;
  assign n22408 = n22152 & n22407;
  assign n31251 = n22144 | n35507;
  assign n31252 = n21837 | n22144;
  assign n35551 = (n31085 & n31251) | (n31085 & n31252) | (n31251 & n31252);
  assign n35552 = (n31084 & n31251) | (n31084 & n31252) | (n31251 & n31252);
  assign n35553 = (n30531 & n35551) | (n30531 & n35552) | (n35551 & n35552);
  assign n22415 = n22145 & n35553;
  assign n22416 = ~n35526 & n22415;
  assign n31254 = n22408 | n22416;
  assign n31290 = n22464 & ~n31254;
  assign n31291 = ~n22416 & n22464;
  assign n31292 = (~n31244 & n31290) | (~n31244 & n31291) | (n31290 & n31291);
  assign n31293 = ~n22464 & n31254;
  assign n31294 = n22416 & ~n22464;
  assign n31295 = (n31244 & n31293) | (n31244 & n31294) | (n31293 & n31294);
  assign n22467 = n31292 | n31295;
  assign n22468 = x133 & x151;
  assign n22469 = n22467 & n22468;
  assign n22470 = n22467 | n22468;
  assign n22471 = ~n22469 & n22470;
  assign n22403 = n22102 | n22152;
  assign n35554 = n22403 | n31076;
  assign n35555 = n22403 | n31077;
  assign n35556 = (n35432 & n35554) | (n35432 & n35555) | (n35554 & n35555);
  assign n35557 = n22408 & n31243;
  assign n35558 = n22405 & n22408;
  assign n35559 = (n35432 & n35557) | (n35432 & n35558) | (n35557 & n35558);
  assign n22410 = n35556 & ~n35559;
  assign n22411 = n22153 & n22410;
  assign n31246 = n22159 | n22411;
  assign n31296 = n22471 | n31246;
  assign n31245 = n22411 | n31237;
  assign n31297 = n22471 | n31245;
  assign n31298 = (n31069 & n31296) | (n31069 & n31297) | (n31296 & n31297);
  assign n31299 = n22471 & n31246;
  assign n31300 = n22471 & n31245;
  assign n31301 = (n31069 & n31299) | (n31069 & n31300) | (n31299 & n31300);
  assign n22474 = n31298 & ~n31301;
  assign n22475 = x132 & x152;
  assign n22476 = n22474 | n22475;
  assign n22477 = n22474 & n22475;
  assign n22478 = n22476 & ~n22477;
  assign n31302 = ~n22401 & n22478;
  assign n31303 = ~n31236 & n31302;
  assign n31304 = n22401 & ~n22478;
  assign n31305 = (~n22478 & n31236) | (~n22478 & n31304) | (n31236 & n31304);
  assign n22481 = n31303 | n31305;
  assign n22482 = x131 & x153;
  assign n22483 = n22481 & n22482;
  assign n22484 = n22481 | n22482;
  assign n22485 = ~n22483 & n22484;
  assign n31306 = n22396 | n22485;
  assign n31307 = n31226 | n31306;
  assign n31308 = n22396 & n22485;
  assign n31309 = (n22485 & n31226) | (n22485 & n31308) | (n31226 & n31308);
  assign n22488 = n31307 & ~n31309;
  assign n22489 = x130 & x154;
  assign n22490 = n22488 | n22489;
  assign n22491 = n22488 & n22489;
  assign n22492 = n22490 & ~n22491;
  assign n31310 = ~n22388 & n22492;
  assign n31311 = ~n31217 & n31310;
  assign n31312 = n22388 & ~n22492;
  assign n31313 = (~n22492 & n31217) | (~n22492 & n31312) | (n31217 & n31312);
  assign n22495 = n31311 | n31313;
  assign n22496 = x129 & x155;
  assign n22497 = n22495 & n22496;
  assign n22498 = n22495 | n22496;
  assign n22499 = ~n22497 & n22498;
  assign n22500 = ~n31223 & n22499;
  assign n22501 = n31223 & ~n22499;
  assign n22502 = n22500 | n22501;
  assign n22503 = x128 & x156;
  assign n22504 = n22502 | n22503;
  assign n22505 = n22502 & n22503;
  assign n22506 = n22504 & ~n22505;
  assign n22507 = ~n31215 & n22506;
  assign n22508 = n31215 & ~n22506;
  assign n22509 = n22507 | n22508;
  assign n22510 = x127 & x157;
  assign n22511 = n22509 & n22510;
  assign n22512 = n22509 | n22510;
  assign n22513 = ~n22511 & n22512;
  assign n22514 = n31207 | n22513;
  assign n22515 = n31207 & n22513;
  assign n22516 = n22514 & ~n22515;
  assign n22517 = x126 & x158;
  assign n22518 = n22516 | n22517;
  assign n22519 = n22516 & n22517;
  assign n22520 = n22518 & ~n22519;
  assign n22521 = ~n31198 & n22520;
  assign n22522 = n31198 & ~n22520;
  assign n22523 = n22521 | n22522;
  assign n22524 = x125 & x159;
  assign n22525 = n22523 & n22524;
  assign n22526 = n22523 | n22524;
  assign n22527 = ~n22525 & n22526;
  assign n22528 = n22357 | n22527;
  assign n22529 = n22357 & n22527;
  assign n22530 = n22528 & ~n22529;
  assign n22531 = x124 & x160;
  assign n22532 = n22530 | n22531;
  assign n22533 = n22530 & n22531;
  assign n22534 = n22532 & ~n22533;
  assign n22535 = n31192 | n22534;
  assign n22536 = n31192 & n22534;
  assign n22537 = n22535 & ~n22536;
  assign n22538 = x123 & x161;
  assign n22539 = n22537 | n22538;
  assign n22540 = n22537 & n22538;
  assign n22541 = n22539 & ~n22540;
  assign n22542 = n31037 | n22345;
  assign n31314 = n22227 & ~n22345;
  assign n31315 = (n22227 & ~n31037) | (n22227 & n31314) | (~n31037 & n31314);
  assign n22544 = n22542 & n31315;
  assign n31316 = n22236 | n22544;
  assign n31317 = (n22544 & n31153) | (n22544 & n31316) | (n31153 & n31316);
  assign n22546 = n22541 | n31317;
  assign n22547 = n22541 & n31317;
  assign n22548 = n22546 & ~n22547;
  assign n22549 = x122 & x162;
  assign n22550 = n22548 | n22549;
  assign n22551 = n22548 & n22549;
  assign n22552 = n22550 & ~n22551;
  assign n22553 = n31190 | n22552;
  assign n22554 = n31190 & n22552;
  assign n22555 = n22553 & ~n22554;
  assign n22556 = x121 & x163;
  assign n22557 = ~n22555 & n22556;
  assign n22558 = n22555 & ~n22556;
  assign n22559 = n22557 | n22558;
  assign n31318 = n22254 & n22262;
  assign n31319 = (n22254 & n31156) | (n22254 & n31318) | (n31156 & n31318);
  assign n31320 = n22029 | n22247;
  assign n31321 = n31031 | n31320;
  assign n35560 = ~n22029 & n22248;
  assign n35561 = (~n22247 & n22248) | (~n22247 & n35560) | (n22248 & n35560);
  assign n31323 = ~n22247 & n22248;
  assign n31324 = (~n31031 & n35561) | (~n31031 & n31323) | (n35561 & n31323);
  assign n22563 = n31321 & n31324;
  assign n22564 = n31319 | n22563;
  assign n22565 = n22559 & n22564;
  assign n22566 = n22559 | n22564;
  assign n22567 = ~n22565 & n22566;
  assign n22568 = x120 & x164;
  assign n22569 = ~n22567 & n22568;
  assign n22570 = n22567 & ~n22568;
  assign n22571 = n22569 | n22570;
  assign n31325 = n22254 | n22262;
  assign n31326 = n31156 | n31325;
  assign n22573 = n22255 & ~n31319;
  assign n22574 = n31326 & n22573;
  assign n22575 = n31181 | n22574;
  assign n22576 = n22571 & n22575;
  assign n22577 = n22571 | n22575;
  assign n22578 = ~n22576 & n22577;
  assign n31327 = ~n22335 & n22578;
  assign n31328 = ~n31178 & n31327;
  assign n31329 = n22335 & ~n22578;
  assign n31330 = (~n22578 & n31178) | (~n22578 & n31329) | (n31178 & n31329);
  assign n22581 = n31328 | n31330;
  assign n22582 = x119 & x165;
  assign n22583 = n22581 & n22582;
  assign n22584 = n22581 | n22582;
  assign n22585 = ~n22583 & n22584;
  assign n31331 = n22282 & n22585;
  assign n31332 = (n22585 & n31170) | (n22585 & n31331) | (n31170 & n31331);
  assign n31333 = n22282 | n22585;
  assign n31334 = n31170 | n31333;
  assign n22588 = ~n31332 & n31334;
  assign n22589 = n22329 | n22588;
  assign n22590 = n22329 & n22588;
  assign n22591 = n22589 & ~n22590;
  assign n31335 = n22288 & n22289;
  assign n31336 = (n22288 & n31174) | (n22288 & n31335) | (n31174 & n31335);
  assign n22594 = n22591 & ~n31336;
  assign n22595 = ~n22591 & n31336;
  assign n22596 = n22594 | n22595;
  assign n22597 = x117 & x167;
  assign n22598 = n22596 | n22597;
  assign n22599 = n22596 & n22597;
  assign n22600 = n22598 & ~n22599;
  assign n31337 = n22297 & n22298;
  assign n31338 = (n22297 & n31176) | (n22297 & n31337) | (n31176 & n31337);
  assign n22603 = n22600 & ~n31338;
  assign n22604 = ~n22600 & n31338;
  assign n22605 = n22603 | n22604;
  assign n22606 = x116 & x168;
  assign n22607 = n22605 | n22606;
  assign n22608 = n22605 & n22606;
  assign n22609 = n22607 & ~n22608;
  assign n31339 = n22306 & n22307;
  assign n31340 = (n22306 & n31024) | (n22306 & n31339) | (n31024 & n31339);
  assign n22612 = n22609 & ~n31340;
  assign n22613 = ~n22609 & n31340;
  assign n22614 = n22612 | n22613;
  assign n22615 = x115 & x169;
  assign n22616 = n22614 | n22615;
  assign n22617 = n22614 & n22615;
  assign n22618 = n22616 & ~n22617;
  assign n22619 = n22010 | n22312;
  assign n22620 = n22313 & n22619;
  assign n22621 = n22618 & ~n22620;
  assign n22622 = ~n22618 & n22620;
  assign n22623 = n22621 | n22622;
  assign n22624 = x114 & x170;
  assign n22625 = n22623 | n22624;
  assign n22626 = n22623 & n22624;
  assign n22627 = n22625 & ~n22626;
  assign n22628 = n22003 | n22319;
  assign n22629 = n22318 & n22628;
  assign n22630 = n22627 & ~n22629;
  assign n22631 = ~n22627 & n22629;
  assign n22632 = n22630 | n22631;
  assign n22633 = n22328 & ~n22632;
  assign n22634 = ~n22328 & n22632;
  assign n22635 = n22633 | n22634;
  assign n22636 = ~n22325 & n22635;
  assign n22637 = n22325 & ~n22635;
  assign n22638 = n22636 | n22637;
  assign n22639 = x112 & x172;
  assign n22640 = n22638 & n22639;
  assign n22641 = n22638 | n22639;
  assign n22642 = ~n22640 & n22641;
  assign n31341 = n22625 & n22626;
  assign n31342 = (n22625 & n22629) | (n22625 & n31341) | (n22629 & n31341);
  assign n22645 = x114 & x171;
  assign n22646 = n31342 & n22645;
  assign n22647 = n31342 | n22645;
  assign n22648 = ~n22646 & n22647;
  assign n22649 = x115 & x170;
  assign n31343 = n22616 & n22617;
  assign n31344 = (n22616 & n22620) | (n22616 & n31343) | (n22620 & n31343);
  assign n22652 = x116 & x169;
  assign n31345 = n22607 & n22608;
  assign n31346 = (n22607 & n31340) | (n22607 & n31345) | (n31340 & n31345);
  assign n22655 = x119 & x166;
  assign n31347 = n22335 & n22578;
  assign n31348 = (n22578 & n31178) | (n22578 & n31347) | (n31178 & n31347);
  assign n31349 = n22567 & n22574;
  assign n31350 = (n22567 & n31181) | (n22567 & n31349) | (n31181 & n31349);
  assign n31351 = n22567 | n22574;
  assign n31352 = n31181 | n31351;
  assign n22660 = n22568 & n31352;
  assign n22661 = ~n31350 & n22660;
  assign n31353 = n22537 & n31316;
  assign n31354 = n22537 & n22544;
  assign n31355 = (n31153 & n31353) | (n31153 & n31354) | (n31353 & n31354);
  assign n31356 = n22537 | n31316;
  assign n31357 = n22537 | n22544;
  assign n31358 = (n31153 & n31356) | (n31153 & n31357) | (n31356 & n31357);
  assign n22666 = n22538 & n31358;
  assign n22667 = ~n31355 & n22666;
  assign n31359 = n22548 | n22667;
  assign n31360 = (n22667 & n31190) | (n22667 & n31359) | (n31190 & n31359);
  assign n22669 = n31192 | n22530;
  assign n22670 = n31037 | n22343;
  assign n37426 = ~n22226 & n22531;
  assign n37427 = ~n22225 & n37426;
  assign n35563 = (~n22530 & n22531) | (~n22530 & n37427) | (n22531 & n37427);
  assign n31362 = (n22531 & ~n22670) | (n22531 & n35563) | (~n22670 & n35563);
  assign n22674 = n22669 & n31362;
  assign n22675 = n31355 | n22674;
  assign n22676 = n22356 | n22523;
  assign n22677 = n31149 | n22676;
  assign n22678 = n22039 | n22356;
  assign n22679 = n30998 | n22678;
  assign n22354 = n22351 & n22353;
  assign n22680 = n22349 & ~n22354;
  assign n22681 = n22052 | n22680;
  assign n22682 = n22523 & n22681;
  assign n22683 = n22679 & n22682;
  assign n22684 = n22677 & ~n22683;
  assign n22685 = n22524 & n22684;
  assign n22671 = n22344 & n22530;
  assign n31363 = n22671 | n22685;
  assign n31364 = (n22670 & n22685) | (n22670 & n31363) | (n22685 & n31363);
  assign n22689 = n31049 | n31205;
  assign n31368 = n22203 | n31201;
  assign n31369 = (n22203 & ~n22367) | (n22203 & n31368) | (~n22367 & n31368);
  assign n22691 = n22509 & n31369;
  assign n22692 = n22689 & n22691;
  assign n31365 = n22509 | n31206;
  assign n31366 = n22509 | n31205;
  assign n31367 = (n31049 & n31365) | (n31049 & n31366) | (n31365 & n31366);
  assign n31370 = n22510 & n31367;
  assign n31371 = ~n22692 & n31370;
  assign n31372 = n22516 | n31371;
  assign n31373 = (n31198 & n31371) | (n31198 & n31372) | (n31371 & n31372);
  assign n22697 = n22383 | n22495;
  assign n31374 = n22697 | n31208;
  assign n31375 = n22191 | n22697;
  assign n31376 = (n31051 & n31374) | (n31051 & n31375) | (n31374 & n31375);
  assign n22700 = n22185 | n22382;
  assign n22701 = n22495 & n22700;
  assign n31377 = n22198 | n22383;
  assign n31379 = n22701 & n31377;
  assign n31380 = (n22701 & n31051) | (n22701 & n31379) | (n31051 & n31379);
  assign n22703 = n31376 & ~n31380;
  assign n22704 = n22496 & n22703;
  assign n31381 = n22502 | n22704;
  assign n35564 = (n22704 & n31381) | (n22704 & n35513) | (n31381 & n35513);
  assign n35565 = (n22374 & n22704) | (n22374 & n31381) | (n22704 & n31381);
  assign n35566 = (n22364 & n35564) | (n22364 & n35565) | (n35564 & n35565);
  assign n31385 = n22396 | n31139;
  assign n31386 = n22180 | n22396;
  assign n31387 = (n31060 & n31385) | (n31060 & n31386) | (n31385 & n31386);
  assign n22720 = x132 & x153;
  assign n22723 = n22153 | n22410;
  assign n22724 = n22467 & n22723;
  assign n22721 = n22093 | n22411;
  assign n31401 = n22721 & n22724;
  assign n35569 = (n22724 & n31068) | (n22724 & n31401) | (n31068 & n31401);
  assign n35570 = (n22084 & n22724) | (n22084 & n31401) | (n22724 & n31401);
  assign n35571 = (n30779 & n35569) | (n30779 & n35570) | (n35569 & n35570);
  assign n31410 = n22416 & n22460;
  assign n35577 = (n22408 & n22460) | (n22408 & n31410) | (n22460 & n31410);
  assign n35578 = (n31243 & n31410) | (n31243 & n35577) | (n31410 & n35577);
  assign n35579 = (n22405 & n31410) | (n22405 & n35577) | (n31410 & n35577);
  assign n35580 = (n35432 & n35578) | (n35432 & n35579) | (n35578 & n35579);
  assign n31413 = n22416 | n22460;
  assign n35581 = n22408 | n31413;
  assign n35582 = (n31243 & n31413) | (n31243 & n35581) | (n31413 & n35581);
  assign n35583 = (n22405 & n31413) | (n22405 & n35581) | (n31413 & n35581);
  assign n35584 = (n35432 & n35582) | (n35432 & n35583) | (n35582 & n35583);
  assign n22732 = n22461 & n35584;
  assign n22733 = ~n35580 & n22732;
  assign n22750 = x141 & x144;
  assign n22751 = x140 & x145;
  assign n22752 = n22750 & n22751;
  assign n22753 = n22750 | n22751;
  assign n22754 = ~n22752 & n22753;
  assign n22755 = x139 & x146;
  assign n22756 = n22754 & n22755;
  assign n22757 = n22754 | n22755;
  assign n22758 = ~n22756 & n22757;
  assign n22745 = n21813 | n22427;
  assign n22746 = n21812 & n22745;
  assign n31424 = n21817 | n22746;
  assign n37428 = n22109 | n22429;
  assign n37429 = (n22429 & n22430) | (n22429 & n37428) | (n22430 & n37428);
  assign n35586 = (n22429 & n31424) | (n22429 & n37429) | (n31424 & n37429);
  assign n31432 = n22758 & ~n35586;
  assign n35587 = n22429 | n22746;
  assign n35588 = (n22429 & n22431) | (n22429 & n35587) | (n22431 & n35587);
  assign n31433 = n22758 & ~n35588;
  assign n31434 = (~n35438 & n31432) | (~n35438 & n31433) | (n31432 & n31433);
  assign n31435 = ~n22758 & n35586;
  assign n31436 = ~n22758 & n35588;
  assign n31437 = (n35438 & n31435) | (n35438 & n31436) | (n31435 & n31436);
  assign n22761 = n31434 | n31437;
  assign n31439 = n22437 | n22761;
  assign n35532 = (n22423 & n31099) | (n22423 & n37417) | (n31099 & n37417);
  assign n35589 = n22439 | n31439;
  assign n35590 = (n31439 & n35532) | (n31439 & n35589) | (n35532 & n35589);
  assign n35531 = (n22423 & n31098) | (n22423 & n37417) | (n31098 & n37417);
  assign n35591 = (n31439 & n35531) | (n31439 & n35589) | (n35531 & n35589);
  assign n35592 = (n35269 & n35590) | (n35269 & n35591) | (n35590 & n35591);
  assign n22764 = n22438 & n22761;
  assign n31441 = n22437 & n22764;
  assign n35593 = (n22764 & n31441) | (n22764 & n35532) | (n31441 & n35532);
  assign n35594 = (n22764 & n31441) | (n22764 & n35531) | (n31441 & n35531);
  assign n35595 = (n35269 & n35593) | (n35269 & n35594) | (n35593 & n35594);
  assign n22766 = n35592 & ~n35595;
  assign n22767 = x138 & x147;
  assign n22768 = n22766 & n22767;
  assign n22769 = n22766 | n22767;
  assign n22770 = ~n22768 & n22769;
  assign n31443 = n22444 | n22770;
  assign n31444 = n35545 | n31443;
  assign n31446 = n22444 | n35542;
  assign n35596 = n22444 | n31105;
  assign n35597 = n31116 | n35596;
  assign n35598 = (n30831 & n31446) | (n30831 & n35597) | (n31446 & n35597);
  assign n35599 = (n31446 & n35400) | (n31446 & n35597) | (n35400 & n35597);
  assign n35600 = (n30333 & n35598) | (n30333 & n35599) | (n35598 & n35599);
  assign n22774 = n22761 & ~n22767;
  assign n22775 = ~n22761 & n22767;
  assign n22776 = n22774 | n22775;
  assign n31422 = n22437 | n22439;
  assign n31448 = n22776 | n31422;
  assign n31449 = n22437 | n22776;
  assign n35601 = (n31448 & n31449) | (n31448 & n35532) | (n31449 & n35532);
  assign n35602 = (n31448 & n31449) | (n31448 & n35531) | (n31449 & n35531);
  assign n35603 = (n35269 & n35601) | (n35269 & n35602) | (n35601 & n35602);
  assign n31451 = n22776 & n31422;
  assign n31452 = n22437 & n22776;
  assign n35604 = (n31451 & n31452) | (n31451 & n35532) | (n31452 & n35532);
  assign n35605 = (n31451 & n31452) | (n31451 & n35531) | (n31452 & n35531);
  assign n35606 = (n35269 & n35604) | (n35269 & n35605) | (n35604 & n35605);
  assign n31454 = n22443 & ~n35606;
  assign n31455 = (n22442 & ~n35606) | (n22442 & n31454) | (~n35606 & n31454);
  assign n22780 = n35603 & n31455;
  assign n22781 = n35600 & n22780;
  assign n22782 = n31444 & ~n22781;
  assign n22783 = x137 & x148;
  assign n22784 = n22782 & n22783;
  assign n22785 = n22782 | n22783;
  assign n22786 = ~n22784 & n22785;
  assign n22787 = x136 & x149;
  assign n22788 = n22786 & n22787;
  assign n22789 = n22786 | n22787;
  assign n22790 = ~n22788 & n22789;
  assign n22739 = n22143 & n22453;
  assign n22737 = n21837 | n22142;
  assign n31415 = n22099 | n22737;
  assign n31417 = n22739 & n31415;
  assign n31418 = n22737 & n22739;
  assign n31419 = (n31086 & n31417) | (n31086 & n31418) | (n31417 & n31418);
  assign n31456 = n22451 & ~n22790;
  assign n31457 = (~n22790 & n31419) | (~n22790 & n31456) | (n31419 & n31456);
  assign n31458 = ~n22451 & n22790;
  assign n31459 = ~n31419 & n31458;
  assign n22794 = n31457 | n31459;
  assign n22795 = x135 & x150;
  assign n22796 = n22794 & n22795;
  assign n22797 = n22794 | n22795;
  assign n22798 = ~n22796 & n22797;
  assign n22735 = n22142 | n22453;
  assign n22736 = n35526 | n22735;
  assign n37851 = ~n22141 & n22454;
  assign n37852 = ~n22140 & n37851;
  assign n37746 = (~n22453 & n22454) | (~n22453 & n37852) | (n22454 & n37852);
  assign n37431 = (n22454 & ~n31415) | (n22454 & n37746) | (~n31415 & n37746);
  assign n37432 = n22454 & ~n22737;
  assign n37433 = (n22454 & ~n22739) | (n22454 & n37432) | (~n22739 & n37432);
  assign n35609 = (~n31086 & n37431) | (~n31086 & n37433) | (n37431 & n37433);
  assign n31421 = n22736 & n35609;
  assign n31460 = n22798 | n31421;
  assign n31461 = n35580 | n31460;
  assign n31462 = n22798 & n31421;
  assign n31463 = (n22798 & n35580) | (n22798 & n31462) | (n35580 & n31462);
  assign n22801 = n31461 & ~n31463;
  assign n22802 = x134 & x151;
  assign n22803 = n22801 | n22802;
  assign n22804 = n22801 & n22802;
  assign n22805 = n22803 & ~n22804;
  assign n31464 = ~n22733 & n22805;
  assign n31465 = ~n35571 & n31464;
  assign n31466 = n22733 & ~n22805;
  assign n31467 = (~n22805 & n35571) | (~n22805 & n31466) | (n35571 & n31466);
  assign n22808 = n31465 | n31467;
  assign n22809 = x133 & x152;
  assign n22810 = n22808 & n22809;
  assign n22811 = n22808 | n22809;
  assign n22812 = ~n22810 & n22811;
  assign n31403 = n22467 | n31246;
  assign n35572 = n22411 | n22467;
  assign n35573 = n31237 | n35572;
  assign n35574 = (n31068 & n31403) | (n31068 & n35573) | (n31403 & n35573);
  assign n35575 = (n22084 & n31403) | (n22084 & n35573) | (n31403 & n35573);
  assign n35576 = (n30779 & n35574) | (n30779 & n35575) | (n35574 & n35575);
  assign n22727 = ~n35571 & n35576;
  assign n22728 = n22468 & n22727;
  assign n31393 = n22401 & n22474;
  assign n31406 = n22728 | n31393;
  assign n35610 = n22812 | n31406;
  assign n31407 = n22474 | n22728;
  assign n35611 = n22812 | n31407;
  assign n35612 = (n31236 & n35610) | (n31236 & n35611) | (n35610 & n35611);
  assign n35613 = n22812 & n31406;
  assign n35614 = n22812 & n31407;
  assign n35615 = (n31236 & n35613) | (n31236 & n35614) | (n35613 & n35614);
  assign n22815 = n35612 & ~n35615;
  assign n22816 = n22720 & n22815;
  assign n22817 = n22720 | n22815;
  assign n22818 = ~n22816 & n22817;
  assign n22708 = n22167 | n22395;
  assign n22709 = n22481 & n22708;
  assign n31394 = (n22474 & n31236) | (n22474 & n31393) | (n31236 & n31393);
  assign n35567 = n22401 & n22475;
  assign n35568 = (n22474 & n22475) | (n22474 & n35567) | (n22475 & n35567);
  assign n31398 = (n22475 & n31236) | (n22475 & n35568) | (n31236 & n35568);
  assign n22718 = ~n31394 & n31398;
  assign n31399 = n22709 | n22718;
  assign n35616 = n22818 & ~n31399;
  assign n35617 = ~n22718 & n22818;
  assign n35618 = (~n31387 & n35616) | (~n31387 & n35617) | (n35616 & n35617);
  assign n35619 = ~n22818 & n31399;
  assign n35620 = n22718 & ~n22818;
  assign n35621 = (n31387 & n35619) | (n31387 & n35620) | (n35619 & n35620);
  assign n22821 = n35618 | n35621;
  assign n22822 = x131 & x154;
  assign n22823 = n22821 & n22822;
  assign n22824 = n22821 | n22822;
  assign n22825 = ~n22823 & n22824;
  assign n22710 = n31387 & n22709;
  assign n31388 = n22396 | n22481;
  assign n31389 = n31226 | n31388;
  assign n22712 = ~n22710 & n31389;
  assign n22713 = n22482 & n22712;
  assign n31391 = n22488 | n22713;
  assign n35622 = n22825 | n31391;
  assign n31383 = n22388 & n22488;
  assign n31390 = n22713 | n31383;
  assign n35623 = n22825 | n31390;
  assign n35624 = (n31217 & n35622) | (n31217 & n35623) | (n35622 & n35623);
  assign n35625 = n22825 & n31391;
  assign n35626 = n22825 & n31390;
  assign n35627 = (n31217 & n35625) | (n31217 & n35626) | (n35625 & n35626);
  assign n22828 = n35624 & ~n35627;
  assign n22829 = x130 & x155;
  assign n22830 = n22828 | n22829;
  assign n22831 = n22828 & n22829;
  assign n22832 = n22830 & ~n22831;
  assign n31468 = n22388 | n22488;
  assign n31469 = n31217 | n31468;
  assign n31470 = n22489 & ~n31383;
  assign n31471 = ~n22488 & n22489;
  assign n31472 = (~n31217 & n31470) | (~n31217 & n31471) | (n31470 & n31471);
  assign n22835 = n31469 & n31472;
  assign n35628 = ~n22832 & n22835;
  assign n35629 = (~n22832 & n31380) | (~n22832 & n35628) | (n31380 & n35628);
  assign n35630 = n22832 & ~n22835;
  assign n35631 = ~n31380 & n35630;
  assign n22839 = n35629 | n35631;
  assign n22840 = x129 & x156;
  assign n22841 = n22839 & n22840;
  assign n22842 = n22839 | n22840;
  assign n22843 = ~n22841 & n22842;
  assign n22844 = n35566 | n22843;
  assign n22845 = n35566 & n22843;
  assign n22846 = n22844 & ~n22845;
  assign n22847 = x128 & x157;
  assign n22848 = ~n22846 & n22847;
  assign n22849 = n22846 & ~n22847;
  assign n22850 = n22848 | n22849;
  assign n35632 = n22502 | n35513;
  assign n35633 = n22374 | n22502;
  assign n35634 = (n22364 & n35632) | (n22364 & n35633) | (n35632 & n35633);
  assign n31473 = ~n22502 & n22503;
  assign n35635 = (n22503 & n31473) | (n22503 & ~n35513) | (n31473 & ~n35513);
  assign n37434 = ~n22374 & n22503;
  assign n37435 = (~n22502 & n22503) | (~n22502 & n37434) | (n22503 & n37434);
  assign n35637 = (~n22364 & n35635) | (~n22364 & n37435) | (n35635 & n37435);
  assign n22853 = n35634 & n35637;
  assign n35638 = n22853 | n31369;
  assign n35639 = (n22509 & n22853) | (n22509 & n35638) | (n22853 & n35638);
  assign n31476 = (n22689 & n22853) | (n22689 & n35639) | (n22853 & n35639);
  assign n22855 = n22850 & ~n31476;
  assign n22856 = ~n22850 & n31476;
  assign n22857 = n22855 | n22856;
  assign n22858 = x127 & x158;
  assign n22859 = n22857 & n22858;
  assign n22860 = n22857 | n22858;
  assign n22861 = ~n22859 & n22860;
  assign n22862 = n31373 | n22861;
  assign n22863 = n31373 & n22861;
  assign n22864 = n22862 & ~n22863;
  assign n22865 = x126 & x159;
  assign n22866 = n22864 | n22865;
  assign n22867 = n22864 & n22865;
  assign n22868 = n22866 & ~n22867;
  assign n22869 = n31198 | n22516;
  assign n31477 = ~n22516 & n22517;
  assign n31478 = (n22517 & ~n31198) | (n22517 & n31477) | (~n31198 & n31477);
  assign n22871 = n22869 & n31478;
  assign n31479 = n22682 | n22871;
  assign n31480 = (n22679 & n22871) | (n22679 & n31479) | (n22871 & n31479);
  assign n22873 = ~n22868 & n31480;
  assign n22874 = n22868 & ~n31480;
  assign n22875 = n22873 | n22874;
  assign n22876 = x125 & x160;
  assign n22877 = n22875 & n22876;
  assign n22878 = n22875 | n22876;
  assign n22879 = ~n22877 & n22878;
  assign n22880 = n31364 | n22879;
  assign n22881 = n31364 & n22879;
  assign n22882 = n22880 & ~n22881;
  assign n22883 = x124 & x161;
  assign n22884 = n22882 | n22883;
  assign n22885 = n22882 & n22883;
  assign n22886 = n22884 & ~n22885;
  assign n22887 = n22675 | n22886;
  assign n22888 = n22675 & n22886;
  assign n22889 = n22887 & ~n22888;
  assign n22890 = x123 & x162;
  assign n22891 = n22889 | n22890;
  assign n22892 = n22889 & n22890;
  assign n22893 = n22891 & ~n22892;
  assign n22894 = n31360 | n22893;
  assign n22895 = n31360 & n22893;
  assign n22896 = n22894 & ~n22895;
  assign n22897 = x122 & x163;
  assign n22898 = ~n22896 & n22897;
  assign n22899 = n22896 & ~n22897;
  assign n22900 = n22898 | n22899;
  assign n22902 = n31190 | n22548;
  assign n31483 = ~n22548 & n22549;
  assign n31484 = (n22549 & ~n31190) | (n22549 & n31483) | (~n31190 & n31483);
  assign n22904 = n22902 & n31484;
  assign n31481 = n22555 & n22563;
  assign n31485 = n22904 | n31481;
  assign n31486 = n22555 | n22904;
  assign n31487 = (n31319 & n31485) | (n31319 & n31486) | (n31485 & n31486);
  assign n22906 = n22900 & n31487;
  assign n22907 = n22900 | n31487;
  assign n22908 = ~n22906 & n22907;
  assign n22909 = x121 & x164;
  assign n22910 = ~n22908 & n22909;
  assign n22911 = n22908 & ~n22909;
  assign n22912 = n22910 | n22911;
  assign n31488 = n22555 | n22563;
  assign n31489 = n31319 | n31488;
  assign n35640 = n22556 & ~n22563;
  assign n35641 = (~n22555 & n22556) | (~n22555 & n35640) | (n22556 & n35640);
  assign n31491 = (n22557 & ~n31319) | (n22557 & n35641) | (~n31319 & n35641);
  assign n22915 = n31489 & n31491;
  assign n22916 = n31350 | n22915;
  assign n22917 = n22912 & n22916;
  assign n22918 = n22912 | n22916;
  assign n22919 = ~n22917 & n22918;
  assign n31492 = ~n22661 & n22919;
  assign n31493 = ~n31348 & n31492;
  assign n31494 = n22661 & ~n22919;
  assign n31495 = (~n22919 & n31348) | (~n22919 & n31494) | (n31348 & n31494);
  assign n22922 = n31493 | n31495;
  assign n22923 = x120 & x165;
  assign n22924 = n22922 & n22923;
  assign n22925 = n22922 | n22923;
  assign n22926 = ~n22924 & n22925;
  assign n31496 = n22583 & n22926;
  assign n31497 = (n22926 & n31332) | (n22926 & n31496) | (n31332 & n31496);
  assign n31498 = n22583 | n22926;
  assign n31499 = n31332 | n31498;
  assign n22929 = ~n31497 & n31499;
  assign n22930 = n22655 | n22929;
  assign n22931 = n22655 & n22929;
  assign n22932 = n22930 & ~n22931;
  assign n31500 = n22589 & n22590;
  assign n31501 = (n22589 & n31336) | (n22589 & n31500) | (n31336 & n31500);
  assign n22935 = n22932 & ~n31501;
  assign n22936 = ~n22932 & n31501;
  assign n22937 = n22935 | n22936;
  assign n22938 = x118 & x167;
  assign n22939 = n22937 | n22938;
  assign n22940 = n22937 & n22938;
  assign n22941 = n22939 & ~n22940;
  assign n31502 = n22598 & n22599;
  assign n31503 = (n22598 & n31338) | (n22598 & n31502) | (n31338 & n31502);
  assign n22944 = n22941 & ~n31503;
  assign n22945 = ~n22941 & n31503;
  assign n22946 = n22944 | n22945;
  assign n22947 = x117 & x168;
  assign n22948 = n22946 | n22947;
  assign n22949 = n22946 & n22947;
  assign n22950 = n22948 & ~n22949;
  assign n22951 = ~n31346 & n22950;
  assign n22952 = n31346 & ~n22950;
  assign n22953 = n22951 | n22952;
  assign n22954 = n22652 & n22953;
  assign n22955 = n22652 | n22953;
  assign n22956 = ~n22954 & n22955;
  assign n22957 = n31344 & n22956;
  assign n22958 = n31344 | n22956;
  assign n22959 = ~n22957 & n22958;
  assign n22960 = n22649 | n22959;
  assign n22961 = n22649 & n22959;
  assign n22962 = n22960 & ~n22961;
  assign n22963 = ~n22648 & n22962;
  assign n22964 = n22648 & ~n22962;
  assign n22965 = n22963 | n22964;
  assign n31504 = n22324 & n22328;
  assign n31505 = n22323 & n31504;
  assign n22967 = n22632 | n31505;
  assign n31506 = n22324 | n22328;
  assign n31507 = (n22323 & n22328) | (n22323 & n31506) | (n22328 & n31506);
  assign n22969 = n22967 & n31507;
  assign n22970 = n22965 & ~n22969;
  assign n22971 = ~n22965 & n22969;
  assign n22972 = n22970 | n22971;
  assign n22973 = x113 & x172;
  assign n22974 = n22972 | n22973;
  assign n22975 = n22972 & n22973;
  assign n22976 = n22974 & ~n22975;
  assign n22977 = ~n22640 & n22976;
  assign n22978 = n22640 & ~n22976;
  assign n22979 = n22977 | n22978;
  assign n22980 = x112 & x173;
  assign n22981 = n22979 & n22980;
  assign n22982 = n22979 | n22980;
  assign n22983 = ~n22981 & n22982;
  assign n31508 = n22948 & n22949;
  assign n31509 = (n22948 & n31346) | (n22948 & n31508) | (n31346 & n31508);
  assign n22986 = x117 & x169;
  assign n22987 = n31509 & n22986;
  assign n22988 = n31509 | n22986;
  assign n22989 = ~n22987 & n22988;
  assign n22990 = x120 & x166;
  assign n31510 = n22661 & n22919;
  assign n31511 = (n22919 & n31348) | (n22919 & n31510) | (n31348 & n31510);
  assign n31512 = n22908 & n22915;
  assign n31513 = (n22908 & n31350) | (n22908 & n31512) | (n31350 & n31512);
  assign n35642 = n22909 & n22915;
  assign n35643 = (n22908 & n22909) | (n22908 & n35642) | (n22909 & n35642);
  assign n31517 = (n22909 & n31350) | (n22909 & n35643) | (n31350 & n35643);
  assign n22996 = ~n31513 & n31517;
  assign n31518 = n22889 & n31359;
  assign n31519 = n22667 & n22889;
  assign n31520 = (n31190 & n31518) | (n31190 & n31519) | (n31518 & n31519);
  assign n31521 = n22674 & n22882;
  assign n31522 = (n22882 & n31355) | (n22882 & n31521) | (n31355 & n31521);
  assign n31523 = n22674 | n22882;
  assign n31524 = n31355 | n31523;
  assign n23001 = n22883 & n31524;
  assign n23002 = ~n31522 & n23001;
  assign n23003 = n31520 | n23002;
  assign n23004 = x125 & x161;
  assign n22346 = n31037 & n22345;
  assign n23007 = n22524 | n22684;
  assign n23008 = n22875 & n23007;
  assign n23005 = n22343 | n22685;
  assign n31525 = n23005 & n23008;
  assign n31526 = (n22346 & n23008) | (n22346 & n31525) | (n23008 & n31525);
  assign n23010 = n22864 & n31480;
  assign n31527 = (n22865 & n22867) | (n22865 & n31480) | (n22867 & n31480);
  assign n23013 = ~n23010 & n31527;
  assign n23014 = n31526 | n23013;
  assign n23016 = n31198 | n31371;
  assign n31531 = n22510 | n31367;
  assign n31532 = (n22510 & ~n22692) | (n22510 & n31531) | (~n22692 & n31531);
  assign n23018 = n22857 & n31532;
  assign n23019 = n23016 & n23018;
  assign n31528 = n22857 | n31372;
  assign n31529 = n22857 | n31371;
  assign n31530 = (n31198 & n31528) | (n31198 & n31529) | (n31528 & n31529);
  assign n31533 = n22858 & n31530;
  assign n31534 = ~n23019 & n31533;
  assign n31535 = n22864 | n31534;
  assign n31536 = (n31480 & n31534) | (n31480 & n31535) | (n31534 & n31535);
  assign n35644 = n22846 & n35639;
  assign n35645 = n22846 & n22853;
  assign n35646 = (n22689 & n35644) | (n22689 & n35645) | (n35644 & n35645);
  assign n31537 = n22846 & n22847;
  assign n35647 = (n22847 & n31537) | (n22847 & n35639) | (n31537 & n35639);
  assign n37436 = n22847 & n22853;
  assign n37437 = (n22846 & n22847) | (n22846 & n37436) | (n22847 & n37436);
  assign n35649 = (n22689 & n35647) | (n22689 & n37437) | (n35647 & n37437);
  assign n23026 = ~n35646 & n35649;
  assign n35650 = n23026 | n31532;
  assign n35651 = (n22857 & n23026) | (n22857 & n35650) | (n23026 & n35650);
  assign n31540 = (n23016 & n23026) | (n23016 & n35651) | (n23026 & n35651);
  assign n23028 = n22374 | n22704;
  assign n31541 = n22366 | n23028;
  assign n31542 = (n22364 & n23028) | (n22364 & n31541) | (n23028 & n31541);
  assign n23030 = n22496 | n22703;
  assign n23031 = n22839 & n23030;
  assign n23032 = n31542 & n23031;
  assign n31543 = n22839 | n31381;
  assign n31544 = n22704 | n22839;
  assign n31545 = (n31215 & n31543) | (n31215 & n31544) | (n31543 & n31544);
  assign n23034 = ~n23032 & n31545;
  assign n23035 = n22840 & n23034;
  assign n31546 = n22846 | n23035;
  assign n31547 = (n23035 & n31476) | (n23035 & n31546) | (n31476 & n31546);
  assign n31548 = n22828 & n22835;
  assign n31549 = (n22828 & n31380) | (n22828 & n31548) | (n31380 & n31548);
  assign n31550 = n22828 | n22835;
  assign n31552 = n22829 & n31550;
  assign n31553 = (n22829 & n31380) | (n22829 & n31552) | (n31380 & n31552);
  assign n23040 = ~n31549 & n31553;
  assign n31554 = n23031 | n23040;
  assign n31555 = (n23040 & n31542) | (n23040 & n31554) | (n31542 & n31554);
  assign n35652 = n22488 | n22821;
  assign n35653 = n22713 | n35652;
  assign n31557 = n22821 | n31390;
  assign n31558 = (n31217 & n35653) | (n31217 & n31557) | (n35653 & n31557);
  assign n23044 = n22482 | n22712;
  assign n23045 = n22821 & n23044;
  assign n31559 = n22388 | n22713;
  assign n31561 = n23045 & n31559;
  assign n31562 = (n23045 & n31217) | (n23045 & n31561) | (n31217 & n31561);
  assign n23047 = n31558 & ~n31562;
  assign n23048 = n22822 & n23047;
  assign n31563 = n23048 | n31548;
  assign n31564 = n22828 | n23048;
  assign n31565 = (n31380 & n31563) | (n31380 & n31564) | (n31563 & n31564);
  assign n31567 = n22718 & n22815;
  assign n35654 = (n22709 & n22815) | (n22709 & n31567) | (n22815 & n31567);
  assign n31568 = (n31387 & n35654) | (n31387 & n31567) | (n35654 & n31567);
  assign n23052 = n22468 | n22727;
  assign n23053 = n22808 & n23052;
  assign n31569 = n22401 | n22728;
  assign n31571 = n23053 & n31569;
  assign n31572 = (n23053 & n31236) | (n23053 & n31571) | (n31236 & n31571);
  assign n31573 = n22808 | n31407;
  assign n35655 = n22728 | n22808;
  assign n35656 = n31393 | n35655;
  assign n31575 = (n31236 & n31573) | (n31236 & n35656) | (n31573 & n35656);
  assign n23056 = ~n31572 & n31575;
  assign n23057 = n22809 & n23056;
  assign n31576 = n22733 & n22801;
  assign n31577 = (n22801 & n35571) | (n22801 & n31576) | (n35571 & n31576);
  assign n31578 = n22733 | n22801;
  assign n31580 = n22802 & n31578;
  assign n31581 = (n22802 & n35571) | (n22802 & n31580) | (n35571 & n31580);
  assign n23062 = ~n31577 & n31581;
  assign n37853 = n22141 & ~n22454;
  assign n37854 = (n22140 & ~n22454) | (n22140 & n37853) | (~n22454 & n37853);
  assign n37748 = n22453 & n37854;
  assign n37439 = n31415 & n37748;
  assign n37440 = ~n22454 & n22737;
  assign n37441 = n22739 & n37440;
  assign n35659 = (n31086 & n37439) | (n31086 & n37441) | (n37439 & n37441);
  assign n31585 = (n22454 & n22736) | (n22454 & ~n35659) | (n22736 & ~n35659);
  assign n23069 = n22794 & n31585;
  assign n23066 = n22416 | n31421;
  assign n31582 = n22408 | n23066;
  assign n31586 = n23069 & n31582;
  assign n31587 = n23066 & n23069;
  assign n31588 = (n31244 & n31586) | (n31244 & n31587) | (n31586 & n31587);
  assign n31594 = n22451 & n22786;
  assign n35660 = (n22786 & n31417) | (n22786 & n31594) | (n31417 & n31594);
  assign n35661 = (n22786 & n31418) | (n22786 & n31594) | (n31418 & n31594);
  assign n35662 = (n31086 & n35660) | (n31086 & n35661) | (n35660 & n35661);
  assign n37442 = n22450 & n22787;
  assign n37443 = n22449 & n37442;
  assign n35664 = (n22786 & n22787) | (n22786 & n37443) | (n22787 & n37443);
  assign n35665 = (n22787 & n31417) | (n22787 & n35664) | (n31417 & n35664);
  assign n35666 = (n22787 & n31418) | (n22787 & n35664) | (n31418 & n35664);
  assign n35667 = (n31086 & n35665) | (n31086 & n35666) | (n35665 & n35666);
  assign n23077 = ~n35662 & n35667;
  assign n23086 = x142 & x144;
  assign n23087 = x141 & x145;
  assign n23088 = n23086 & n23087;
  assign n23089 = n23086 | n23087;
  assign n23090 = ~n23088 & n23089;
  assign n23091 = n22752 | n23090;
  assign n35668 = n22754 | n23091;
  assign n35669 = (n23091 & n35586) | (n23091 & n35668) | (n35586 & n35668);
  assign n35670 = (n23091 & n35588) | (n23091 & n35668) | (n35588 & n35668);
  assign n31619 = (n35438 & n35669) | (n35438 & n35670) | (n35669 & n35670);
  assign n23094 = n22753 & n23090;
  assign n37444 = n22752 & n22753;
  assign n37445 = n23090 & n37444;
  assign n37446 = (n23094 & n37429) | (n23094 & n37445) | (n37429 & n37445);
  assign n37447 = (n22429 & n23094) | (n22429 & n37445) | (n23094 & n37445);
  assign n37448 = (n31424 & n37446) | (n31424 & n37447) | (n37446 & n37447);
  assign n35673 = (n23094 & n35588) | (n23094 & n37445) | (n35588 & n37445);
  assign n31625 = (n35438 & n37448) | (n35438 & n35673) | (n37448 & n35673);
  assign n23096 = n31619 & ~n31625;
  assign n23097 = x140 & x146;
  assign n23098 = n23096 & n23097;
  assign n23099 = n23096 | n23097;
  assign n23100 = ~n23098 & n23099;
  assign n37449 = n22754 & n37429;
  assign n37450 = n22429 & n22754;
  assign n37451 = (n31424 & n37449) | (n31424 & n37450) | (n37449 & n37450);
  assign n31606 = n22754 & n35588;
  assign n31607 = (n35438 & n37451) | (n35438 & n31606) | (n37451 & n31606);
  assign n37452 = (n22755 & n22756) | (n22755 & n37429) | (n22756 & n37429);
  assign n37749 = n22429 & n22755;
  assign n37750 = (n22754 & n22755) | (n22754 & n37749) | (n22755 & n37749);
  assign n37454 = (n31424 & n37452) | (n31424 & n37750) | (n37452 & n37750);
  assign n35675 = (n22755 & n22756) | (n22755 & n35588) | (n22756 & n35588);
  assign n31613 = (n35438 & n37454) | (n35438 & n35675) | (n37454 & n35675);
  assign n23084 = ~n31607 & n31613;
  assign n35676 = n22437 | n23084;
  assign n35677 = (n22764 & n23084) | (n22764 & n35676) | (n23084 & n35676);
  assign n31626 = n23100 & ~n35677;
  assign n35678 = n22761 | n23084;
  assign n35679 = (n22438 & n23084) | (n22438 & n35678) | (n23084 & n35678);
  assign n31627 = n23100 & ~n35679;
  assign n35680 = (n31626 & n31627) | (n31626 & ~n35532) | (n31627 & ~n35532);
  assign n35681 = (n31626 & n31627) | (n31626 & ~n35531) | (n31627 & ~n35531);
  assign n35682 = (~n35269 & n35680) | (~n35269 & n35681) | (n35680 & n35681);
  assign n31629 = ~n23100 & n35677;
  assign n31630 = ~n23100 & n35679;
  assign n35683 = (n31629 & n31630) | (n31629 & n35532) | (n31630 & n35532);
  assign n35684 = (n31629 & n31630) | (n31629 & n35531) | (n31630 & n35531);
  assign n35685 = (n35269 & n35683) | (n35269 & n35684) | (n35683 & n35684);
  assign n23103 = n35682 | n35685;
  assign n23104 = x139 & x147;
  assign n23105 = n23103 & n23104;
  assign n23106 = n23103 | n23104;
  assign n23107 = ~n23105 & n23106;
  assign n31603 = n22768 | n22780;
  assign n31632 = n23107 | n31603;
  assign n31633 = n22768 | n23107;
  assign n31634 = (n35600 & n31632) | (n35600 & n31633) | (n31632 & n31633);
  assign n31635 = n23107 & n31603;
  assign n31636 = n22768 & n23107;
  assign n31637 = (n35600 & n31635) | (n35600 & n31636) | (n31635 & n31636);
  assign n23110 = n31634 & ~n31637;
  assign n23111 = x138 & x148;
  assign n23112 = n23110 | n23111;
  assign n23113 = n23110 & n23111;
  assign n23114 = n23112 & ~n23113;
  assign n23115 = x137 & x149;
  assign n23116 = n23114 & n23115;
  assign n23117 = n23114 | n23115;
  assign n23118 = ~n23116 & n23117;
  assign n31787 = n22451 | n22784;
  assign n35686 = (n22784 & n22786) | (n22784 & n31787) | (n22786 & n31787);
  assign n31638 = n23118 | n35686;
  assign n31601 = n22784 | n22786;
  assign n31639 = n23118 | n31601;
  assign n31640 = (n31419 & n31638) | (n31419 & n31639) | (n31638 & n31639);
  assign n31641 = n23118 & n35686;
  assign n31642 = n23118 & n31601;
  assign n31643 = (n31419 & n31641) | (n31419 & n31642) | (n31641 & n31642);
  assign n23121 = n31640 & ~n31643;
  assign n23122 = x136 & x150;
  assign n23123 = n23121 | n23122;
  assign n23124 = n23121 & n23122;
  assign n23125 = n23123 & ~n23124;
  assign n31644 = ~n23077 & n23125;
  assign n31645 = ~n31588 & n31644;
  assign n31646 = n23077 & ~n23125;
  assign n31647 = (~n23125 & n31588) | (~n23125 & n31646) | (n31588 & n31646);
  assign n23128 = n31645 | n31647;
  assign n23129 = x135 & x151;
  assign n23130 = n23128 & n23129;
  assign n23131 = n23128 | n23129;
  assign n23132 = ~n23130 & n23131;
  assign n23064 = n31421 | n22794;
  assign n23065 = n35580 | n23064;
  assign n37455 = n22795 & ~n23066;
  assign n37456 = (n22795 & ~n23069) | (n22795 & n37455) | (~n23069 & n37455);
  assign n35688 = n22795 & ~n31586;
  assign n35689 = (~n31244 & n37456) | (~n31244 & n35688) | (n37456 & n35688);
  assign n31590 = n23065 & n35689;
  assign n31591 = n31576 | n31590;
  assign n31648 = n23132 | n31591;
  assign n31592 = n22801 | n31590;
  assign n31649 = n23132 | n31592;
  assign n31650 = (n35571 & n31648) | (n35571 & n31649) | (n31648 & n31649);
  assign n31651 = n23132 & n31591;
  assign n31652 = n23132 & n31592;
  assign n31653 = (n35571 & n31651) | (n35571 & n31652) | (n31651 & n31652);
  assign n23135 = n31650 & ~n31653;
  assign n23136 = x134 & x152;
  assign n23137 = n23135 | n23136;
  assign n23138 = n23135 & n23136;
  assign n23139 = n23137 & ~n23138;
  assign n31654 = ~n23062 & n23139;
  assign n31655 = ~n31572 & n31654;
  assign n31656 = n23062 & ~n23139;
  assign n31657 = (~n23139 & n31572) | (~n23139 & n31656) | (n31572 & n31656);
  assign n23142 = n31655 | n31657;
  assign n23143 = x133 & x153;
  assign n23144 = n23142 & n23143;
  assign n23145 = n23142 | n23143;
  assign n23146 = ~n23144 & n23145;
  assign n31658 = n23057 | n23146;
  assign n31659 = n31568 | n31658;
  assign n31660 = n23057 & n23146;
  assign n31661 = (n23146 & n31568) | (n23146 & n31660) | (n31568 & n31660);
  assign n23149 = n31659 & ~n31661;
  assign n23150 = x132 & x154;
  assign n23151 = n23149 | n23150;
  assign n23152 = n23149 & n23150;
  assign n23153 = n23151 & ~n23152;
  assign n31663 = n22718 | n22815;
  assign n35690 = n22709 | n31663;
  assign n31664 = (n31387 & n35690) | (n31387 & n31663) | (n35690 & n31663);
  assign n35691 = n22720 & ~n35654;
  assign n35692 = n22720 & ~n31567;
  assign n35693 = (~n31387 & n35691) | (~n31387 & n35692) | (n35691 & n35692);
  assign n23156 = n31664 & n35693;
  assign n31665 = ~n23153 & n23156;
  assign n31666 = (~n23153 & n31562) | (~n23153 & n31665) | (n31562 & n31665);
  assign n31667 = n23153 & ~n23156;
  assign n31668 = ~n31562 & n31667;
  assign n23160 = n31666 | n31668;
  assign n23161 = x131 & x155;
  assign n23162 = n23160 & n23161;
  assign n23163 = n23160 | n23161;
  assign n23164 = ~n23162 & n23163;
  assign n23165 = n31565 | n23164;
  assign n23166 = n31565 & n23164;
  assign n23167 = n23165 & ~n23166;
  assign n23168 = x130 & x156;
  assign n23169 = n23167 | n23168;
  assign n23170 = n23167 & n23168;
  assign n23171 = n23169 & ~n23170;
  assign n23172 = ~n31555 & n23171;
  assign n23173 = n31555 & ~n23171;
  assign n23174 = n23172 | n23173;
  assign n23175 = x129 & x157;
  assign n23176 = n23174 & n23175;
  assign n23177 = n23174 | n23175;
  assign n23178 = ~n23176 & n23177;
  assign n23179 = n31547 | n23178;
  assign n23180 = n31547 & n23178;
  assign n23181 = n23179 & ~n23180;
  assign n23182 = x128 & x158;
  assign n23183 = ~n23181 & n23182;
  assign n23184 = n23181 & ~n23182;
  assign n23185 = n23183 | n23184;
  assign n23186 = ~n31540 & n23185;
  assign n23187 = n31540 & ~n23185;
  assign n23188 = n23186 | n23187;
  assign n23189 = x127 & x159;
  assign n23190 = n23188 & n23189;
  assign n23191 = n23188 | n23189;
  assign n23192 = ~n23190 & n23191;
  assign n23193 = n31536 | n23192;
  assign n23194 = n31536 & n23192;
  assign n23195 = n23193 & ~n23194;
  assign n23196 = x126 & x160;
  assign n23197 = ~n23195 & n23196;
  assign n23198 = n23195 & ~n23196;
  assign n23199 = n23197 | n23198;
  assign n23200 = n23014 | n23199;
  assign n23201 = n23014 & n23199;
  assign n23202 = n23200 & ~n23201;
  assign n23203 = n23004 & n23202;
  assign n23204 = n23004 | n23202;
  assign n23205 = ~n23203 & n23204;
  assign n23206 = n22685 | n22875;
  assign n31669 = n22671 | n23206;
  assign n31670 = (n22670 & n23206) | (n22670 & n31669) | (n23206 & n31669);
  assign n23208 = ~n31526 & n31670;
  assign n23209 = n22876 & n23208;
  assign n23210 = n31522 | n23209;
  assign n23211 = n23205 | n23210;
  assign n23212 = n23205 & n23210;
  assign n23213 = n23211 & ~n23212;
  assign n23214 = x124 & x162;
  assign n23215 = n23213 | n23214;
  assign n23216 = n23213 & n23214;
  assign n23217 = n23215 & ~n23216;
  assign n23218 = n23003 | n23217;
  assign n23219 = n23003 & n23217;
  assign n23220 = n23218 & ~n23219;
  assign n23221 = x123 & x163;
  assign n23222 = n23220 | n23221;
  assign n23223 = n23220 & n23221;
  assign n23224 = n23222 & ~n23223;
  assign n31671 = n22889 | n31359;
  assign n31672 = n22667 | n22889;
  assign n31673 = (n31190 & n31671) | (n31190 & n31672) | (n31671 & n31672);
  assign n23227 = n22890 & ~n31520;
  assign n23228 = n31673 & n23227;
  assign n31674 = n22896 | n23228;
  assign n31675 = (n23228 & n31487) | (n23228 & n31674) | (n31487 & n31674);
  assign n23230 = ~n23224 & n31675;
  assign n23231 = n23224 & ~n31675;
  assign n23232 = n23230 | n23231;
  assign n23233 = x122 & x164;
  assign n23234 = n23232 & ~n23233;
  assign n23235 = ~n23232 & n23233;
  assign n23236 = n23234 | n23235;
  assign n23237 = n22896 | n31487;
  assign n31676 = (n22897 & n22898) | (n22897 & ~n31487) | (n22898 & ~n31487);
  assign n23239 = n23237 & n31676;
  assign n31677 = n23239 | n31512;
  assign n31678 = n22908 | n23239;
  assign n31679 = (n31350 & n31677) | (n31350 & n31678) | (n31677 & n31678);
  assign n23241 = n23236 & n31679;
  assign n23242 = n23236 | n31679;
  assign n23243 = ~n23241 & n23242;
  assign n31680 = ~n22996 & n23243;
  assign n31681 = ~n31511 & n31680;
  assign n31682 = n22996 & ~n23243;
  assign n31683 = (~n23243 & n31511) | (~n23243 & n31682) | (n31511 & n31682);
  assign n23246 = n31681 | n31683;
  assign n23247 = x121 & x165;
  assign n23248 = n23246 & n23247;
  assign n23249 = n23246 | n23247;
  assign n23250 = ~n23248 & n23249;
  assign n31684 = n22924 & n23250;
  assign n31685 = (n23250 & n31497) | (n23250 & n31684) | (n31497 & n31684);
  assign n31686 = n22924 | n23250;
  assign n31687 = n31497 | n31686;
  assign n23253 = ~n31685 & n31687;
  assign n23254 = n22990 | n23253;
  assign n23255 = n22990 & n23253;
  assign n23256 = n23254 & ~n23255;
  assign n31688 = n22930 & n22931;
  assign n31689 = (n22930 & n31501) | (n22930 & n31688) | (n31501 & n31688);
  assign n23259 = n23256 & ~n31689;
  assign n23260 = ~n23256 & n31689;
  assign n23261 = n23259 | n23260;
  assign n23262 = x119 & x167;
  assign n23263 = n23261 | n23262;
  assign n23264 = n23261 & n23262;
  assign n23265 = n23263 & ~n23264;
  assign n31690 = n22939 & n22940;
  assign n31691 = (n22939 & n31503) | (n22939 & n31690) | (n31503 & n31690);
  assign n23268 = n23265 & ~n31691;
  assign n23269 = ~n23265 & n31691;
  assign n23270 = n23268 | n23269;
  assign n23271 = x118 & x168;
  assign n23272 = n23270 | n23271;
  assign n23273 = n23270 & n23271;
  assign n23274 = n23272 & ~n23273;
  assign n23275 = ~n22989 & n23274;
  assign n23276 = n22989 & ~n23274;
  assign n23277 = n23275 | n23276;
  assign n31692 = n22954 & n22955;
  assign n31693 = (n22955 & n31344) | (n22955 & n31692) | (n31344 & n31692);
  assign n23280 = n23277 & ~n31693;
  assign n23281 = ~n23277 & n31693;
  assign n23282 = n23280 | n23281;
  assign n23283 = x116 & x170;
  assign n23284 = n23282 | n23283;
  assign n23285 = n23282 & n23283;
  assign n23286 = n23284 & ~n23285;
  assign n31694 = n22960 & n22961;
  assign n31695 = (n22960 & n31342) | (n22960 & n31694) | (n31342 & n31694);
  assign n23289 = n23286 & ~n31695;
  assign n23290 = ~n23286 & n31695;
  assign n23291 = n23289 | n23290;
  assign n23292 = x115 & x171;
  assign n23293 = n23291 | n23292;
  assign n23294 = n23291 & n23292;
  assign n23295 = n23293 & ~n23294;
  assign n23296 = ~n31342 & n22962;
  assign n23297 = n31342 & ~n22962;
  assign n23298 = n23296 | n23297;
  assign n23299 = n22645 & n23298;
  assign n23300 = n22969 | n23299;
  assign n23301 = n22645 | n23298;
  assign n23302 = n23300 & n23301;
  assign n23303 = n23295 & ~n23302;
  assign n23304 = ~n23295 & n23302;
  assign n23305 = n23303 | n23304;
  assign n23306 = x114 & x172;
  assign n23307 = n23305 | n23306;
  assign n23308 = n23305 & n23306;
  assign n23309 = n23307 & ~n23308;
  assign n23310 = n22640 | n22975;
  assign n23311 = n22974 & n23310;
  assign n23312 = n23309 & ~n23311;
  assign n23313 = ~n23309 & n23311;
  assign n23314 = n23312 | n23313;
  assign n23315 = x113 & x173;
  assign n23316 = n23314 | n23315;
  assign n23317 = n23314 & n23315;
  assign n23318 = n23316 & ~n23317;
  assign n23319 = ~n22981 & n23318;
  assign n23320 = n22981 & ~n23318;
  assign n23321 = n23319 | n23320;
  assign n23322 = x112 & x174;
  assign n23323 = n23321 & n23322;
  assign n23324 = n23321 | n23322;
  assign n23325 = ~n23323 & n23324;
  assign n31696 = n23284 & n23285;
  assign n31697 = (n23284 & n31695) | (n23284 & n31696) | (n31695 & n31696);
  assign n23328 = x116 & x171;
  assign n23329 = n31697 & n23328;
  assign n23330 = n31697 | n23328;
  assign n23331 = ~n23329 & n23330;
  assign n23332 = x117 & x170;
  assign n23333 = ~n31509 & n23274;
  assign n23334 = n31509 & ~n23274;
  assign n23335 = n23333 | n23334;
  assign n23338 = n22986 | n23335;
  assign n23336 = n22986 & n23335;
  assign n31698 = n23336 & n23338;
  assign n31699 = (n23338 & n31693) | (n23338 & n31698) | (n31693 & n31698);
  assign n23340 = x118 & x169;
  assign n31700 = n23272 & n23273;
  assign n31701 = (n23272 & n31509) | (n23272 & n31700) | (n31509 & n31700);
  assign n23343 = x121 & x166;
  assign n23345 = x122 & x165;
  assign n23347 = n23232 | n31679;
  assign n31704 = (n23233 & n23235) | (n23233 & ~n31679) | (n23235 & ~n31679);
  assign n23350 = n23347 & n31704;
  assign n31702 = n22996 & n23243;
  assign n31705 = n23350 | n31702;
  assign n31706 = n23243 | n23350;
  assign n31707 = (n31511 & n31705) | (n31511 & n31706) | (n31705 & n31706);
  assign n31708 = n23002 & n23213;
  assign n31709 = (n23213 & n31520) | (n23213 & n31708) | (n31520 & n31708);
  assign n31710 = n23202 | n23209;
  assign n31711 = n31522 | n31710;
  assign n23354 = n22674 | n23209;
  assign n23355 = n31355 | n23354;
  assign n23356 = n22876 | n23208;
  assign n23357 = n23202 & n23356;
  assign n23358 = n23355 & n23357;
  assign n23359 = n31711 & ~n23358;
  assign n23360 = n23004 & n23359;
  assign n23361 = n31709 | n23360;
  assign n31712 = n23013 & n23195;
  assign n23367 = n31480 | n31534;
  assign n31718 = n22858 | n31530;
  assign n31719 = (n22858 & ~n23019) | (n22858 & n31718) | (~n23019 & n31718);
  assign n23369 = n23188 & n31719;
  assign n23370 = n23367 & n23369;
  assign n31720 = n23188 | n31535;
  assign n31721 = n23188 | n31534;
  assign n31722 = (n31480 & n31720) | (n31480 & n31721) | (n31720 & n31721);
  assign n31723 = n23189 & n31722;
  assign n31724 = ~n23370 & n31723;
  assign n31725 = n31712 | n31724;
  assign n31726 = n23195 | n31724;
  assign n31727 = (n31526 & n31725) | (n31526 & n31726) | (n31725 & n31726);
  assign n23376 = n23035 | n23174;
  assign n31728 = n22846 | n23376;
  assign n31729 = (n23376 & n31476) | (n23376 & n31728) | (n31476 & n31728);
  assign n23379 = n22840 | n23034;
  assign n23380 = n23174 & n23379;
  assign n31730 = n23035 & n23380;
  assign n31731 = (n23380 & n31476) | (n23380 & n31730) | (n31476 & n31730);
  assign n23382 = n31729 & ~n31731;
  assign n23383 = n23175 & n23382;
  assign n31732 = n23181 | n23383;
  assign n31733 = (n23383 & n31540) | (n23383 & n31732) | (n31540 & n31732);
  assign n23385 = x129 & x158;
  assign n35694 = n23167 & n31554;
  assign n35695 = n23040 & n23167;
  assign n35696 = (n31542 & n35694) | (n31542 & n35695) | (n35694 & n35695);
  assign n35697 = (n23168 & n23170) | (n23168 & n31554) | (n23170 & n31554);
  assign n37457 = n23040 & n23168;
  assign n37458 = (n23167 & n23168) | (n23167 & n37457) | (n23168 & n37457);
  assign n35699 = (n31542 & n35697) | (n31542 & n37458) | (n35697 & n37458);
  assign n23389 = ~n35696 & n35699;
  assign n35700 = n23160 | n31564;
  assign n35701 = n23160 | n31563;
  assign n35702 = (n31380 & n35700) | (n31380 & n35701) | (n35700 & n35701);
  assign n23392 = n22822 | n23047;
  assign n23393 = n23160 & n23392;
  assign n31735 = n22835 | n23048;
  assign n31737 = n23393 & n31735;
  assign n31738 = (n23393 & n31380) | (n23393 & n31737) | (n31380 & n31737);
  assign n31739 = n23161 & ~n31738;
  assign n31740 = n35702 & n31739;
  assign n31741 = n23167 | n31740;
  assign n35703 = (n31554 & n31740) | (n31554 & n31741) | (n31740 & n31741);
  assign n35704 = (n23040 & n31740) | (n23040 & n31741) | (n31740 & n31741);
  assign n35705 = (n31542 & n35703) | (n31542 & n35704) | (n35703 & n35704);
  assign n31743 = n23149 & n23156;
  assign n31744 = (n23149 & n31562) | (n23149 & n31743) | (n31562 & n31743);
  assign n35706 = n23150 & n23156;
  assign n35707 = (n23149 & n23150) | (n23149 & n35706) | (n23150 & n35706);
  assign n31748 = (n23150 & n31562) | (n23150 & n35707) | (n31562 & n35707);
  assign n23402 = ~n31744 & n31748;
  assign n31749 = n23057 | n31399;
  assign n31750 = n22718 | n23057;
  assign n31751 = (n31387 & n31749) | (n31387 & n31750) | (n31749 & n31750);
  assign n23417 = n31590 | n23128;
  assign n31765 = n23417 | n31576;
  assign n35719 = n23128 | n31592;
  assign n31767 = (n35571 & n31765) | (n35571 & n35719) | (n31765 & n35719);
  assign n37459 = ~n22795 & n23066;
  assign n37460 = n23069 & n37459;
  assign n35721 = ~n22795 & n31586;
  assign n35722 = (n31244 & n37460) | (n31244 & n35721) | (n37460 & n35721);
  assign n31769 = (n22795 & n23065) | (n22795 & ~n35722) | (n23065 & ~n35722);
  assign n23422 = n23128 & n31769;
  assign n23419 = n22733 | n31590;
  assign n31770 = n23419 & n23422;
  assign n31771 = (n23422 & n35571) | (n23422 & n31770) | (n35571 & n31770);
  assign n23424 = n31767 & ~n31771;
  assign n23425 = n23129 & n23424;
  assign n31757 = n23062 & n23135;
  assign n31772 = n23425 | n31757;
  assign n31773 = n23135 | n23425;
  assign n35723 = (n31571 & n31772) | (n31571 & n31773) | (n31772 & n31773);
  assign n35724 = (n23053 & n31772) | (n23053 & n31773) | (n31772 & n31773);
  assign n35725 = (n31236 & n35723) | (n31236 & n35724) | (n35723 & n35724);
  assign n35738 = n23098 | n23099;
  assign n35739 = (n23098 & n35677) | (n23098 & n35738) | (n35677 & n35738);
  assign n35740 = (n23098 & n35679) | (n23098 & n35738) | (n35679 & n35738);
  assign n35741 = (n35532 & n35739) | (n35532 & n35740) | (n35739 & n35740);
  assign n35742 = (n35531 & n35739) | (n35531 & n35740) | (n35739 & n35740);
  assign n35743 = (n35269 & n35741) | (n35269 & n35742) | (n35741 & n35742);
  assign n23441 = x140 & x147;
  assign n23442 = x141 & x146;
  assign n23444 = x143 & x144;
  assign n23445 = x142 & x145;
  assign n23446 = n23444 & ~n23445;
  assign n23447 = ~n23444 & n23445;
  assign n23448 = n23446 | n23447;
  assign n35747 = n23088 & n23448;
  assign n37466 = (n23448 & n35747) | (n23448 & n37445) | (n35747 & n37445);
  assign n37461 = n22753 | n23088;
  assign n37462 = (n23088 & n23090) | (n23088 & n37461) | (n23090 & n37461);
  assign n37464 = n23448 & n37462;
  assign n37465 = (n35586 & n37466) | (n35586 & n37464) | (n37466 & n37464);
  assign n37467 = (n23094 & n23448) | (n23094 & n35747) | (n23448 & n35747);
  assign n37468 = (n35588 & n37466) | (n35588 & n37467) | (n37466 & n37467);
  assign n31805 = (n35438 & n37465) | (n35438 & n37468) | (n37465 & n37468);
  assign n35749 = n23088 | n23448;
  assign n37472 = n35749 | n37445;
  assign n37470 = n23448 | n37462;
  assign n37471 = (n35586 & n37472) | (n35586 & n37470) | (n37472 & n37470);
  assign n37473 = n23094 | n35749;
  assign n37474 = (n35588 & n37472) | (n35588 & n37473) | (n37472 & n37473);
  assign n31808 = (n35438 & n37471) | (n35438 & n37474) | (n37471 & n37474);
  assign n23451 = ~n31805 & n31808;
  assign n23452 = n23442 & n23451;
  assign n23453 = n23442 | n23451;
  assign n23454 = ~n23452 & n23453;
  assign n23455 = ~n23441 & n23454;
  assign n23456 = n23441 & ~n23454;
  assign n23457 = n23455 | n23456;
  assign n23458 = n35743 & n23457;
  assign n23459 = n35743 | n23457;
  assign n23460 = ~n23458 & n23459;
  assign n23461 = n23105 | n23460;
  assign n35751 = n23107 | n23461;
  assign n35752 = (n23461 & n31603) | (n23461 & n35751) | (n31603 & n35751);
  assign n31810 = n23461 | n31636;
  assign n31811 = (n35600 & n35752) | (n35600 & n31810) | (n35752 & n31810);
  assign n23464 = n23106 & n23460;
  assign n31813 = n22768 | n23105;
  assign n35753 = n22780 | n31813;
  assign n31815 = n23464 & n35753;
  assign n31816 = n23464 & n31813;
  assign n31817 = (n35600 & n31815) | (n35600 & n31816) | (n31815 & n31816);
  assign n23466 = n31811 & ~n31817;
  assign n23467 = x139 & x148;
  assign n23468 = n23466 & n23467;
  assign n23469 = n23466 | n23467;
  assign n23470 = ~n23468 & n23469;
  assign n23471 = x138 & x149;
  assign n23472 = n23470 & n23471;
  assign n23473 = n23470 | n23471;
  assign n23474 = ~n23472 & n23473;
  assign n23434 = n22785 & n23114;
  assign n35754 = n23113 | n31787;
  assign n35755 = (n23113 & n23434) | (n23113 & n35754) | (n23434 & n35754);
  assign n35756 = n22785 | n23113;
  assign n35757 = (n23113 & n23114) | (n23113 & n35756) | (n23114 & n35756);
  assign n35758 = (n31417 & n35755) | (n31417 & n35757) | (n35755 & n35757);
  assign n35759 = (n31418 & n35755) | (n31418 & n35757) | (n35755 & n35757);
  assign n35760 = (n31086 & n35758) | (n31086 & n35759) | (n35758 & n35759);
  assign n23476 = ~n23474 & n35760;
  assign n23477 = n23474 & ~n35760;
  assign n23478 = n23476 | n23477;
  assign n23479 = x137 & x150;
  assign n23480 = n23478 & n23479;
  assign n23481 = n23478 | n23479;
  assign n23482 = ~n23480 & n23481;
  assign n31784 = n23114 | n35686;
  assign n31785 = n23114 | n31601;
  assign n35761 = (n31417 & n31784) | (n31417 & n31785) | (n31784 & n31785);
  assign n35762 = (n31418 & n31784) | (n31418 & n31785) | (n31784 & n31785);
  assign n35763 = (n31086 & n35761) | (n31086 & n35762) | (n35761 & n35762);
  assign n31789 = n23434 & n31787;
  assign n35764 = (n23434 & n31417) | (n23434 & n31789) | (n31417 & n31789);
  assign n35765 = (n23434 & n31418) | (n23434 & n31789) | (n31418 & n31789);
  assign n35766 = (n31086 & n35764) | (n31086 & n35765) | (n35764 & n35765);
  assign n23436 = n35763 & ~n35766;
  assign n23437 = n23115 & n23436;
  assign n31792 = n23121 | n23437;
  assign n31821 = n23482 & ~n31792;
  assign n31775 = n23077 & n23121;
  assign n31791 = n23437 | n31775;
  assign n31822 = n23482 & ~n31791;
  assign n31823 = (~n31588 & n31821) | (~n31588 & n31822) | (n31821 & n31822);
  assign n31824 = ~n23482 & n31792;
  assign n31825 = ~n23482 & n31791;
  assign n31826 = (n31588 & n31824) | (n31588 & n31825) | (n31824 & n31825);
  assign n23485 = n31823 | n31826;
  assign n23486 = x136 & x151;
  assign n23487 = n23485 | n23486;
  assign n23488 = n23485 & n23486;
  assign n23489 = n23487 & ~n23488;
  assign n35726 = (n23121 & n31587) | (n23121 & n31775) | (n31587 & n31775);
  assign n35727 = (n23121 & n31586) | (n23121 & n31775) | (n31586 & n31775);
  assign n35728 = (n31244 & n35726) | (n31244 & n35727) | (n35726 & n35727);
  assign n35729 = n23077 & n23122;
  assign n35730 = (n23121 & n23122) | (n23121 & n35729) | (n23122 & n35729);
  assign n35731 = (n23122 & n31587) | (n23122 & n35730) | (n31587 & n35730);
  assign n35732 = (n23122 & n31586) | (n23122 & n35730) | (n31586 & n35730);
  assign n35733 = (n31244 & n35731) | (n31244 & n35732) | (n35731 & n35732);
  assign n23430 = ~n35728 & n35733;
  assign n35734 = n23419 | n23430;
  assign n35735 = (n23422 & n23430) | (n23422 & n35734) | (n23430 & n35734);
  assign n35767 = n23489 & ~n35735;
  assign n35736 = n23430 | n31769;
  assign n35737 = (n23128 & n23430) | (n23128 & n35736) | (n23430 & n35736);
  assign n35768 = n23489 & ~n35737;
  assign n35769 = (~n35571 & n35767) | (~n35571 & n35768) | (n35767 & n35768);
  assign n35770 = ~n23489 & n35735;
  assign n35771 = ~n23489 & n35737;
  assign n35772 = (n35571 & n35770) | (n35571 & n35771) | (n35770 & n35771);
  assign n23492 = n35769 | n35772;
  assign n23493 = x135 & x152;
  assign n23494 = n23492 & n23493;
  assign n23495 = n23492 | n23493;
  assign n23496 = ~n23494 & n23495;
  assign n23497 = n35725 | n23496;
  assign n23498 = n35725 & n23496;
  assign n23499 = n23497 & ~n23498;
  assign n23500 = x134 & x153;
  assign n23501 = n23499 | n23500;
  assign n23502 = n23499 & n23500;
  assign n23503 = n23501 & ~n23502;
  assign n23405 = n22809 | n23056;
  assign n23406 = n23142 & n23405;
  assign n35713 = (n23135 & n31571) | (n23135 & n31757) | (n31571 & n31757);
  assign n35714 = (n23053 & n23135) | (n23053 & n31757) | (n23135 & n31757);
  assign n35715 = (n31236 & n35713) | (n31236 & n35714) | (n35713 & n35714);
  assign n31759 = n23062 | n23135;
  assign n31761 = n23136 & n31759;
  assign n35716 = (n23136 & n31571) | (n23136 & n31761) | (n31571 & n31761);
  assign n35717 = (n23053 & n23136) | (n23053 & n31761) | (n23136 & n31761);
  assign n35718 = (n31236 & n35716) | (n31236 & n35717) | (n35716 & n35717);
  assign n23415 = ~n35715 & n35718;
  assign n31763 = n23406 | n23415;
  assign n35773 = n23503 & ~n31763;
  assign n35774 = ~n23415 & n23503;
  assign n35775 = (~n31751 & n35773) | (~n31751 & n35774) | (n35773 & n35774);
  assign n35776 = ~n23503 & n31763;
  assign n35777 = n23415 & ~n23503;
  assign n35778 = (n31751 & n35776) | (n31751 & n35777) | (n35776 & n35777);
  assign n23506 = n35775 | n35778;
  assign n23507 = x133 & x154;
  assign n23508 = n23506 & n23507;
  assign n23509 = n23506 | n23507;
  assign n23510 = ~n23508 & n23509;
  assign n23407 = n31751 & n23406;
  assign n31752 = n23057 | n23142;
  assign n35708 = n31752 | n35654;
  assign n35709 = n31567 | n31752;
  assign n35710 = (n31387 & n35708) | (n31387 & n35709) | (n35708 & n35709);
  assign n35711 = n23143 & n35710;
  assign n35712 = ~n23407 & n35711;
  assign n31754 = n35712 | n31743;
  assign n35779 = n23510 | n31754;
  assign n31755 = n23149 | n35712;
  assign n35780 = n23510 | n31755;
  assign n35781 = (n31562 & n35779) | (n31562 & n35780) | (n35779 & n35780);
  assign n35782 = n23510 & n31754;
  assign n35783 = n23510 & n31755;
  assign n35784 = (n31562 & n35782) | (n31562 & n35783) | (n35782 & n35783);
  assign n23513 = n35781 & ~n35784;
  assign n23514 = x132 & x155;
  assign n23515 = n23513 | n23514;
  assign n23516 = n23513 & n23514;
  assign n23517 = n23515 & ~n23516;
  assign n35785 = ~n23402 & n23517;
  assign n35786 = ~n31738 & n35785;
  assign n35787 = n23402 & ~n23517;
  assign n35788 = (~n23517 & n31738) | (~n23517 & n35787) | (n31738 & n35787);
  assign n23520 = n35786 | n35788;
  assign n23521 = x131 & x156;
  assign n23522 = n23520 & n23521;
  assign n23523 = n23520 | n23521;
  assign n23524 = ~n23522 & n23523;
  assign n23525 = n35705 | n23524;
  assign n23526 = n35705 & n23524;
  assign n23527 = n23525 & ~n23526;
  assign n23528 = x130 & x157;
  assign n23529 = ~n23527 & n23528;
  assign n23530 = n23527 & ~n23528;
  assign n23531 = n23529 | n23530;
  assign n35789 = n23389 | n23531;
  assign n35790 = n31731 | n35789;
  assign n35791 = n23389 & n23531;
  assign n35792 = (n23531 & n31731) | (n23531 & n35791) | (n31731 & n35791);
  assign n23534 = n35790 & ~n35792;
  assign n23535 = n23385 & n23534;
  assign n23536 = n23385 | n23534;
  assign n23537 = ~n23535 & n23536;
  assign n23538 = ~n31733 & n23537;
  assign n23539 = n31733 & ~n23537;
  assign n23540 = n23538 | n23539;
  assign n23541 = x128 & x159;
  assign n23542 = n23540 | n23541;
  assign n23543 = n23540 & n23541;
  assign n23544 = n23542 & ~n23543;
  assign n35793 = n23181 | n35651;
  assign n35794 = n23026 | n23181;
  assign n35795 = (n23016 & n35793) | (n23016 & n35794) | (n35793 & n35794);
  assign n31827 = (n23182 & n23183) | (n23182 & ~n31540) | (n23183 & ~n31540);
  assign n23547 = n35795 & n31827;
  assign n31828 = n23369 | n23547;
  assign n31829 = (n23367 & n23547) | (n23367 & n31828) | (n23547 & n31828);
  assign n23549 = ~n23544 & n31829;
  assign n23550 = n23544 & ~n31829;
  assign n23551 = n23549 | n23550;
  assign n23552 = x127 & x160;
  assign n23553 = ~n23551 & n23552;
  assign n23554 = n23551 & ~n23552;
  assign n23555 = n23553 | n23554;
  assign n23556 = n31727 & ~n23555;
  assign n23557 = ~n31727 & n23555;
  assign n23558 = n23556 | n23557;
  assign n31713 = (n23195 & n31526) | (n23195 & n31712) | (n31526 & n31712);
  assign n35796 = n23013 & n23196;
  assign n35797 = (n23195 & n23196) | (n23195 & n35796) | (n23196 & n35796);
  assign n31717 = (n23196 & n31526) | (n23196 & n35797) | (n31526 & n35797);
  assign n23365 = ~n31713 & n31717;
  assign n31830 = n23365 & n23558;
  assign n31831 = (n23358 & n23558) | (n23358 & n31830) | (n23558 & n31830);
  assign n31832 = n23365 | n23558;
  assign n31833 = n23358 | n31832;
  assign n23561 = ~n31831 & n31833;
  assign n23562 = x126 & x161;
  assign n23563 = n23561 & n23562;
  assign n23564 = n23561 | n23562;
  assign n23565 = ~n23563 & n23564;
  assign n23566 = x125 & x162;
  assign n23567 = n23565 & n23566;
  assign n23568 = n23565 | n23566;
  assign n23569 = ~n23567 & n23568;
  assign n23570 = n23361 | n23569;
  assign n23571 = n23361 & n23569;
  assign n23572 = n23570 & ~n23571;
  assign n23573 = x124 & x163;
  assign n23574 = n23572 | n23573;
  assign n23575 = n23572 & n23573;
  assign n23576 = n23574 & ~n23575;
  assign n31834 = n23220 & n31674;
  assign n31835 = n23220 & n23228;
  assign n31836 = (n31487 & n31834) | (n31487 & n31835) | (n31834 & n31835);
  assign n31837 = n23002 | n23213;
  assign n31838 = n31520 | n31837;
  assign n23579 = n23214 & ~n31709;
  assign n23580 = n31838 & n23579;
  assign n23581 = n31836 | n23580;
  assign n23582 = ~n23576 & n23581;
  assign n23583 = n23576 & ~n23581;
  assign n23584 = n23582 | n23583;
  assign n23585 = x123 & x164;
  assign n23586 = n23584 & n23585;
  assign n23587 = n23584 | n23585;
  assign n23588 = ~n23586 & n23587;
  assign n31839 = n23220 | n31674;
  assign n31840 = n23220 | n23228;
  assign n31841 = (n31487 & n31839) | (n31487 & n31840) | (n31839 & n31840);
  assign n23590 = n23221 & ~n31836;
  assign n23591 = n31841 & n23590;
  assign n31842 = n23232 | n23591;
  assign n31843 = (n23591 & n31679) | (n23591 & n31842) | (n31679 & n31842);
  assign n23593 = ~n23588 & n31843;
  assign n23594 = n23588 & ~n31843;
  assign n23595 = n23593 | n23594;
  assign n23596 = n31707 & n23595;
  assign n23597 = n31707 | n23595;
  assign n23598 = ~n23596 & n23597;
  assign n23599 = ~n23345 & n23598;
  assign n23600 = n23345 & ~n23598;
  assign n23601 = n23599 | n23600;
  assign n31844 = n23248 & n23601;
  assign n31845 = (n23601 & n31685) | (n23601 & n31844) | (n31685 & n31844);
  assign n31846 = n23248 | n23601;
  assign n31847 = n31685 | n31846;
  assign n23604 = ~n31845 & n31847;
  assign n23605 = n23343 | n23604;
  assign n23606 = n23343 & n23604;
  assign n23607 = n23605 & ~n23606;
  assign n31848 = n23254 & n23255;
  assign n31849 = (n23254 & n31689) | (n23254 & n31848) | (n31689 & n31848);
  assign n23610 = n23607 & ~n31849;
  assign n23611 = ~n23607 & n31849;
  assign n23612 = n23610 | n23611;
  assign n23613 = x120 & x167;
  assign n23614 = n23612 | n23613;
  assign n23615 = n23612 & n23613;
  assign n23616 = n23614 & ~n23615;
  assign n31850 = n23263 & n23264;
  assign n31851 = (n23263 & n31691) | (n23263 & n31850) | (n31691 & n31850);
  assign n23619 = n23616 & ~n31851;
  assign n23620 = ~n23616 & n31851;
  assign n23621 = n23619 | n23620;
  assign n23622 = x119 & x168;
  assign n23623 = n23621 | n23622;
  assign n23624 = n23621 & n23622;
  assign n23625 = n23623 & ~n23624;
  assign n23626 = ~n31701 & n23625;
  assign n23627 = n31701 & ~n23625;
  assign n23628 = n23626 | n23627;
  assign n23629 = n23340 & n23628;
  assign n23630 = n23340 | n23628;
  assign n23631 = ~n23629 & n23630;
  assign n23632 = n31699 & n23631;
  assign n23633 = n31699 | n23631;
  assign n23634 = ~n23632 & n23633;
  assign n23635 = n23332 | n23634;
  assign n23636 = n23332 & n23634;
  assign n23637 = n23635 & ~n23636;
  assign n23638 = ~n23331 & n23637;
  assign n23639 = n23331 & ~n23637;
  assign n23640 = n23638 | n23639;
  assign n31852 = n23293 & n23294;
  assign n31853 = (n23293 & n23302) | (n23293 & n31852) | (n23302 & n31852);
  assign n23643 = n23640 & ~n31853;
  assign n23644 = ~n23640 & n31853;
  assign n23645 = n23643 | n23644;
  assign n23646 = x115 & x172;
  assign n23647 = n23645 | n23646;
  assign n23648 = n23645 & n23646;
  assign n23649 = n23647 & ~n23648;
  assign n31854 = n23307 & n23308;
  assign n31855 = (n23307 & n23311) | (n23307 & n31854) | (n23311 & n31854);
  assign n23652 = n23649 & ~n31855;
  assign n23653 = ~n23649 & n31855;
  assign n23654 = n23652 | n23653;
  assign n23655 = x114 & x173;
  assign n23656 = n23654 | n23655;
  assign n23657 = n23654 & n23655;
  assign n23658 = n23656 & ~n23657;
  assign n23659 = n22981 | n23317;
  assign n23660 = n23316 & n23659;
  assign n23661 = n23658 & ~n23660;
  assign n23662 = ~n23658 & n23660;
  assign n23663 = n23661 | n23662;
  assign n23664 = x113 & x174;
  assign n23665 = n23663 | n23664;
  assign n23666 = n23663 & n23664;
  assign n23667 = n23665 & ~n23666;
  assign n23668 = ~n23323 & n23667;
  assign n23669 = n23323 & ~n23667;
  assign n23670 = n23668 | n23669;
  assign n23671 = x112 & x175;
  assign n23672 = n23670 & n23671;
  assign n23673 = n23670 | n23671;
  assign n23674 = ~n23672 & n23673;
  assign n23675 = n23323 | n23666;
  assign n23676 = n23665 & n23675;
  assign n23677 = x114 & x174;
  assign n31856 = n23656 & n23657;
  assign n31857 = (n23656 & n23660) | (n23656 & n31856) | (n23660 & n31856);
  assign n23680 = x116 & x172;
  assign n23681 = ~n31697 & n23637;
  assign n23682 = n31697 & ~n23637;
  assign n23683 = n23681 | n23682;
  assign n23686 = n23328 | n23683;
  assign n23684 = n23328 & n23683;
  assign n31858 = n23684 & n23686;
  assign n31859 = (n23686 & n31853) | (n23686 & n31858) | (n31853 & n31858);
  assign n31860 = n23635 & n23636;
  assign n31861 = (n23635 & n31697) | (n23635 & n31860) | (n31697 & n31860);
  assign n23690 = x118 & x170;
  assign n31862 = n23629 & n23630;
  assign n31863 = (n23630 & n31699) | (n23630 & n31862) | (n31699 & n31862);
  assign n31864 = n23623 & n23624;
  assign n31865 = (n23623 & n31701) | (n23623 & n31864) | (n31701 & n31864);
  assign n31866 = n23614 & n23615;
  assign n31867 = (n23614 & n31851) | (n23614 & n31866) | (n31851 & n31866);
  assign n23697 = x121 & x167;
  assign n23698 = x120 & x168;
  assign n23699 = n23697 & n23698;
  assign n23700 = n23697 | n23698;
  assign n23701 = ~n23699 & n23700;
  assign n31868 = n23605 & n23606;
  assign n31869 = (n23605 & n31849) | (n23605 & n31868) | (n31849 & n31868);
  assign n23704 = x122 & x166;
  assign n23707 = n23584 | n31843;
  assign n31870 = ~n23584 & n23585;
  assign n31871 = (n23585 & ~n31843) | (n23585 & n31870) | (~n31843 & n31870);
  assign n23710 = n23707 & n31871;
  assign n31872 = n23595 | n23710;
  assign n31873 = (n23710 & n31707) | (n23710 & n31872) | (n31707 & n31872);
  assign n23712 = n23572 & n23581;
  assign n23713 = n23572 | n23581;
  assign n23714 = ~n23712 & n23713;
  assign n23715 = n23573 & n23714;
  assign n31874 = n23584 | n23715;
  assign n31875 = (n23715 & n31843) | (n23715 & n31874) | (n31843 & n31874);
  assign n23717 = n23361 | n23565;
  assign n23719 = n23004 | n23359;
  assign n23720 = n23565 & n23719;
  assign n31876 = n23002 | n23360;
  assign n31877 = n31520 | n31876;
  assign n31878 = n23566 & ~n31877;
  assign n31879 = (n23566 & ~n23720) | (n23566 & n31878) | (~n23720 & n31878);
  assign n23723 = n23717 & n31879;
  assign n31880 = n23572 | n23723;
  assign n31881 = (n23581 & n23723) | (n23581 & n31880) | (n23723 & n31880);
  assign n23729 = n23540 & n31829;
  assign n31886 = (n23541 & n23543) | (n23541 & n31829) | (n23543 & n31829);
  assign n23732 = ~n23729 & n31886;
  assign n31882 = n23013 | n31724;
  assign n31883 = n31526 | n31882;
  assign n31884 = n23189 | n31722;
  assign n31885 = (n23189 & ~n23370) | (n23189 & n31884) | (~n23370 & n31884);
  assign n23727 = n23551 & n31885;
  assign n31887 = n23727 | n23732;
  assign n31888 = (n23732 & n31883) | (n23732 & n31887) | (n31883 & n31887);
  assign n31889 = n23389 & n23527;
  assign n31890 = (n23527 & n31731) | (n23527 & n31889) | (n31731 & n31889);
  assign n35798 = n23389 & n23528;
  assign n35799 = (n23527 & n23528) | (n23527 & n35798) | (n23528 & n35798);
  assign n31894 = (n23528 & n31731) | (n23528 & n35799) | (n31731 & n35799);
  assign n23737 = ~n31890 & n31894;
  assign n35800 = n23026 | n23175;
  assign n35801 = (n23026 & n23382) | (n23026 & n35800) | (n23382 & n35800);
  assign n35802 = n23018 | n35801;
  assign n35803 = (n23016 & n35801) | (n23016 & n35802) | (n35801 & n35802);
  assign n23740 = n23175 | n23382;
  assign n23741 = n23534 & n23740;
  assign n31895 = n23737 | n23741;
  assign n31896 = (n23737 & n35803) | (n23737 & n31895) | (n35803 & n31895);
  assign n31897 = n23520 | n31741;
  assign n31898 = n23520 | n31740;
  assign n31899 = (n31555 & n31897) | (n31555 & n31898) | (n31897 & n31898);
  assign n31900 = ~n23161 & n31738;
  assign n31901 = (n23161 & n35702) | (n23161 & ~n31900) | (n35702 & ~n31900);
  assign n23747 = n23520 & n31901;
  assign n31902 = n23747 & n31740;
  assign n31903 = (n23747 & n31555) | (n23747 & n31902) | (n31555 & n31902);
  assign n23749 = n31899 & ~n31903;
  assign n23750 = n23521 & n23749;
  assign n31904 = n23750 | n31889;
  assign n31905 = n23527 | n23750;
  assign n31906 = (n31731 & n31904) | (n31731 & n31905) | (n31904 & n31905);
  assign n23753 = n35712 | n23506;
  assign n31909 = n23753 | n31743;
  assign n31910 = n23149 | n23753;
  assign n31911 = (n31562 & n31909) | (n31562 & n31910) | (n31909 & n31910);
  assign n35804 = n23143 | n35710;
  assign n35805 = (n23143 & ~n23407) | (n23143 & n35804) | (~n23407 & n35804);
  assign n23757 = n23506 & n35805;
  assign n31912 = n23156 | n35712;
  assign n31914 = n23757 & n31912;
  assign n31915 = (n23757 & n31562) | (n23757 & n31914) | (n31562 & n31914);
  assign n23759 = n31911 & ~n31915;
  assign n23760 = n23507 & n23759;
  assign n31907 = n23402 & n23513;
  assign n31916 = n23760 | n31907;
  assign n31917 = n23513 | n23760;
  assign n31918 = (n31738 & n31916) | (n31738 & n31917) | (n31916 & n31917);
  assign n31920 = n23415 & n23499;
  assign n35806 = (n23406 & n23499) | (n23406 & n31920) | (n23499 & n31920);
  assign n31921 = (n31751 & n35806) | (n31751 & n31920) | (n35806 & n31920);
  assign n31923 = n23415 | n23499;
  assign n35807 = n23406 | n31923;
  assign n35808 = n23500 & n35807;
  assign n37475 = n23415 & n23500;
  assign n37476 = (n23499 & n23500) | (n23499 & n37475) | (n23500 & n37475);
  assign n35810 = (n31751 & n35808) | (n31751 & n37476) | (n35808 & n37476);
  assign n23765 = ~n31921 & n35810;
  assign n23767 = n23425 | n23492;
  assign n31925 = n23767 | n31757;
  assign n35811 = n23135 | n23492;
  assign n35812 = n23425 | n35811;
  assign n31927 = (n31572 & n31925) | (n31572 & n35812) | (n31925 & n35812);
  assign n23771 = n23129 | n23424;
  assign n23772 = n23492 & n23771;
  assign n23769 = n23062 | n23425;
  assign n31928 = n23769 & n23772;
  assign n31929 = (n23772 & n31572) | (n23772 & n31928) | (n31572 & n31928);
  assign n23774 = n31927 & ~n31929;
  assign n23775 = n23493 & n23774;
  assign n35813 = n23775 | n35806;
  assign n35814 = n23775 | n31920;
  assign n35815 = (n31751 & n35813) | (n31751 & n35814) | (n35813 & n35814);
  assign n35816 = n23485 & n35735;
  assign n35817 = n23485 & n35737;
  assign n35818 = (n35571 & n35816) | (n35571 & n35817) | (n35816 & n35817);
  assign n35819 = (n23486 & n23488) | (n23486 & n35735) | (n23488 & n35735);
  assign n35820 = (n23486 & n23488) | (n23486 & n35737) | (n23488 & n35737);
  assign n35821 = (n35571 & n35819) | (n35571 & n35820) | (n35819 & n35820);
  assign n23780 = ~n35818 & n35821;
  assign n31783 = (n35571 & n35735) | (n35571 & n35737) | (n35735 & n35737);
  assign n23798 = x140 & x148;
  assign n23804 = x141 & x147;
  assign n23808 = x143 & x145;
  assign n23806 = n23444 & n23445;
  assign n31950 = n23806 & n23808;
  assign n37855 = (n23448 & n23808) | (n23448 & n31950) | (n23808 & n31950);
  assign n37857 = (n37462 & n37855) | (n37462 & n31950) | (n37855 & n31950);
  assign n37752 = (n23808 & n31950) | (n23808 & n37466) | (n31950 & n37466);
  assign n37753 = (n35586 & n37857) | (n35586 & n37752) | (n37857 & n37752);
  assign n35823 = (n23808 & n31950) | (n23808 & n37468) | (n31950 & n37468);
  assign n35824 = (n35438 & n37753) | (n35438 & n35823) | (n37753 & n35823);
  assign n31952 = n23806 | n23808;
  assign n37858 = n23448 | n31952;
  assign n37859 = (n31952 & n37462) | (n31952 & n37858) | (n37462 & n37858);
  assign n37755 = n31952 | n37466;
  assign n37756 = (n35586 & n37859) | (n35586 & n37755) | (n37859 & n37755);
  assign n35826 = n31952 | n37468;
  assign n35827 = (n35438 & n37756) | (n35438 & n35826) | (n37756 & n35826);
  assign n23811 = ~n35824 & n35827;
  assign n23812 = x142 & x146;
  assign n23813 = n23811 & n23812;
  assign n23814 = n23811 | n23812;
  assign n23815 = ~n23813 & n23814;
  assign n31948 = n23452 | n23454;
  assign n31954 = n23815 & n31948;
  assign n31955 = n23452 & n23815;
  assign n31956 = (n35743 & n31954) | (n35743 & n31955) | (n31954 & n31955);
  assign n31957 = n23815 | n31948;
  assign n31958 = n23452 | n23815;
  assign n31959 = (n35743 & n31957) | (n35743 & n31958) | (n31957 & n31958);
  assign n23818 = ~n31956 & n31959;
  assign n23819 = n23804 & n23818;
  assign n23820 = n23804 | n23818;
  assign n23821 = ~n23819 & n23820;
  assign n23799 = n35743 & n23454;
  assign n31946 = n23441 & n23454;
  assign n31947 = (n23441 & n35743) | (n23441 & n31946) | (n35743 & n31946);
  assign n23802 = ~n23799 & n31947;
  assign n31960 = n23802 & n23821;
  assign n35828 = (n23821 & n31815) | (n23821 & n31960) | (n31815 & n31960);
  assign n35829 = (n23821 & n31816) | (n23821 & n31960) | (n31816 & n31960);
  assign n35830 = (n35600 & n35828) | (n35600 & n35829) | (n35828 & n35829);
  assign n31962 = n23802 | n23821;
  assign n35831 = n31815 | n31962;
  assign n35832 = n31816 | n31962;
  assign n35833 = (n35600 & n35831) | (n35600 & n35832) | (n35831 & n35832);
  assign n23824 = ~n35830 & n35833;
  assign n23825 = n23798 | n23824;
  assign n23826 = n23798 & n23824;
  assign n23827 = n23825 & ~n23826;
  assign n23828 = x139 & x149;
  assign n23829 = n23827 & n23828;
  assign n23830 = n23827 | n23828;
  assign n23831 = ~n23829 & n23830;
  assign n31944 = n23468 & n23469;
  assign n31964 = n23831 & n31944;
  assign n31965 = n23469 & n23831;
  assign n31966 = (n35760 & n31964) | (n35760 & n31965) | (n31964 & n31965);
  assign n31967 = n23831 | n31944;
  assign n31968 = n23469 | n23831;
  assign n31969 = (n35760 & n31967) | (n35760 & n31968) | (n31967 & n31968);
  assign n23834 = ~n31966 & n31969;
  assign n23835 = x138 & x150;
  assign n23836 = n23834 | n23835;
  assign n23837 = n23834 & n23835;
  assign n23838 = n23836 & ~n23837;
  assign n23791 = n23470 & n35760;
  assign n31940 = (n23471 & n23472) | (n23471 & n35760) | (n23472 & n35760);
  assign n23794 = ~n23791 & n31940;
  assign n23783 = n23115 | n23436;
  assign n23784 = n23478 & n23783;
  assign n31931 = n23077 | n23437;
  assign n31933 = n23784 & n31931;
  assign n31941 = n23794 | n31933;
  assign n35834 = n23838 | n31941;
  assign n31942 = n23784 | n23794;
  assign n35835 = n23838 | n31942;
  assign n35836 = (n31588 & n35834) | (n31588 & n35835) | (n35834 & n35835);
  assign n35837 = n23838 & n31941;
  assign n35838 = n23838 & n31942;
  assign n35839 = (n31588 & n35837) | (n31588 & n35838) | (n35837 & n35838);
  assign n23841 = n35836 & ~n35839;
  assign n23842 = x137 & x151;
  assign n23843 = n23841 | n23842;
  assign n23844 = n23841 & n23842;
  assign n23845 = n23843 & ~n23844;
  assign n35840 = (n23784 & n31587) | (n23784 & n31933) | (n31587 & n31933);
  assign n35841 = (n23784 & n31586) | (n23784 & n31933) | (n31586 & n31933);
  assign n35842 = (n31244 & n35840) | (n31244 & n35841) | (n35840 & n35841);
  assign n23786 = n23437 | n23478;
  assign n31935 = n23786 | n31775;
  assign n31936 = n23121 | n23786;
  assign n35843 = (n31587 & n31935) | (n31587 & n31936) | (n31935 & n31936);
  assign n35844 = (n31586 & n31935) | (n31586 & n31936) | (n31935 & n31936);
  assign n35845 = (n31244 & n35843) | (n31244 & n35844) | (n35843 & n35844);
  assign n23788 = ~n35842 & n35845;
  assign n23789 = n23479 & n23788;
  assign n31938 = n23485 | n23789;
  assign n31970 = n23845 & ~n31938;
  assign n31971 = ~n23789 & n23845;
  assign n31972 = (~n31783 & n31970) | (~n31783 & n31971) | (n31970 & n31971);
  assign n31973 = ~n23845 & n31938;
  assign n31974 = n23789 & ~n23845;
  assign n31975 = (n31783 & n31973) | (n31783 & n31974) | (n31973 & n31974);
  assign n23848 = n31972 | n31975;
  assign n23849 = x136 & x152;
  assign n23850 = n23848 | n23849;
  assign n23851 = n23848 & n23849;
  assign n23852 = n23850 & ~n23851;
  assign n31976 = ~n23780 & n23852;
  assign n31977 = ~n31929 & n31976;
  assign n31978 = n23780 & ~n23852;
  assign n31979 = (~n23852 & n31929) | (~n23852 & n31978) | (n31929 & n31978);
  assign n23855 = n31977 | n31979;
  assign n23856 = x135 & x153;
  assign n23857 = n23855 & n23856;
  assign n23858 = n23855 | n23856;
  assign n23859 = ~n23857 & n23858;
  assign n23860 = x134 & x154;
  assign n23861 = n23859 & ~n23860;
  assign n23862 = ~n23859 & n23860;
  assign n23863 = n23861 | n23862;
  assign n23864 = n35815 | n23863;
  assign n23865 = n35815 & n23863;
  assign n23866 = n23864 & ~n23865;
  assign n31980 = ~n23765 & n23866;
  assign n31981 = ~n31915 & n31980;
  assign n31982 = n23765 & ~n23866;
  assign n31983 = (~n23866 & n31915) | (~n23866 & n31982) | (n31915 & n31982);
  assign n23869 = n31981 | n31983;
  assign n23870 = x133 & x155;
  assign n23871 = n23869 & n23870;
  assign n23872 = n23869 | n23870;
  assign n23873 = ~n23871 & n23872;
  assign n23874 = n31918 | n23873;
  assign n23875 = n31918 & n23873;
  assign n23876 = n23874 & ~n23875;
  assign n23877 = x132 & x156;
  assign n23878 = n23876 | n23877;
  assign n23879 = n23876 & n23877;
  assign n23880 = n23878 & ~n23879;
  assign n31984 = n23402 | n23513;
  assign n31985 = n31738 | n31984;
  assign n31986 = n23514 & ~n31907;
  assign n31987 = ~n23513 & n23514;
  assign n31988 = (~n31738 & n31986) | (~n31738 & n31987) | (n31986 & n31987);
  assign n23883 = n31985 & n31988;
  assign n31989 = ~n23880 & n23883;
  assign n31990 = (~n23880 & n31903) | (~n23880 & n31989) | (n31903 & n31989);
  assign n31991 = n23880 & ~n23883;
  assign n31992 = ~n31903 & n31991;
  assign n23887 = n31990 | n31992;
  assign n23888 = x131 & x157;
  assign n23889 = n23887 & n23888;
  assign n23890 = n23887 | n23888;
  assign n23891 = ~n23889 & n23890;
  assign n23892 = n31906 | n23891;
  assign n23893 = n31906 & n23891;
  assign n23894 = n23892 & ~n23893;
  assign n23895 = x130 & x158;
  assign n23896 = n23894 | n23895;
  assign n23897 = n23894 & n23895;
  assign n23898 = n23896 & ~n23897;
  assign n23899 = ~n31896 & n23898;
  assign n23900 = n31896 & ~n23898;
  assign n23901 = n23899 | n23900;
  assign n23742 = n35803 & n23741;
  assign n31993 = n23534 | n31732;
  assign n31994 = n23383 | n23534;
  assign n31995 = (n31540 & n31993) | (n31540 & n31994) | (n31993 & n31994);
  assign n31996 = n23385 & n31995;
  assign n31997 = ~n23742 & n31996;
  assign n23905 = n23901 | n31997;
  assign n35846 = n23540 | n23905;
  assign n35847 = (n23905 & n31829) | (n23905 & n35846) | (n31829 & n35846);
  assign n31998 = n23385 | n31995;
  assign n31999 = (n23385 & ~n23742) | (n23385 & n31998) | (~n23742 & n31998);
  assign n23909 = n23901 & n31999;
  assign n35848 = n23909 & n31997;
  assign n35849 = (n23909 & n31829) | (n23909 & n35848) | (n31829 & n35848);
  assign n23911 = n35847 & ~n35849;
  assign n23912 = x129 & x159;
  assign n23913 = n23911 & n23912;
  assign n23914 = n23911 | n23912;
  assign n23915 = ~n23913 & n23914;
  assign n23916 = n31888 & n23915;
  assign n23917 = n31888 | n23915;
  assign n23918 = ~n23916 & n23917;
  assign n23919 = x128 & x160;
  assign n23920 = n23918 & n23919;
  assign n23921 = n23918 | n23919;
  assign n23922 = ~n23920 & n23921;
  assign n23728 = n31883 & n23727;
  assign n23923 = n31727 | n23551;
  assign n23924 = ~n23728 & n23923;
  assign n23925 = n23552 & n23924;
  assign n32000 = n23925 | n31830;
  assign n32001 = n23558 | n23925;
  assign n32002 = (n23358 & n32000) | (n23358 & n32001) | (n32000 & n32001);
  assign n23927 = n23922 | n32002;
  assign n23928 = n23922 & n32002;
  assign n23929 = n23927 & ~n23928;
  assign n23930 = x127 & x161;
  assign n23931 = n23929 & ~n23930;
  assign n23932 = ~n23929 & n23930;
  assign n23933 = n23931 | n23932;
  assign n23934 = x126 & x162;
  assign n23935 = n23933 & n23934;
  assign n23936 = n23933 | n23934;
  assign n23937 = ~n23935 & n23936;
  assign n32003 = n23563 | n31877;
  assign n32004 = (n23563 & n23720) | (n23563 & n32003) | (n23720 & n32003);
  assign n23939 = n23937 | n32004;
  assign n23940 = n23937 & n32004;
  assign n23941 = n23939 & ~n23940;
  assign n23942 = x125 & x163;
  assign n23943 = n23941 | n23942;
  assign n23944 = n23941 & n23942;
  assign n23945 = n23943 & ~n23944;
  assign n23946 = n31881 | n23945;
  assign n23947 = n31881 & n23945;
  assign n23948 = n23946 & ~n23947;
  assign n23949 = x124 & x164;
  assign n23950 = n23948 | n23949;
  assign n23951 = n23948 & n23949;
  assign n23952 = n23950 & ~n23951;
  assign n23953 = n31875 | n23952;
  assign n23954 = n31875 & n23952;
  assign n23955 = n23953 & ~n23954;
  assign n23956 = ~n31873 & n23955;
  assign n23957 = n31873 & ~n23955;
  assign n23958 = n23956 | n23957;
  assign n23959 = x123 & x165;
  assign n23960 = n23958 & n23959;
  assign n23961 = n23958 | n23959;
  assign n23962 = ~n23960 & n23961;
  assign n23705 = n23345 & n23598;
  assign n32005 = n23705 & n23962;
  assign n32006 = (n23962 & n31845) | (n23962 & n32005) | (n31845 & n32005);
  assign n32007 = n23705 | n23962;
  assign n32008 = n31845 | n32007;
  assign n23965 = ~n32006 & n32008;
  assign n23966 = n23704 & n23965;
  assign n23967 = n23704 | n23965;
  assign n23968 = ~n23966 & n23967;
  assign n23969 = n31869 & n23968;
  assign n23970 = n31869 | n23968;
  assign n23971 = ~n23969 & n23970;
  assign n23972 = n23701 & n23971;
  assign n23973 = n23701 | n23971;
  assign n23974 = ~n23972 & n23973;
  assign n23975 = n31867 & n23974;
  assign n23976 = n31867 | n23974;
  assign n23977 = ~n23975 & n23976;
  assign n23978 = n31865 & ~n23977;
  assign n23979 = ~n31865 & n23977;
  assign n23980 = n23978 | n23979;
  assign n23981 = x119 & x169;
  assign n23982 = n23980 & n23981;
  assign n23983 = n23980 | n23981;
  assign n23984 = ~n23982 & n23983;
  assign n23985 = n31863 | n23984;
  assign n23986 = n31863 & n23984;
  assign n23987 = n23985 & ~n23986;
  assign n23988 = n23690 & n23987;
  assign n23989 = n23690 | n23987;
  assign n23990 = ~n23988 & n23989;
  assign n23991 = n31861 & ~n23990;
  assign n23992 = ~n31861 & n23990;
  assign n23993 = n23991 | n23992;
  assign n23994 = x117 & x171;
  assign n23995 = n23993 & n23994;
  assign n23996 = n23993 | n23994;
  assign n23997 = ~n23995 & n23996;
  assign n23998 = n31859 & n23997;
  assign n23999 = n31859 | n23997;
  assign n24000 = ~n23998 & n23999;
  assign n24001 = n23680 | n24000;
  assign n24002 = n23680 & n24000;
  assign n24003 = n24001 & ~n24002;
  assign n32009 = n23647 & n23648;
  assign n32010 = (n23647 & n31855) | (n23647 & n32009) | (n31855 & n32009);
  assign n24006 = n24003 & ~n32010;
  assign n24007 = ~n24003 & n32010;
  assign n24008 = n24006 | n24007;
  assign n24009 = x115 & x173;
  assign n24010 = n24008 & n24009;
  assign n24011 = n24008 | n24009;
  assign n24012 = ~n24010 & n24011;
  assign n24013 = n31857 & n24012;
  assign n24014 = n31857 | n24012;
  assign n24015 = ~n24013 & n24014;
  assign n24016 = n23677 & n24015;
  assign n24017 = n23677 | n24015;
  assign n24018 = ~n24016 & n24017;
  assign n24019 = ~n23676 & n24018;
  assign n24020 = n23676 & ~n24018;
  assign n24021 = n24019 | n24020;
  assign n24022 = x113 & x175;
  assign n24023 = n24021 | n24022;
  assign n24024 = n24021 & n24022;
  assign n24025 = n24023 & ~n24024;
  assign n24026 = ~n23672 & n24025;
  assign n24027 = n23672 & ~n24025;
  assign n24028 = n24026 | n24027;
  assign n24029 = x114 & x175;
  assign n24030 = n23676 & n24018;
  assign n24031 = n24016 | n24030;
  assign n24032 = x115 & x174;
  assign n24033 = n24010 | n24013;
  assign n24034 = x117 & x172;
  assign n24035 = n23995 | n23998;
  assign n24036 = x118 & x171;
  assign n24037 = n31861 & n23990;
  assign n24038 = n23988 | n24037;
  assign n24039 = x119 & x170;
  assign n24040 = n23982 | n23986;
  assign n24042 = n23697 & n23968;
  assign n24043 = n23697 | n23968;
  assign n24044 = ~n24042 & n24043;
  assign n24045 = n31869 | n24044;
  assign n24046 = n31869 & n24044;
  assign n24047 = n24045 & ~n24046;
  assign n24048 = n31867 & n24047;
  assign n24049 = n31867 | n24047;
  assign n24050 = n23698 & n24049;
  assign n24051 = ~n24048 & n24050;
  assign n32011 = n23977 | n24051;
  assign n32012 = (n24051 & n31865) | (n24051 & n32011) | (n31865 & n32011);
  assign n24053 = n23697 & n23971;
  assign n24054 = n24048 | n24053;
  assign n24055 = x122 & x167;
  assign n24056 = x121 & x168;
  assign n24057 = n24055 & n24056;
  assign n24058 = n24055 | n24056;
  assign n24059 = ~n24057 & n24058;
  assign n24060 = n23966 | n23969;
  assign n24061 = x123 & x166;
  assign n24062 = n23960 | n32006;
  assign n24064 = n31875 | n23948;
  assign n24065 = n31843 | n23715;
  assign n24066 = n23573 | n23714;
  assign n24067 = n23948 & n24066;
  assign n24068 = n24065 & n24067;
  assign n24069 = n23949 & ~n24068;
  assign n24070 = n24064 & n24069;
  assign n32013 = n23955 | n24070;
  assign n32014 = (n24070 & n31873) | (n24070 & n32013) | (n31873 & n32013);
  assign n24072 = x125 & x164;
  assign n24074 = n23933 & n32004;
  assign n32015 = (n23934 & n23935) | (n23934 & n32004) | (n23935 & n32004);
  assign n24077 = ~n24074 & n32015;
  assign n32016 = n23941 | n24077;
  assign n32017 = (n24077 & n31881) | (n24077 & n32016) | (n31881 & n32016);
  assign n35850 = n23365 | n23552;
  assign n35851 = (n23365 & n23924) | (n23365 & n35850) | (n23924 & n35850);
  assign n32019 = n23358 | n35851;
  assign n24080 = n23552 | n23924;
  assign n24081 = ~n23912 & n23919;
  assign n24082 = n23912 & ~n23919;
  assign n24083 = n24081 | n24082;
  assign n24084 = n23911 & ~n24083;
  assign n24085 = ~n23911 & n24083;
  assign n24086 = n24084 | n24085;
  assign n24087 = n31888 & n24086;
  assign n24088 = n31888 | n24086;
  assign n24089 = ~n24087 & n24088;
  assign n24090 = n24080 & n24089;
  assign n24091 = n32019 & n24090;
  assign n24092 = n23927 & ~n24091;
  assign n24093 = n23930 & n24092;
  assign n24094 = n32004 | n24093;
  assign n24095 = n23930 | n24092;
  assign n24096 = x128 & x161;
  assign n24099 = n23521 | n23749;
  assign n24100 = n23887 & n24099;
  assign n35852 = n23389 | n23521;
  assign n35853 = (n23389 & n23749) | (n23389 & n35852) | (n23749 & n35852);
  assign n32022 = n24100 & n35853;
  assign n32023 = (n24100 & n31731) | (n24100 & n32022) | (n31731 & n32022);
  assign n32028 = n23876 & n23883;
  assign n35854 = (n23876 & n31902) | (n23876 & n32028) | (n31902 & n32028);
  assign n35855 = (n23747 & n23876) | (n23747 & n32028) | (n23876 & n32028);
  assign n35856 = (n31555 & n35854) | (n31555 & n35855) | (n35854 & n35855);
  assign n35857 = n23877 & n23883;
  assign n35858 = (n23876 & n23877) | (n23876 & n35857) | (n23877 & n35857);
  assign n35859 = (n23877 & n31902) | (n23877 & n35858) | (n31902 & n35858);
  assign n35860 = (n23747 & n23877) | (n23747 & n35858) | (n23877 & n35858);
  assign n35861 = (n31555 & n35859) | (n31555 & n35860) | (n35859 & n35860);
  assign n24109 = ~n35856 & n35861;
  assign n24115 = n23507 | n23759;
  assign n24116 = n23869 & n24115;
  assign n24113 = n23402 | n23760;
  assign n32037 = n24113 & n24116;
  assign n32038 = (n24116 & n31738) | (n24116 & n32037) | (n31738 & n32037);
  assign n32042 = n23775 | n23859;
  assign n32043 = n31921 | n32042;
  assign n32044 = n23775 & n23859;
  assign n32045 = (n23859 & n31921) | (n23859 & n32044) | (n31921 & n32044);
  assign n24123 = n32043 & ~n32045;
  assign n32046 = n23765 & n24123;
  assign n35862 = (n24123 & n31914) | (n24123 & n32046) | (n31914 & n32046);
  assign n35863 = (n23757 & n24123) | (n23757 & n32046) | (n24123 & n32046);
  assign n35864 = (n31562 & n35862) | (n31562 & n35863) | (n35862 & n35863);
  assign n35865 = n23765 & n23860;
  assign n35866 = (n23860 & n24123) | (n23860 & n35865) | (n24123 & n35865);
  assign n35867 = (n23860 & n31914) | (n23860 & n35866) | (n31914 & n35866);
  assign n35868 = (n23757 & n23860) | (n23757 & n35866) | (n23860 & n35866);
  assign n35869 = (n31562 & n35867) | (n31562 & n35868) | (n35867 & n35868);
  assign n24127 = ~n35864 & n35869;
  assign n24129 = n23775 | n23855;
  assign n35870 = n24129 | n35806;
  assign n35871 = n24129 | n31920;
  assign n35872 = (n31751 & n35870) | (n31751 & n35871) | (n35870 & n35871);
  assign n35873 = n23415 | n23493;
  assign n35874 = (n23415 & n23774) | (n23415 & n35873) | (n23774 & n35873);
  assign n32052 = n23406 | n35874;
  assign n32053 = (n35874 & n31751) | (n35874 & n32052) | (n31751 & n32052);
  assign n24133 = n23493 | n23774;
  assign n24134 = n23855 & n24133;
  assign n32054 = n23856 & ~n24134;
  assign n32055 = (n23856 & ~n32053) | (n23856 & n32054) | (~n32053 & n32054);
  assign n24137 = n35872 & n32055;
  assign n32056 = n24137 | n32046;
  assign n32057 = n24123 | n24137;
  assign n32058 = (n31915 & n32056) | (n31915 & n32057) | (n32056 & n32057);
  assign n24146 = n23430 | n23789;
  assign n32069 = n24146 | n31770;
  assign n32070 = n23422 | n24146;
  assign n32071 = (n35571 & n32069) | (n35571 & n32070) | (n32069 & n32070);
  assign n24162 = x141 & x148;
  assign n24164 = x142 & x147;
  assign n24166 = x143 & x146;
  assign n32095 = n23808 & ~n24166;
  assign n35875 = n23806 & n32095;
  assign n37860 = (n23448 & n32095) | (n23448 & n35875) | (n32095 & n35875);
  assign n37861 = n32095 & n35875;
  assign n37862 = (n37462 & n37860) | (n37462 & n37861) | (n37860 & n37861);
  assign n37758 = (n32095 & n35875) | (n32095 & n37466) | (n35875 & n37466);
  assign n37759 = (n35586 & n37862) | (n35586 & n37758) | (n37862 & n37758);
  assign n35877 = (n32095 & n37468) | (n32095 & n35875) | (n37468 & n35875);
  assign n35878 = (n35438 & n37759) | (n35438 & n35877) | (n37759 & n35877);
  assign n32098 = ~n23808 & n24166;
  assign n35879 = (~n23806 & n24166) | (~n23806 & n32098) | (n24166 & n32098);
  assign n37863 = (~n23448 & n32098) | (~n23448 & n35879) | (n32098 & n35879);
  assign n37864 = n32098 | n35879;
  assign n37865 = (~n37462 & n37863) | (~n37462 & n37864) | (n37863 & n37864);
  assign n37761 = (n32098 & n35879) | (n32098 & ~n37466) | (n35879 & ~n37466);
  assign n37762 = (~n35586 & n37865) | (~n35586 & n37761) | (n37865 & n37761);
  assign n35881 = (n32098 & ~n37468) | (n32098 & n35879) | (~n37468 & n35879);
  assign n35882 = (~n35438 & n37762) | (~n35438 & n35881) | (n37762 & n35881);
  assign n24169 = n35878 | n35882;
  assign n35883 = n23813 | n23815;
  assign n35884 = (n23813 & n31948) | (n23813 & n35883) | (n31948 & n35883);
  assign n32100 = n24169 & n35884;
  assign n35885 = n23452 | n23813;
  assign n35886 = (n23813 & n23815) | (n23813 & n35885) | (n23815 & n35885);
  assign n32101 = n24169 & n35886;
  assign n32102 = (n35743 & n32100) | (n35743 & n32101) | (n32100 & n32101);
  assign n32103 = n24169 | n35884;
  assign n32104 = n24169 | n35886;
  assign n32105 = (n35743 & n32103) | (n35743 & n32104) | (n32103 & n32104);
  assign n24172 = ~n32102 & n32105;
  assign n24173 = n24164 & n24172;
  assign n24174 = n24164 | n24172;
  assign n24175 = ~n24173 & n24174;
  assign n35887 = n23802 | n23819;
  assign n35888 = (n23819 & n23821) | (n23819 & n35887) | (n23821 & n35887);
  assign n32106 = n24175 & n35888;
  assign n32089 = n23819 | n23821;
  assign n32107 = n24175 & n32089;
  assign n35889 = (n31815 & n32106) | (n31815 & n32107) | (n32106 & n32107);
  assign n35890 = (n31816 & n32106) | (n31816 & n32107) | (n32106 & n32107);
  assign n35891 = (n35600 & n35889) | (n35600 & n35890) | (n35889 & n35890);
  assign n32109 = n24175 | n35888;
  assign n32110 = n24175 | n32089;
  assign n35892 = (n31815 & n32109) | (n31815 & n32110) | (n32109 & n32110);
  assign n35893 = (n31816 & n32109) | (n31816 & n32110) | (n32109 & n32110);
  assign n35894 = (n35600 & n35892) | (n35600 & n35893) | (n35892 & n35893);
  assign n24178 = ~n35891 & n35894;
  assign n24179 = n24162 & n24178;
  assign n24180 = n24162 | n24178;
  assign n24181 = ~n24179 & n24180;
  assign n24182 = x140 & x149;
  assign n24183 = n24181 & n24182;
  assign n24184 = n24181 | n24182;
  assign n24185 = ~n24183 & n24184;
  assign n32075 = n23827 & n31944;
  assign n32086 = n23826 | n32075;
  assign n32112 = n24185 | n32086;
  assign n35895 = n23469 | n23826;
  assign n35896 = (n23826 & n23827) | (n23826 & n35895) | (n23827 & n35895);
  assign n32113 = n24185 | n35896;
  assign n32114 = (n35760 & n32112) | (n35760 & n32113) | (n32112 & n32113);
  assign n32115 = n24185 & n32086;
  assign n32116 = n24185 & n35896;
  assign n32117 = (n35760 & n32115) | (n35760 & n32116) | (n32115 & n32116);
  assign n24188 = n32114 & ~n32117;
  assign n24189 = x139 & x150;
  assign n24190 = n24188 | n24189;
  assign n24191 = n24188 & n24189;
  assign n24192 = n24190 & ~n24191;
  assign n32076 = n23469 & n23827;
  assign n32077 = (n35760 & n32075) | (n35760 & n32076) | (n32075 & n32076);
  assign n24156 = n23468 | n23827;
  assign n35897 = n23470 & n23828;
  assign n35898 = (n23828 & n24156) | (n23828 & n35897) | (n24156 & n35897);
  assign n37477 = n23467 & n23828;
  assign n37478 = n23466 & n37477;
  assign n35900 = (n23827 & n23828) | (n23827 & n37478) | (n23828 & n37478);
  assign n32082 = (n35760 & n35898) | (n35760 & n35900) | (n35898 & n35900);
  assign n24159 = ~n32077 & n32082;
  assign n32083 = n23834 | n24159;
  assign n32118 = n24192 | n32083;
  assign n32119 = n24159 | n24192;
  assign n35901 = (n31941 & n32118) | (n31941 & n32119) | (n32118 & n32119);
  assign n35902 = (n31942 & n32118) | (n31942 & n32119) | (n32118 & n32119);
  assign n35903 = (n31588 & n35901) | (n31588 & n35902) | (n35901 & n35902);
  assign n32121 = n24192 & n32083;
  assign n32122 = n24159 & n24192;
  assign n35904 = (n31941 & n32121) | (n31941 & n32122) | (n32121 & n32122);
  assign n35905 = (n31942 & n32121) | (n31942 & n32122) | (n32121 & n32122);
  assign n35906 = (n31588 & n35904) | (n31588 & n35905) | (n35904 & n35905);
  assign n24195 = n35903 & ~n35906;
  assign n24196 = x138 & x151;
  assign n24197 = n24195 | n24196;
  assign n24198 = n24195 & n24196;
  assign n24199 = n24197 & ~n24198;
  assign n24148 = n23479 | n23788;
  assign n24149 = n23841 & n24148;
  assign n37479 = n23794 | n23834;
  assign n37480 = n31933 | n37479;
  assign n37481 = n23784 | n37479;
  assign n35909 = (n31588 & n37480) | (n31588 & n37481) | (n37480 & n37481);
  assign n32124 = ~n23834 & n23835;
  assign n37482 = (~n23794 & n23835) | (~n23794 & n32124) | (n23835 & n32124);
  assign n37484 = (~n31933 & n37482) | (~n31933 & n32124) | (n37482 & n32124);
  assign n35911 = (n23835 & ~n31942) | (n23835 & n32124) | (~n31942 & n32124);
  assign n35912 = (~n31588 & n37484) | (~n31588 & n35911) | (n37484 & n35911);
  assign n24202 = n35909 & n35912;
  assign n32126 = n24149 | n24202;
  assign n32128 = ~n24199 & n32126;
  assign n32129 = ~n24199 & n24202;
  assign n32130 = (n32071 & n32128) | (n32071 & n32129) | (n32128 & n32129);
  assign n32131 = n24199 & ~n32126;
  assign n32132 = n24199 & ~n24202;
  assign n32133 = (~n32071 & n32131) | (~n32071 & n32132) | (n32131 & n32132);
  assign n24206 = n32130 | n32133;
  assign n24207 = x137 & x152;
  assign n24208 = n24206 & n24207;
  assign n24209 = n24206 | n24207;
  assign n24210 = ~n24208 & n24209;
  assign n24150 = n32071 & n24149;
  assign n24144 = n23789 | n23841;
  assign n32067 = n23485 | n24144;
  assign n35913 = (n24144 & n32067) | (n24144 & n35735) | (n32067 & n35735);
  assign n35914 = (n24144 & n32067) | (n24144 & n35737) | (n32067 & n35737);
  assign n35915 = (n35571 & n35913) | (n35571 & n35914) | (n35913 & n35914);
  assign n35916 = n23842 & n35915;
  assign n35917 = ~n24150 & n35916;
  assign n32073 = n23848 | n35917;
  assign n32134 = n24210 & ~n32073;
  assign n32059 = n23780 & n23848;
  assign n32072 = n35917 | n32059;
  assign n32135 = n24210 & ~n32072;
  assign n32136 = (~n31929 & n32134) | (~n31929 & n32135) | (n32134 & n32135);
  assign n32137 = ~n24210 & n32073;
  assign n32138 = ~n24210 & n32072;
  assign n32139 = (n31929 & n32137) | (n31929 & n32138) | (n32137 & n32138);
  assign n24213 = n32136 | n32139;
  assign n24214 = x136 & x153;
  assign n24215 = n24213 | n24214;
  assign n24216 = n24213 & n24214;
  assign n24217 = n24215 & ~n24216;
  assign n35918 = (n23848 & n31928) | (n23848 & n32059) | (n31928 & n32059);
  assign n35919 = (n23772 & n23848) | (n23772 & n32059) | (n23848 & n32059);
  assign n35920 = (n31572 & n35918) | (n31572 & n35919) | (n35918 & n35919);
  assign n35921 = n23780 & n23849;
  assign n35922 = (n23848 & n23849) | (n23848 & n35921) | (n23849 & n35921);
  assign n35923 = (n23849 & n31928) | (n23849 & n35922) | (n31928 & n35922);
  assign n35924 = (n23772 & n23849) | (n23772 & n35922) | (n23849 & n35922);
  assign n35925 = (n31572 & n35923) | (n31572 & n35924) | (n35923 & n35924);
  assign n24142 = ~n35920 & n35925;
  assign n32065 = n24134 | n24142;
  assign n32140 = n24217 & ~n32065;
  assign n32141 = ~n24142 & n24217;
  assign n32142 = (~n32053 & n32140) | (~n32053 & n32141) | (n32140 & n32141);
  assign n32143 = ~n24217 & n32065;
  assign n32144 = n24142 & ~n24217;
  assign n32145 = (n32053 & n32143) | (n32053 & n32144) | (n32143 & n32144);
  assign n24220 = n32142 | n32145;
  assign n24221 = x135 & x154;
  assign n24222 = n24220 & n24221;
  assign n24223 = n24220 | n24221;
  assign n24224 = ~n24222 & n24223;
  assign n24225 = x134 & x155;
  assign n24226 = n24224 & ~n24225;
  assign n24227 = ~n24224 & n24225;
  assign n24228 = n24226 | n24227;
  assign n24229 = n32058 | n24228;
  assign n24230 = n32058 & n24228;
  assign n24231 = n24229 & ~n24230;
  assign n32146 = ~n24127 & n24231;
  assign n32147 = ~n32038 & n32146;
  assign n32148 = n24127 & ~n24231;
  assign n32149 = (~n24231 & n32038) | (~n24231 & n32148) | (n32038 & n32148);
  assign n24234 = n32147 | n32149;
  assign n24235 = x133 & x156;
  assign n24236 = n24234 & n24235;
  assign n24237 = n24234 | n24235;
  assign n24238 = ~n24236 & n24237;
  assign n24111 = n23760 | n23869;
  assign n32034 = n24111 | n31907;
  assign n32035 = n23513 | n24111;
  assign n32036 = (n31738 & n32034) | (n31738 & n32035) | (n32034 & n32035);
  assign n24118 = n23870 & ~n32038;
  assign n24119 = n32036 & n24118;
  assign n32039 = n24119 | n32028;
  assign n32150 = n24238 | n32039;
  assign n32040 = n23876 | n24119;
  assign n32151 = n24238 | n32040;
  assign n32152 = (n31903 & n32150) | (n31903 & n32151) | (n32150 & n32151);
  assign n32153 = n24238 & n32039;
  assign n32154 = n24238 & n32040;
  assign n32155 = (n31903 & n32153) | (n31903 & n32154) | (n32153 & n32154);
  assign n24241 = n32152 & ~n32155;
  assign n24242 = x132 & x157;
  assign n24243 = ~n24241 & n24242;
  assign n24244 = n24241 & ~n24242;
  assign n24245 = n24243 | n24244;
  assign n32156 = ~n24109 & n24245;
  assign n32157 = ~n32023 & n32156;
  assign n32158 = n24109 & ~n24245;
  assign n32159 = (~n24245 & n32023) | (~n24245 & n32158) | (n32023 & n32158);
  assign n24248 = n32157 | n32159;
  assign n24249 = x131 & x158;
  assign n24250 = n24248 & n24249;
  assign n24251 = n24248 | n24249;
  assign n24252 = ~n24250 & n24251;
  assign n35926 = n23887 | n31905;
  assign n35927 = n23887 | n31904;
  assign n35928 = (n31731 & n35926) | (n31731 & n35927) | (n35926 & n35927);
  assign n32024 = n23888 & ~n32023;
  assign n32025 = n35928 & n32024;
  assign n32026 = n23894 | n32025;
  assign n32160 = n24252 | n32026;
  assign n32161 = n24252 | n32025;
  assign n32162 = (n31896 & n32160) | (n31896 & n32161) | (n32160 & n32161);
  assign n32163 = n24252 & n32026;
  assign n32164 = n24252 & n32025;
  assign n32165 = (n31896 & n32163) | (n31896 & n32164) | (n32163 & n32164);
  assign n24255 = n32162 & ~n32165;
  assign n24256 = x130 & x159;
  assign n24257 = n24255 | n24256;
  assign n24258 = n24255 & n24256;
  assign n24259 = n24257 & ~n24258;
  assign n23907 = n31829 | n31997;
  assign n24260 = n31896 | n23894;
  assign n32166 = ~n23894 & n23895;
  assign n32167 = (n23895 & ~n31896) | (n23895 & n32166) | (~n31896 & n32166);
  assign n24262 = n24260 & n32167;
  assign n32168 = n23909 | n24262;
  assign n32169 = (n23907 & n24262) | (n23907 & n32168) | (n24262 & n32168);
  assign n24264 = ~n24259 & n32169;
  assign n24265 = n24259 & ~n32169;
  assign n24266 = n24264 | n24265;
  assign n24267 = n23913 | n24266;
  assign n24268 = n23916 | n24267;
  assign n24269 = n31888 | n23913;
  assign n24270 = n23914 & n24266;
  assign n24271 = n24269 & n24270;
  assign n24272 = n24268 & ~n24271;
  assign n24273 = x129 & x160;
  assign n24274 = n24272 | n24273;
  assign n24275 = n24272 & n24273;
  assign n24276 = n24274 & ~n24275;
  assign n32170 = n23920 | n24090;
  assign n32171 = (n23920 & n32019) | (n23920 & n32170) | (n32019 & n32170);
  assign n24278 = n24276 | n32171;
  assign n24279 = n24276 & n32171;
  assign n24280 = n24278 & ~n24279;
  assign n24281 = n24096 & n24280;
  assign n24282 = n24096 | n24280;
  assign n24283 = ~n24281 & n24282;
  assign n24284 = n24095 & n24283;
  assign n24285 = n24094 & n24284;
  assign n24286 = n24093 | n24283;
  assign n24287 = n24074 | n24286;
  assign n24288 = ~n24285 & n24287;
  assign n24289 = x127 & x162;
  assign n24290 = n24288 & n24289;
  assign n24291 = n24288 | n24289;
  assign n24292 = ~n24290 & n24291;
  assign n24293 = x126 & x163;
  assign n24294 = n24292 & n24293;
  assign n24295 = n24292 | n24293;
  assign n24296 = ~n24294 & n24295;
  assign n24297 = n32017 | n24296;
  assign n24298 = n32017 & n24296;
  assign n24299 = n24297 & ~n24298;
  assign n24300 = n31881 | n23941;
  assign n32172 = ~n23941 & n23942;
  assign n32173 = (n23942 & ~n31881) | (n23942 & n32172) | (~n31881 & n32172);
  assign n24302 = n24300 & n32173;
  assign n24303 = n24068 | n24302;
  assign n24304 = n24299 | n24303;
  assign n24305 = n24299 & n24303;
  assign n24306 = n24304 & ~n24305;
  assign n24307 = n24072 & n24306;
  assign n24308 = n24072 | n24306;
  assign n24309 = ~n24307 & n24308;
  assign n24310 = ~n32014 & n24309;
  assign n24311 = n32014 & ~n24309;
  assign n24312 = n24310 | n24311;
  assign n24313 = x124 & x165;
  assign n24314 = n24312 & n24313;
  assign n24315 = n24312 | n24313;
  assign n24316 = ~n24314 & n24315;
  assign n24317 = n24062 & n24316;
  assign n24318 = n24062 | n24316;
  assign n24319 = ~n24317 & n24318;
  assign n24320 = n24061 & n24319;
  assign n24321 = n24061 | n24319;
  assign n24322 = ~n24320 & n24321;
  assign n24323 = n24060 & n24322;
  assign n24324 = n24060 | n24322;
  assign n24325 = ~n24323 & n24324;
  assign n24326 = n24059 & n24325;
  assign n24327 = n24059 | n24325;
  assign n24328 = ~n24326 & n24327;
  assign n24329 = n24054 | n24328;
  assign n24330 = n24054 & n24328;
  assign n24331 = n24329 & ~n24330;
  assign n24332 = ~n32012 & n24331;
  assign n24333 = n32012 & ~n24331;
  assign n24334 = n24332 | n24333;
  assign n24335 = x120 & x169;
  assign n24336 = n24334 & n24335;
  assign n24337 = n24334 | n24335;
  assign n24338 = ~n24336 & n24337;
  assign n24339 = n24040 & n24338;
  assign n24340 = n24040 | n24338;
  assign n24341 = ~n24339 & n24340;
  assign n24342 = n24039 & n24341;
  assign n24343 = n24039 | n24341;
  assign n24344 = ~n24342 & n24343;
  assign n24345 = n24038 & n24344;
  assign n24346 = n24038 | n24344;
  assign n24347 = ~n24345 & n24346;
  assign n24348 = n24036 & n24347;
  assign n24349 = n24036 | n24347;
  assign n24350 = ~n24348 & n24349;
  assign n24351 = n24035 & n24350;
  assign n24352 = n24035 | n24350;
  assign n24353 = ~n24351 & n24352;
  assign n24354 = n24034 | n24353;
  assign n24355 = n24034 & n24353;
  assign n24356 = n24354 & ~n24355;
  assign n32174 = n24001 & n24002;
  assign n32175 = (n24001 & n32010) | (n24001 & n32174) | (n32010 & n32174);
  assign n24359 = n24356 & ~n32175;
  assign n24360 = ~n24356 & n32175;
  assign n24361 = n24359 | n24360;
  assign n24362 = x116 & x173;
  assign n24363 = n24361 & n24362;
  assign n24364 = n24361 | n24362;
  assign n24365 = ~n24363 & n24364;
  assign n24366 = n24033 & n24365;
  assign n24367 = n24033 | n24365;
  assign n24368 = ~n24366 & n24367;
  assign n24369 = n24032 & n24368;
  assign n24370 = n24032 | n24368;
  assign n24371 = ~n24369 & n24370;
  assign n24372 = n24031 & n24371;
  assign n24373 = n24031 | n24371;
  assign n24374 = ~n24372 & n24373;
  assign n24375 = n24029 | n24374;
  assign n24376 = n24029 & n24374;
  assign n24377 = n24375 & ~n24376;
  assign n24378 = n23672 | n24024;
  assign n24379 = n24023 & n24378;
  assign n24380 = n24377 & ~n24379;
  assign n24381 = ~n24377 & n24379;
  assign n24382 = n24380 | n24381;
  assign n24383 = x115 & x175;
  assign n24384 = n24369 | n24372;
  assign n24385 = x116 & x174;
  assign n24386 = n24363 | n24366;
  assign n24387 = x118 & x172;
  assign n24388 = n24348 | n24351;
  assign n24389 = x119 & x171;
  assign n24390 = n24342 | n24345;
  assign n24391 = x120 & x170;
  assign n32176 = n24336 | n24338;
  assign n32177 = (n24040 & n24336) | (n24040 & n32176) | (n24336 & n32176);
  assign n24393 = n32012 & n24331;
  assign n24394 = n24055 & n24325;
  assign n24395 = n24055 | n24325;
  assign n24396 = ~n24394 & n24395;
  assign n24397 = n24054 & n24396;
  assign n24398 = n24054 | n24396;
  assign n24399 = n24056 & n24398;
  assign n24400 = ~n24397 & n24399;
  assign n24401 = n24393 | n24400;
  assign n24402 = n24394 | n24397;
  assign n24403 = n24320 | n24323;
  assign n32178 = n24314 | n24316;
  assign n32179 = (n24062 & n24314) | (n24062 & n32178) | (n24314 & n32178);
  assign n32180 = n24307 | n32014;
  assign n32181 = (n24307 & n24309) | (n24307 & n32180) | (n24309 & n32180);
  assign n24407 = n32017 & n24292;
  assign n24408 = n32017 | n24292;
  assign n24409 = n24293 & n24408;
  assign n24410 = ~n24407 & n24409;
  assign n32182 = n24299 | n24410;
  assign n32183 = (n24303 & n24410) | (n24303 & n32182) | (n24410 & n32182);
  assign n24412 = n24281 | n24285;
  assign n35929 = n24255 & n32168;
  assign n35930 = n24255 & n24262;
  assign n35931 = (n23907 & n35929) | (n23907 & n35930) | (n35929 & n35930);
  assign n35932 = (n24256 & n24258) | (n24256 & n32168) | (n24258 & n32168);
  assign n37485 = n24256 & n24262;
  assign n37486 = (n24255 & n24256) | (n24255 & n37485) | (n24256 & n37485);
  assign n35934 = (n23907 & n35932) | (n23907 & n37486) | (n35932 & n37486);
  assign n24416 = ~n35931 & n35934;
  assign n35935 = n23914 | n24416;
  assign n35936 = (n24266 & n24416) | (n24266 & n35935) | (n24416 & n35935);
  assign n32186 = (n24269 & n24416) | (n24269 & n35936) | (n24416 & n35936);
  assign n32187 = n24248 | n32026;
  assign n32188 = n24248 | n32025;
  assign n32189 = (n31896 & n32187) | (n31896 & n32188) | (n32187 & n32188);
  assign n32190 = ~n23888 & n32023;
  assign n32191 = (n23888 & n35928) | (n23888 & ~n32190) | (n35928 & ~n32190);
  assign n24421 = n24248 & n32191;
  assign n32192 = n24421 & n32025;
  assign n32193 = (n24421 & n31896) | (n24421 & n32192) | (n31896 & n32192);
  assign n24423 = n32189 & ~n32193;
  assign n24426 = n24249 | n24423;
  assign n24428 = n24119 | n24234;
  assign n32196 = n24428 | n32028;
  assign n32197 = n23876 | n24428;
  assign n32198 = (n31903 & n32196) | (n31903 & n32197) | (n32196 & n32197);
  assign n24432 = n32036 & ~n32038;
  assign n24433 = n23870 | n24432;
  assign n24434 = n24234 & n24433;
  assign n24430 = n23883 | n24119;
  assign n32199 = n24430 & n24434;
  assign n32200 = (n24434 & n31903) | (n24434 & n32199) | (n31903 & n32199);
  assign n24436 = n32198 & ~n32200;
  assign n24437 = n24235 & n24436;
  assign n32194 = n24109 & n24241;
  assign n32201 = n24437 | n32194;
  assign n32202 = n24241 | n24437;
  assign n32203 = (n32023 & n32201) | (n32023 & n32202) | (n32201 & n32202);
  assign n35937 = n24134 & n32052;
  assign n35938 = n24134 & n35874;
  assign n35939 = (n31751 & n35937) | (n31751 & n35938) | (n35937 & n35938);
  assign n24445 = n35872 & ~n35939;
  assign n24446 = n23856 | n24445;
  assign n24447 = n24220 & n24446;
  assign n24443 = n23765 | n24137;
  assign n32212 = n24443 & n24447;
  assign n32213 = (n24447 & n31915) | (n24447 & n32212) | (n31915 & n32212);
  assign n35940 = n24137 | n24220;
  assign n35941 = n32046 | n35940;
  assign n32215 = n24220 | n32057;
  assign n32216 = (n31915 & n35941) | (n31915 & n32215) | (n35941 & n32215);
  assign n24450 = ~n32213 & n32216;
  assign n24451 = n24221 & n24450;
  assign n32204 = n24224 | n32056;
  assign n32205 = n24224 | n32057;
  assign n32206 = (n31915 & n32204) | (n31915 & n32205) | (n32204 & n32205);
  assign n32207 = n24224 & n32056;
  assign n32208 = n24224 & n32057;
  assign n32209 = (n31915 & n32207) | (n31915 & n32208) | (n32207 & n32208);
  assign n24441 = n32206 & ~n32209;
  assign n32210 = n24127 & n24441;
  assign n32217 = n24451 | n32210;
  assign n32218 = n24441 | n24451;
  assign n32219 = (n32038 & n32217) | (n32038 & n32218) | (n32217 & n32218);
  assign n32221 = n24142 & n24213;
  assign n35942 = (n24134 & n24213) | (n24134 & n32221) | (n24213 & n32221);
  assign n32222 = (n32053 & n35942) | (n32053 & n32221) | (n35942 & n32221);
  assign n24454 = n35917 | n24206;
  assign n32223 = n24454 | n32059;
  assign n32224 = n23848 | n24454;
  assign n35943 = (n31928 & n32223) | (n31928 & n32224) | (n32223 & n32224);
  assign n35944 = (n23772 & n32223) | (n23772 & n32224) | (n32223 & n32224);
  assign n35945 = (n31572 & n35943) | (n31572 & n35944) | (n35943 & n35944);
  assign n35946 = n23842 | n35915;
  assign n35947 = (n23842 & ~n24150) | (n23842 & n35946) | (~n24150 & n35946);
  assign n24459 = n24206 & n35947;
  assign n24456 = n23780 | n35917;
  assign n32226 = n24456 & n24459;
  assign n35948 = (n24459 & n31928) | (n24459 & n32226) | (n31928 & n32226);
  assign n35949 = (n23772 & n24459) | (n23772 & n32226) | (n24459 & n32226);
  assign n35950 = (n31572 & n35948) | (n31572 & n35949) | (n35948 & n35949);
  assign n24461 = n35945 & ~n35950;
  assign n24462 = n24207 & n24461;
  assign n32262 = n24195 & n24202;
  assign n35951 = (n24149 & n24195) | (n24149 & n32262) | (n24195 & n32262);
  assign n32263 = (n32071 & n35951) | (n32071 & n32262) | (n35951 & n32262);
  assign n31943 = (n31588 & n31941) | (n31588 & n31942) | (n31941 & n31942);
  assign n24473 = x141 & x149;
  assign n24474 = x142 & x148;
  assign n24478 = x143 & x147;
  assign n32243 = n23808 & n24166;
  assign n35952 = n23806 & n32243;
  assign n37866 = n24478 & n35952;
  assign n37867 = n24478 & n32243;
  assign n37868 = (n37468 & n37866) | (n37468 & n37867) | (n37866 & n37867);
  assign n37869 = (n23448 & n32243) | (n23448 & n35952) | (n32243 & n35952);
  assign n37870 = n32243 & n35952;
  assign n37871 = (n37462 & n37869) | (n37462 & n37870) | (n37869 & n37870);
  assign n37764 = (n32243 & n35952) | (n32243 & n37466) | (n35952 & n37466);
  assign n37765 = (n35586 & n37871) | (n35586 & n37764) | (n37871 & n37764);
  assign n37768 = n24478 & n37765;
  assign n37769 = (n35438 & n37868) | (n35438 & n37768) | (n37868 & n37768);
  assign n37766 = (n24169 & n24478) | (n24169 & n37769) | (n24478 & n37769);
  assign n37489 = (n35884 & n37766) | (n35884 & n37769) | (n37766 & n37769);
  assign n37490 = (n35886 & n37766) | (n35886 & n37769) | (n37766 & n37769);
  assign n35961 = (n35743 & n37489) | (n35743 & n37490) | (n37489 & n37490);
  assign n37872 = n24478 | n35952;
  assign n37873 = n24478 | n32243;
  assign n37874 = (n37468 & n37872) | (n37468 & n37873) | (n37872 & n37873);
  assign n37772 = n24478 | n37765;
  assign n37773 = (n35438 & n37874) | (n35438 & n37772) | (n37874 & n37772);
  assign n37770 = n24169 | n37773;
  assign n37493 = (n35884 & n37770) | (n35884 & n37773) | (n37770 & n37773);
  assign n37494 = (n35886 & n37770) | (n35886 & n37773) | (n37770 & n37773);
  assign n35964 = (n35743 & n37493) | (n35743 & n37494) | (n37493 & n37494);
  assign n24481 = ~n35961 & n35964;
  assign n32248 = n24173 & n24481;
  assign n32249 = (n24481 & n35891) | (n24481 & n32248) | (n35891 & n32248);
  assign n32250 = n24173 | n24481;
  assign n32251 = n35891 | n32250;
  assign n24484 = ~n32249 & n32251;
  assign n24485 = n24474 & n24484;
  assign n24486 = n24474 | n24484;
  assign n24487 = ~n24485 & n24486;
  assign n24488 = n24473 & n24487;
  assign n24489 = n24473 | n24487;
  assign n24490 = ~n24488 & n24489;
  assign n24468 = n23825 & n24181;
  assign n24466 = n23468 | n23826;
  assign n32234 = n23470 | n24466;
  assign n32236 = n24468 & n32234;
  assign n32253 = n24179 | n32236;
  assign n35967 = ~n24490 & n32253;
  assign n35965 = n24179 | n24466;
  assign n35966 = (n24179 & n24468) | (n24179 & n35965) | (n24468 & n35965);
  assign n35968 = ~n24490 & n35966;
  assign n35969 = (n35760 & n35967) | (n35760 & n35968) | (n35967 & n35968);
  assign n35970 = n24490 & ~n32253;
  assign n35971 = n24490 & ~n35966;
  assign n35972 = (~n35760 & n35970) | (~n35760 & n35971) | (n35970 & n35971);
  assign n24494 = n35969 | n35972;
  assign n24495 = x140 & x150;
  assign n24496 = n24494 & n24495;
  assign n24497 = n24494 | n24495;
  assign n24498 = ~n24496 & n24497;
  assign n35973 = n23826 | n24181;
  assign n35974 = n32075 | n35973;
  assign n32232 = n24181 | n35896;
  assign n32233 = (n35760 & n35974) | (n35760 & n32232) | (n35974 & n32232);
  assign n32237 = n24466 & n24468;
  assign n32238 = (n35760 & n32236) | (n35760 & n32237) | (n32236 & n32237);
  assign n24470 = n32233 & ~n32238;
  assign n24471 = n24182 & n24470;
  assign n32228 = n24188 & n32083;
  assign n32239 = n24471 | n32228;
  assign n32255 = n24498 & ~n32239;
  assign n32229 = n24159 & n24188;
  assign n32240 = n24471 | n32229;
  assign n32256 = n24498 & ~n32240;
  assign n32257 = (~n31943 & n32255) | (~n31943 & n32256) | (n32255 & n32256);
  assign n32258 = ~n24498 & n32239;
  assign n32259 = ~n24498 & n32240;
  assign n32260 = (n31943 & n32258) | (n31943 & n32259) | (n32258 & n32259);
  assign n24501 = n32257 | n32260;
  assign n24502 = x139 & x151;
  assign n24503 = n24501 | n24502;
  assign n24504 = n24501 & n24502;
  assign n24505 = n24503 & ~n24504;
  assign n32264 = n24188 | n32083;
  assign n32265 = n24159 | n24188;
  assign n35975 = (n31941 & n32264) | (n31941 & n32265) | (n32264 & n32265);
  assign n35976 = (n31942 & n32264) | (n31942 & n32265) | (n32264 & n32265);
  assign n35977 = (n31588 & n35975) | (n31588 & n35976) | (n35975 & n35976);
  assign n32268 = n24189 & ~n32229;
  assign n35978 = ~n24188 & n24189;
  assign n35979 = (n24189 & ~n32083) | (n24189 & n35978) | (~n32083 & n35978);
  assign n35980 = (~n31941 & n32268) | (~n31941 & n35979) | (n32268 & n35979);
  assign n35981 = (~n31942 & n32268) | (~n31942 & n35979) | (n32268 & n35979);
  assign n35982 = (~n31588 & n35980) | (~n31588 & n35981) | (n35980 & n35981);
  assign n24509 = n35977 & n35982;
  assign n32270 = n24505 | n24509;
  assign n32271 = n32263 | n32270;
  assign n32272 = n24505 & n24509;
  assign n32273 = (n24505 & n32263) | (n24505 & n32272) | (n32263 & n32272);
  assign n24513 = n32271 & ~n32273;
  assign n24514 = x138 & x152;
  assign n24515 = n24513 | n24514;
  assign n24516 = n24513 & n24514;
  assign n24517 = n24515 & ~n24516;
  assign n32275 = n24195 | n24202;
  assign n35983 = n24149 | n32275;
  assign n32276 = (n32071 & n35983) | (n32071 & n32275) | (n35983 & n32275);
  assign n35984 = n24196 & ~n35951;
  assign n35985 = n24196 & ~n32262;
  assign n35986 = (~n32071 & n35984) | (~n32071 & n35985) | (n35984 & n35985);
  assign n24520 = n32276 & n35986;
  assign n32277 = ~n24517 & n24520;
  assign n32278 = (~n24517 & n35950) | (~n24517 & n32277) | (n35950 & n32277);
  assign n32279 = n24517 & ~n24520;
  assign n32280 = ~n35950 & n32279;
  assign n24524 = n32278 | n32280;
  assign n24525 = x137 & x153;
  assign n24526 = n24524 & n24525;
  assign n24527 = n24524 | n24525;
  assign n24528 = ~n24526 & n24527;
  assign n32281 = ~n24462 & n24528;
  assign n32282 = ~n32222 & n32281;
  assign n32283 = n24462 & ~n24528;
  assign n32284 = (~n24528 & n32222) | (~n24528 & n32283) | (n32222 & n32283);
  assign n24531 = n32282 | n32284;
  assign n24532 = x136 & x154;
  assign n24533 = n24531 | n24532;
  assign n24534 = n24531 & n24532;
  assign n24535 = n24533 & ~n24534;
  assign n32286 = n24142 | n24213;
  assign n35987 = n24134 | n32286;
  assign n32287 = (n32053 & n35987) | (n32053 & n32286) | (n35987 & n32286);
  assign n35988 = n24214 & ~n35942;
  assign n37495 = ~n24142 & n24214;
  assign n37496 = (~n24213 & n24214) | (~n24213 & n37495) | (n24214 & n37495);
  assign n35990 = (~n32053 & n35988) | (~n32053 & n37496) | (n35988 & n37496);
  assign n24538 = n32287 & n35990;
  assign n32288 = ~n24535 & n24538;
  assign n32289 = (~n24535 & n32213) | (~n24535 & n32288) | (n32213 & n32288);
  assign n32290 = n24535 & ~n24538;
  assign n32291 = ~n32213 & n32290;
  assign n24542 = n32289 | n32291;
  assign n24543 = x135 & x155;
  assign n24544 = n24542 & n24543;
  assign n24545 = n24542 | n24543;
  assign n24546 = ~n24544 & n24545;
  assign n24547 = n32219 | n24546;
  assign n24548 = n32219 & n24546;
  assign n24549 = n24547 & ~n24548;
  assign n24550 = x134 & x156;
  assign n24551 = n24549 | n24550;
  assign n24552 = n24549 & n24550;
  assign n24553 = n24551 & ~n24552;
  assign n32292 = n24127 | n24441;
  assign n32293 = n32038 | n32292;
  assign n35991 = ~n24127 & n24225;
  assign n35992 = (n24225 & ~n24441) | (n24225 & n35991) | (~n24441 & n35991);
  assign n32295 = n24225 & ~n24441;
  assign n32296 = (~n32038 & n35992) | (~n32038 & n32295) | (n35992 & n32295);
  assign n24556 = n32293 & n32296;
  assign n32297 = n24556 | n32199;
  assign n32298 = n24434 | n24556;
  assign n32299 = (n31903 & n32297) | (n31903 & n32298) | (n32297 & n32298);
  assign n24558 = ~n24553 & n32299;
  assign n24559 = n24553 & ~n32299;
  assign n24560 = n24558 | n24559;
  assign n24561 = x133 & x157;
  assign n24562 = n24560 & n24561;
  assign n24563 = n24560 | n24561;
  assign n24564 = ~n24562 & n24563;
  assign n24565 = n32203 | n24564;
  assign n24566 = n32203 & n24564;
  assign n24567 = n24565 & ~n24566;
  assign n24568 = x132 & x158;
  assign n24569 = ~n24567 & n24568;
  assign n24570 = n24567 & ~n24568;
  assign n24571 = n24569 | n24570;
  assign n32300 = n24109 | n24241;
  assign n32301 = n32023 | n32300;
  assign n35993 = ~n24109 & n24242;
  assign n35994 = (~n24241 & n24242) | (~n24241 & n35993) | (n24242 & n35993);
  assign n32303 = (n24243 & ~n32023) | (n24243 & n35994) | (~n32023 & n35994);
  assign n24574 = n32301 & n32303;
  assign n35995 = n24574 | n32025;
  assign n35996 = (n24421 & n24574) | (n24421 & n35995) | (n24574 & n35995);
  assign n32305 = n24421 | n24574;
  assign n32306 = (n31896 & n35996) | (n31896 & n32305) | (n35996 & n32305);
  assign n24576 = n24571 & n32306;
  assign n24577 = n24571 | n32306;
  assign n24578 = ~n24576 & n24577;
  assign n24579 = n24426 & n24578;
  assign n24424 = n24249 & n24423;
  assign n32307 = n24424 & n24579;
  assign n32308 = (n24579 & n32169) | (n24579 & n32307) | (n32169 & n32307);
  assign n24581 = n24424 | n24578;
  assign n32309 = n24255 | n24581;
  assign n32310 = (n24581 & n32169) | (n24581 & n32309) | (n32169 & n32309);
  assign n24583 = ~n32308 & n32310;
  assign n24584 = x131 & x159;
  assign n24585 = x130 & x160;
  assign n24586 = n24584 | n24585;
  assign n24587 = n24584 & n24585;
  assign n24588 = n24586 & ~n24587;
  assign n24589 = n24583 | n24588;
  assign n24590 = n24583 & n24588;
  assign n24591 = n24589 & ~n24590;
  assign n24592 = ~n32186 & n24591;
  assign n24593 = n32186 & ~n24591;
  assign n24594 = n24592 | n24593;
  assign n24595 = n24275 | n24594;
  assign n24596 = n24279 | n24595;
  assign n24597 = n24275 | n32171;
  assign n24598 = n24274 & n24594;
  assign n24599 = n24597 & n24598;
  assign n24600 = n24596 & ~n24599;
  assign n24601 = x129 & x161;
  assign n24602 = n24600 & n24601;
  assign n24603 = n24600 | n24601;
  assign n24604 = ~n24602 & n24603;
  assign n24605 = x128 & x162;
  assign n24606 = n24604 & n24605;
  assign n24607 = n24604 | n24605;
  assign n24608 = ~n24606 & n24607;
  assign n24609 = ~n24412 & n24608;
  assign n24610 = n24412 & ~n24608;
  assign n24611 = n24609 | n24610;
  assign n24612 = n24290 | n24611;
  assign n24613 = n24407 | n24612;
  assign n24073 = n31881 & n23941;
  assign n32311 = n24077 | n24289;
  assign n32312 = (n24077 & n24288) | (n24077 & n32311) | (n24288 & n32311);
  assign n24615 = n24073 | n32312;
  assign n24616 = n24291 & n24611;
  assign n24617 = n24615 & n24616;
  assign n24618 = n24613 & ~n24617;
  assign n24619 = x127 & x163;
  assign n24620 = n24618 & n24619;
  assign n24621 = n24618 | n24619;
  assign n24622 = ~n24620 & n24621;
  assign n24623 = n32183 | n24622;
  assign n24624 = n32183 & n24622;
  assign n24625 = n24623 & ~n24624;
  assign n24626 = x126 & x164;
  assign n24627 = x125 & x165;
  assign n24628 = n24626 & n24627;
  assign n24629 = n24626 | n24627;
  assign n24630 = ~n24628 & n24629;
  assign n24631 = n24625 & n24630;
  assign n24632 = n24625 | n24630;
  assign n24633 = ~n24631 & n24632;
  assign n24634 = n32181 | n24633;
  assign n24635 = n32181 & n24633;
  assign n24636 = n24634 & ~n24635;
  assign n24637 = x124 & x166;
  assign n24638 = n24636 | n24637;
  assign n24639 = n24636 & n24637;
  assign n24640 = n24638 & ~n24639;
  assign n24641 = n32179 | n24640;
  assign n24642 = n32179 & n24640;
  assign n24643 = n24641 & ~n24642;
  assign n24644 = x123 & x167;
  assign n24645 = n24643 | n24644;
  assign n24646 = n24643 & n24644;
  assign n24647 = n24645 & ~n24646;
  assign n24648 = n24403 | n24647;
  assign n24649 = n24403 & n24647;
  assign n24650 = n24648 & ~n24649;
  assign n24651 = x122 & x168;
  assign n24652 = n24650 | n24651;
  assign n24653 = n24650 & n24651;
  assign n24654 = n24652 & ~n24653;
  assign n24655 = n24402 | n24654;
  assign n24656 = n24402 & n24654;
  assign n24657 = n24655 & ~n24656;
  assign n24658 = ~n24401 & n24657;
  assign n24659 = n24401 & ~n24657;
  assign n24660 = n24658 | n24659;
  assign n24661 = x121 & x169;
  assign n24662 = n24660 & n24661;
  assign n24663 = n24660 | n24661;
  assign n24664 = ~n24662 & n24663;
  assign n24665 = n32177 & n24664;
  assign n24666 = n32177 | n24664;
  assign n24667 = ~n24665 & n24666;
  assign n24668 = n24391 & n24667;
  assign n24669 = n24391 | n24667;
  assign n24670 = ~n24668 & n24669;
  assign n24671 = n24390 & n24670;
  assign n24672 = n24390 | n24670;
  assign n24673 = ~n24671 & n24672;
  assign n24674 = n24389 & n24673;
  assign n24675 = n24389 | n24673;
  assign n24676 = ~n24674 & n24675;
  assign n24677 = n24388 & n24676;
  assign n24678 = n24388 | n24676;
  assign n24679 = ~n24677 & n24678;
  assign n24680 = n24387 | n24679;
  assign n24681 = n24387 & n24679;
  assign n24682 = n24680 & ~n24681;
  assign n24683 = n24355 | n32175;
  assign n24684 = n24354 & n24683;
  assign n24685 = n24682 & ~n24684;
  assign n24686 = ~n24682 & n24684;
  assign n24687 = n24685 | n24686;
  assign n24688 = x117 & x173;
  assign n24689 = n24687 & n24688;
  assign n24690 = n24687 | n24688;
  assign n24691 = ~n24689 & n24690;
  assign n24692 = n24386 & n24691;
  assign n24693 = n24386 | n24691;
  assign n24694 = ~n24692 & n24693;
  assign n24695 = n24385 & n24694;
  assign n24696 = n24385 | n24694;
  assign n24697 = ~n24695 & n24696;
  assign n24698 = n24384 & n24697;
  assign n24699 = n24384 | n24697;
  assign n24700 = ~n24698 & n24699;
  assign n24701 = n24383 | n24700;
  assign n24702 = n24383 & n24700;
  assign n24703 = n24701 & ~n24702;
  assign n24704 = n24376 | n24379;
  assign n24705 = n24375 & n24704;
  assign n24706 = n24703 & ~n24705;
  assign n24707 = ~n24703 & n24705;
  assign n24708 = n24706 | n24707;
  assign n24709 = x116 & x175;
  assign n24710 = n24695 | n24698;
  assign n24711 = x117 & x174;
  assign n24712 = n24689 | n24692;
  assign n24713 = x119 & x172;
  assign n24714 = n24674 | n24677;
  assign n24715 = x120 & x171;
  assign n32313 = n24668 | n24670;
  assign n32314 = (n24390 & n24668) | (n24390 & n32313) | (n24668 & n32313);
  assign n24717 = x121 & x170;
  assign n24718 = n24662 | n24665;
  assign n32315 = n24394 & n24650;
  assign n32316 = (n24397 & n24650) | (n24397 & n32315) | (n24650 & n32315);
  assign n32317 = n24394 | n24650;
  assign n32318 = n24397 | n32317;
  assign n24722 = n24651 & n32318;
  assign n24723 = ~n32316 & n24722;
  assign n32319 = n24657 | n24723;
  assign n32320 = (n24401 & n24723) | (n24401 & n32319) | (n24723 & n32319);
  assign n32321 = n24320 & n24643;
  assign n32322 = (n24323 & n24643) | (n24323 & n32321) | (n24643 & n32321);
  assign n32323 = n24320 | n24643;
  assign n32325 = n24644 & n32323;
  assign n32326 = (n24323 & n24644) | (n24323 & n32325) | (n24644 & n32325);
  assign n24728 = ~n32322 & n32326;
  assign n24729 = n32316 | n24728;
  assign n24730 = x124 & x167;
  assign n24731 = x123 & x168;
  assign n24732 = n24730 & n24731;
  assign n24733 = n24730 | n24731;
  assign n24734 = ~n24732 & n24733;
  assign n24735 = n32179 & n24636;
  assign n32327 = (n24637 & n24639) | (n24637 & n32179) | (n24639 & n32179);
  assign n24738 = ~n24735 & n32327;
  assign n32328 = n24738 | n32321;
  assign n32329 = n24643 | n24738;
  assign n32330 = (n24323 & n32328) | (n24323 & n32329) | (n32328 & n32329);
  assign n24740 = n24625 & n24626;
  assign n24741 = n24625 | n24626;
  assign n24742 = ~n24740 & n24741;
  assign n24743 = n32181 & n24742;
  assign n24744 = n32181 | n24742;
  assign n24745 = n24627 & n24744;
  assign n24746 = ~n24743 & n24745;
  assign n32331 = n24636 | n24746;
  assign n32332 = (n24746 & n32179) | (n24746 & n32331) | (n32179 & n32331);
  assign n24748 = n24740 | n24743;
  assign n24749 = x128 & x163;
  assign n32333 = n24281 & n24604;
  assign n32334 = (n24285 & n24604) | (n24285 & n32333) | (n24604 & n32333);
  assign n24751 = x130 & x161;
  assign n24752 = n24583 & n24584;
  assign n24756 = n24567 & n32306;
  assign n32335 = n24567 & n24568;
  assign n32336 = (n24568 & n32306) | (n24568 & n32335) | (n32306 & n32335);
  assign n24759 = ~n24756 & n32336;
  assign n24765 = n24235 | n24436;
  assign n24766 = n24560 & n24765;
  assign n35997 = n24109 | n24235;
  assign n35998 = (n24109 & n24436) | (n24109 & n35997) | (n24436 & n35997);
  assign n32340 = n35998 & n24766;
  assign n32341 = (n24766 & n32023) | (n24766 & n32340) | (n32023 & n32340);
  assign n24771 = n24549 & n32299;
  assign n32344 = (n24550 & n24552) | (n24550 & n32299) | (n24552 & n32299);
  assign n24774 = ~n24771 & n32344;
  assign n24778 = n24221 | n24450;
  assign n24779 = n24542 & n24778;
  assign n35999 = n24127 | n24221;
  assign n36000 = (n24127 & n24450) | (n24127 & n35999) | (n24450 & n35999);
  assign n32350 = n24779 & n36000;
  assign n32351 = (n24779 & n32038) | (n24779 & n32350) | (n32038 & n32350);
  assign n32354 = n24531 & n24538;
  assign n36001 = (n24531 & n32212) | (n24531 & n32354) | (n32212 & n32354);
  assign n36002 = (n24447 & n24531) | (n24447 & n32354) | (n24531 & n32354);
  assign n36003 = (n31915 & n36001) | (n31915 & n36002) | (n36001 & n36002);
  assign n36004 = n24532 & n24538;
  assign n36005 = (n24531 & n24532) | (n24531 & n36004) | (n24532 & n36004);
  assign n36006 = (n24532 & n32212) | (n24532 & n36005) | (n32212 & n36005);
  assign n36007 = (n24447 & n24532) | (n24447 & n36005) | (n24532 & n36005);
  assign n36008 = (n31915 & n36006) | (n31915 & n36007) | (n36006 & n36007);
  assign n24787 = ~n36003 & n36008;
  assign n24791 = n24142 | n24462;
  assign n32360 = n24134 | n24791;
  assign n32361 = (n24791 & n32053) | (n24791 & n32360) | (n32053 & n32360);
  assign n24811 = n24182 | n24470;
  assign n24812 = n24494 & n24811;
  assign n32388 = n24159 | n24471;
  assign n32390 = n24812 & n32388;
  assign n37503 = n24179 & n24487;
  assign n37504 = (n24487 & n32236) | (n24487 & n37503) | (n32236 & n37503);
  assign n36010 = n24487 & n35966;
  assign n36011 = (n35760 & n37504) | (n35760 & n36010) | (n37504 & n36010);
  assign n36012 = (n24473 & n24488) | (n24473 & n32253) | (n24488 & n32253);
  assign n36013 = (n24473 & n24488) | (n24473 & n35966) | (n24488 & n35966);
  assign n36014 = (n35760 & n36012) | (n35760 & n36013) | (n36012 & n36013);
  assign n24820 = ~n36011 & n36014;
  assign n24823 = x142 & x149;
  assign n24825 = x143 & x148;
  assign n36015 = n24481 | n35961;
  assign n36016 = (n24173 & n35961) | (n24173 & n36015) | (n35961 & n36015);
  assign n32405 = n24825 & n36016;
  assign n37875 = n24478 & n24825;
  assign n37912 = n37765 & n37875;
  assign n37929 = n35952 & n37875;
  assign n37930 = n32243 & n37875;
  assign n37915 = (n37468 & n37929) | (n37468 & n37930) | (n37929 & n37930);
  assign n37879 = (n35438 & n37912) | (n35438 & n37915) | (n37912 & n37915);
  assign n37876 = (n24169 & n37879) | (n24169 & n37875) | (n37879 & n37875);
  assign n37776 = (n35884 & n37876) | (n35884 & n37879) | (n37876 & n37879);
  assign n37777 = (n35886 & n37876) | (n35886 & n37879) | (n37876 & n37879);
  assign n37499 = (n35743 & n37776) | (n35743 & n37777) | (n37776 & n37777);
  assign n36018 = (n24481 & n24825) | (n24481 & n37499) | (n24825 & n37499);
  assign n32407 = (n35891 & n32405) | (n35891 & n36018) | (n32405 & n36018);
  assign n32408 = n24825 | n36016;
  assign n37880 = n24478 | n24825;
  assign n37916 = (n24825 & n37765) | (n24825 & n37880) | (n37765 & n37880);
  assign n37931 = (n24825 & n35952) | (n24825 & n37880) | (n35952 & n37880);
  assign n37932 = (n24825 & n32243) | (n24825 & n37880) | (n32243 & n37880);
  assign n37919 = (n37468 & n37931) | (n37468 & n37932) | (n37931 & n37932);
  assign n37884 = (n35438 & n37916) | (n35438 & n37919) | (n37916 & n37919);
  assign n37881 = (n24169 & n37884) | (n24169 & n37880) | (n37884 & n37880);
  assign n37780 = (n35884 & n37881) | (n35884 & n37884) | (n37881 & n37884);
  assign n37781 = (n35886 & n37881) | (n35886 & n37884) | (n37881 & n37884);
  assign n37502 = (n35743 & n37780) | (n35743 & n37781) | (n37780 & n37781);
  assign n36020 = n24481 | n37502;
  assign n32410 = (n35891 & n32408) | (n35891 & n36020) | (n32408 & n36020);
  assign n24828 = ~n32407 & n32410;
  assign n24829 = n24823 & n24828;
  assign n24830 = n24823 | n24828;
  assign n24831 = ~n24829 & n24830;
  assign n32400 = n24485 | n24487;
  assign n32411 = n24831 | n32400;
  assign n32412 = n24485 | n24831;
  assign n36021 = (n32253 & n32411) | (n32253 & n32412) | (n32411 & n32412);
  assign n36022 = (n32411 & n32412) | (n32411 & n35966) | (n32412 & n35966);
  assign n36023 = (n35760 & n36021) | (n35760 & n36022) | (n36021 & n36022);
  assign n32414 = n24831 & n32400;
  assign n32415 = n24485 & n24831;
  assign n36024 = (n32253 & n32414) | (n32253 & n32415) | (n32414 & n32415);
  assign n36025 = (n32414 & n32415) | (n32414 & n35966) | (n32415 & n35966);
  assign n36026 = (n35760 & n36024) | (n35760 & n36025) | (n36024 & n36025);
  assign n24834 = n36023 & ~n36026;
  assign n24835 = x141 & x150;
  assign n24836 = n24834 | n24835;
  assign n24837 = n24834 & n24835;
  assign n24838 = n24836 & ~n24837;
  assign n37505 = ~n24820 & n24838;
  assign n37506 = ~n32390 & n37505;
  assign n32387 = n24471 | n32083;
  assign n32391 = n24812 & n32387;
  assign n37507 = ~n32391 & n37505;
  assign n36029 = (~n31943 & n37506) | (~n31943 & n37507) | (n37506 & n37507);
  assign n37508 = n24820 & ~n24838;
  assign n37509 = (~n24838 & n32390) | (~n24838 & n37508) | (n32390 & n37508);
  assign n37510 = (~n24838 & n32391) | (~n24838 & n37508) | (n32391 & n37508);
  assign n36032 = (n31943 & n37509) | (n31943 & n37510) | (n37509 & n37510);
  assign n24841 = n36029 | n36032;
  assign n24842 = x140 & x151;
  assign n24843 = n24841 & n24842;
  assign n24844 = n24841 | n24842;
  assign n24845 = ~n24843 & n24844;
  assign n32385 = n24494 | n32240;
  assign n36033 = n24471 | n24494;
  assign n36034 = n32228 | n36033;
  assign n36035 = (n31941 & n32385) | (n31941 & n36034) | (n32385 & n36034);
  assign n36036 = (n31942 & n32385) | (n31942 & n36034) | (n32385 & n36034);
  assign n36037 = (n31588 & n36035) | (n31588 & n36036) | (n36035 & n36036);
  assign n36038 = (n31941 & n32390) | (n31941 & n32391) | (n32390 & n32391);
  assign n36039 = (n31942 & n32390) | (n31942 & n32391) | (n32390 & n32391);
  assign n36040 = (n31588 & n36038) | (n31588 & n36039) | (n36038 & n36039);
  assign n24814 = n36037 & ~n36040;
  assign n24815 = n24495 & n24814;
  assign n32394 = n24501 | n24815;
  assign n32417 = n24845 | n32394;
  assign n32375 = n24501 & n24509;
  assign n32393 = n24815 | n32375;
  assign n32418 = n24845 | n32393;
  assign n32419 = (n32263 & n32417) | (n32263 & n32418) | (n32417 & n32418);
  assign n32420 = n24845 & n32394;
  assign n32421 = n24845 & n32393;
  assign n32422 = (n32263 & n32420) | (n32263 & n32421) | (n32420 & n32421);
  assign n24848 = n32419 & ~n32422;
  assign n24849 = x139 & x152;
  assign n24850 = n24848 | n24849;
  assign n24851 = n24848 & n24849;
  assign n24852 = n24850 & ~n24851;
  assign n36041 = (n24501 & n32375) | (n24501 & n35951) | (n32375 & n35951);
  assign n36042 = (n24501 & n32262) | (n24501 & n32375) | (n32262 & n32375);
  assign n36043 = (n32071 & n36041) | (n32071 & n36042) | (n36041 & n36042);
  assign n36044 = n24502 & n24509;
  assign n36045 = (n24501 & n24502) | (n24501 & n36044) | (n24502 & n36044);
  assign n36046 = (n24502 & n35951) | (n24502 & n36045) | (n35951 & n36045);
  assign n36047 = (n24502 & n32262) | (n24502 & n36045) | (n32262 & n36045);
  assign n36048 = (n32071 & n36046) | (n32071 & n36047) | (n36046 & n36047);
  assign n24807 = ~n36043 & n36048;
  assign n36049 = n24520 | n24807;
  assign n36050 = (n24513 & n24807) | (n24513 & n36049) | (n24807 & n36049);
  assign n32423 = n24852 | n36050;
  assign n32382 = n24513 | n24807;
  assign n32424 = n24852 | n32382;
  assign n32425 = (n35950 & n32423) | (n35950 & n32424) | (n32423 & n32424);
  assign n32426 = n24852 & n36050;
  assign n32427 = n24852 & n32382;
  assign n32428 = (n35950 & n32426) | (n35950 & n32427) | (n32426 & n32427);
  assign n24855 = n32425 & ~n32428;
  assign n24856 = x138 & x153;
  assign n24857 = n24855 | n24856;
  assign n24858 = n24855 & n24856;
  assign n24859 = n24857 & ~n24858;
  assign n24793 = n24207 | n24461;
  assign n24794 = n24524 & n24793;
  assign n32367 = n24513 & n24520;
  assign n32368 = (n24513 & n35950) | (n24513 & n32367) | (n35950 & n32367);
  assign n36051 = n24514 & n24520;
  assign n36052 = (n24513 & n24514) | (n24513 & n36051) | (n24514 & n36051);
  assign n32372 = (n24514 & n35950) | (n24514 & n36052) | (n35950 & n36052);
  assign n24802 = ~n32368 & n32372;
  assign n32373 = n24794 | n24802;
  assign n32429 = n24859 & ~n32373;
  assign n32430 = ~n24802 & n24859;
  assign n32431 = (~n32361 & n32429) | (~n32361 & n32430) | (n32429 & n32430);
  assign n32432 = ~n24859 & n32373;
  assign n32433 = n24802 & ~n24859;
  assign n32434 = (n32361 & n32432) | (n32361 & n32433) | (n32432 & n32433);
  assign n24862 = n32431 | n32434;
  assign n24863 = x137 & x154;
  assign n24864 = n24862 & n24863;
  assign n24865 = n24862 | n24863;
  assign n24866 = ~n24864 & n24865;
  assign n24789 = n24462 | n24524;
  assign n36053 = n24789 | n35942;
  assign n36054 = n24789 | n32221;
  assign n36055 = (n32053 & n36053) | (n32053 & n36054) | (n36053 & n36054);
  assign n32362 = n24525 & ~n24794;
  assign n36056 = (n24525 & ~n32360) | (n24525 & n32362) | (~n32360 & n32362);
  assign n36057 = (n24525 & ~n24791) | (n24525 & n32362) | (~n24791 & n32362);
  assign n36058 = (~n32053 & n36056) | (~n32053 & n36057) | (n36056 & n36057);
  assign n24797 = n36055 & n36058;
  assign n25070 = n24538 | n24797;
  assign n36059 = (n24531 & n24797) | (n24531 & n25070) | (n24797 & n25070);
  assign n32435 = n24866 & ~n36059;
  assign n32365 = n24531 | n24797;
  assign n32436 = n24866 & ~n32365;
  assign n32437 = (~n32213 & n32435) | (~n32213 & n32436) | (n32435 & n32436);
  assign n32438 = ~n24866 & n36059;
  assign n32439 = ~n24866 & n32365;
  assign n32440 = (n32213 & n32438) | (n32213 & n32439) | (n32438 & n32439);
  assign n24869 = n32437 | n32440;
  assign n24870 = x136 & x155;
  assign n24871 = n24869 | n24870;
  assign n24872 = n24869 & n24870;
  assign n24873 = n24871 & ~n24872;
  assign n32441 = ~n24787 & n24873;
  assign n32442 = ~n32351 & n32441;
  assign n32443 = n24787 & ~n24873;
  assign n32444 = (~n24873 & n32351) | (~n24873 & n32443) | (n32351 & n32443);
  assign n24876 = n32442 | n32444;
  assign n24877 = x135 & x156;
  assign n24878 = n24876 & n24877;
  assign n24879 = n24876 | n24877;
  assign n24880 = ~n24878 & n24879;
  assign n32345 = n24542 | n32218;
  assign n32346 = n24542 | n32217;
  assign n32347 = (n32038 & n32345) | (n32038 & n32346) | (n32345 & n32346);
  assign n24781 = n32347 & ~n32351;
  assign n24782 = n24543 & n24781;
  assign n32352 = n24549 | n24782;
  assign n32445 = n24880 | n32352;
  assign n32446 = n24782 | n24880;
  assign n32447 = (n32299 & n32445) | (n32299 & n32446) | (n32445 & n32446);
  assign n32448 = n24880 & n32352;
  assign n32449 = n24782 & n24880;
  assign n32450 = (n32299 & n32448) | (n32299 & n32449) | (n32448 & n32449);
  assign n24883 = n32447 & ~n32450;
  assign n24884 = x134 & x157;
  assign n24885 = ~n24883 & n24884;
  assign n24886 = n24883 & ~n24884;
  assign n24887 = n24885 | n24886;
  assign n32451 = ~n24774 & n24887;
  assign n32452 = ~n32341 & n32451;
  assign n32453 = n24774 & ~n24887;
  assign n32454 = (~n24887 & n32341) | (~n24887 & n32453) | (n32341 & n32453);
  assign n24890 = n32452 | n32454;
  assign n24891 = x133 & x158;
  assign n24892 = n24890 & n24891;
  assign n24893 = n24890 | n24891;
  assign n24894 = ~n24892 & n24893;
  assign n24761 = n24437 | n24560;
  assign n32337 = n24761 | n32194;
  assign n32338 = n24241 | n24761;
  assign n32339 = (n32023 & n32337) | (n32023 & n32338) | (n32337 & n32338);
  assign n24768 = n24561 & ~n32341;
  assign n24769 = n32339 & n24768;
  assign n32342 = n24567 | n24769;
  assign n32455 = n24894 | n32342;
  assign n32456 = n24769 | n24894;
  assign n32457 = (n32306 & n32455) | (n32306 & n32456) | (n32455 & n32456);
  assign n32458 = n24894 & n32342;
  assign n32459 = n24769 & n24894;
  assign n32460 = (n32306 & n32458) | (n32306 & n32459) | (n32458 & n32459);
  assign n24897 = n32457 & ~n32460;
  assign n24898 = x132 & x159;
  assign n24899 = n24897 | n24898;
  assign n24900 = n24897 & n24898;
  assign n24901 = n24899 & ~n24900;
  assign n32461 = ~n24759 & n24901;
  assign n32462 = ~n32308 & n32461;
  assign n32463 = n24759 & ~n24901;
  assign n32464 = (~n24901 & n32308) | (~n24901 & n32463) | (n32308 & n32463);
  assign n24904 = n32462 | n32464;
  assign n24905 = n24752 | n24904;
  assign n24753 = n24583 | n24584;
  assign n24754 = ~n24752 & n24753;
  assign n32465 = n24754 | n24905;
  assign n32466 = (n24905 & n32186) | (n24905 & n32465) | (n32186 & n32465);
  assign n24909 = n24753 & n24904;
  assign n36060 = n24416 | n24584;
  assign n36061 = (n24416 & n24583) | (n24416 & n36060) | (n24583 & n36060);
  assign n32467 = n36061 & n24909;
  assign n32468 = (n24271 & n24909) | (n24271 & n32467) | (n24909 & n32467);
  assign n24911 = n32466 & ~n32468;
  assign n24912 = x131 & x160;
  assign n24913 = n24911 | n24912;
  assign n24914 = ~n32468 & n24912;
  assign n24915 = n32466 & n24914;
  assign n24916 = n24913 & ~n24915;
  assign n24917 = n32186 | n24754;
  assign n32469 = n24585 & ~n24754;
  assign n32470 = (n24585 & ~n32186) | (n24585 & n32469) | (~n32186 & n32469);
  assign n24919 = n24917 & n32470;
  assign n32471 = n24598 | n24919;
  assign n32472 = (n24597 & n24919) | (n24597 & n32471) | (n24919 & n32471);
  assign n24921 = n24916 | n32472;
  assign n24922 = n24916 & n32472;
  assign n24923 = n24921 & ~n24922;
  assign n24924 = n24751 & n24923;
  assign n24925 = n24751 | n24923;
  assign n24926 = ~n24924 & n24925;
  assign n24927 = n24602 | n24926;
  assign n24928 = n32334 | n24927;
  assign n24929 = n24281 | n24602;
  assign n24930 = n24285 | n24929;
  assign n24931 = n24603 & n24926;
  assign n24932 = n24930 & n24931;
  assign n24933 = n24928 & ~n24932;
  assign n24934 = x129 & x162;
  assign n24935 = n24933 & n24934;
  assign n24936 = n24933 | n24934;
  assign n24937 = ~n24935 & n24936;
  assign n32473 = n24281 | n24604;
  assign n32474 = n24285 | n32473;
  assign n24939 = n24605 & ~n32334;
  assign n24940 = n32474 & n24939;
  assign n24941 = n24617 | n24940;
  assign n24942 = n24937 & n24941;
  assign n24943 = n24937 | n24941;
  assign n24944 = ~n24942 & n24943;
  assign n24945 = n24749 & n24944;
  assign n24946 = n24749 | n24944;
  assign n24947 = ~n24945 & n24946;
  assign n32475 = n24620 & n24621;
  assign n32476 = (n24621 & n32183) | (n24621 & n32475) | (n32183 & n32475);
  assign n24950 = n24947 & n32476;
  assign n24951 = n24947 | n32476;
  assign n24952 = ~n24950 & n24951;
  assign n24953 = x127 & x164;
  assign n24954 = n24952 & n24953;
  assign n24955 = n24952 | n24953;
  assign n24956 = ~n24954 & n24955;
  assign n24957 = n24748 & n24956;
  assign n24958 = n24748 | n24956;
  assign n24959 = ~n24957 & n24958;
  assign n24960 = x126 & x165;
  assign n24961 = n24959 & n24960;
  assign n24962 = n24959 | n24960;
  assign n24963 = ~n24961 & n24962;
  assign n24964 = n32332 & n24963;
  assign n24965 = n32332 | n24963;
  assign n24966 = ~n24964 & n24965;
  assign n24967 = x125 & x166;
  assign n24968 = n24966 & n24967;
  assign n24969 = n24966 | n24967;
  assign n24970 = ~n24968 & n24969;
  assign n24971 = n32330 & n24970;
  assign n24972 = n32330 | n24970;
  assign n24973 = ~n24971 & n24972;
  assign n24974 = n24734 & n24973;
  assign n24975 = n24734 | n24973;
  assign n24976 = ~n24974 & n24975;
  assign n24977 = n24729 | n24976;
  assign n24978 = n24729 & n24976;
  assign n24979 = n24977 & ~n24978;
  assign n24980 = ~n32320 & n24979;
  assign n24981 = n32320 & ~n24979;
  assign n24982 = n24980 | n24981;
  assign n24983 = x122 & x169;
  assign n24984 = n24982 & n24983;
  assign n24985 = n24982 | n24983;
  assign n24986 = ~n24984 & n24985;
  assign n24987 = n24718 & n24986;
  assign n24988 = n24718 | n24986;
  assign n24989 = ~n24987 & n24988;
  assign n24990 = n24717 & n24989;
  assign n24991 = n24717 | n24989;
  assign n24992 = ~n24990 & n24991;
  assign n24993 = n32314 & n24992;
  assign n24994 = n32314 | n24992;
  assign n24995 = ~n24993 & n24994;
  assign n24996 = n24715 & n24995;
  assign n24997 = n24715 | n24995;
  assign n24998 = ~n24996 & n24997;
  assign n24999 = n24714 & n24998;
  assign n25000 = n24714 | n24998;
  assign n25001 = ~n24999 & n25000;
  assign n25002 = n24713 & n25001;
  assign n25003 = n24713 | n25001;
  assign n25004 = ~n25002 & n25003;
  assign n25005 = n24681 | n24684;
  assign n25006 = n24680 & n25005;
  assign n25007 = n25004 & ~n25006;
  assign n25008 = ~n25004 & n25006;
  assign n25009 = n25007 | n25008;
  assign n25010 = x118 & x173;
  assign n25011 = n25009 & n25010;
  assign n25012 = n25009 | n25010;
  assign n25013 = ~n25011 & n25012;
  assign n25014 = n24712 & n25013;
  assign n25015 = n24712 | n25013;
  assign n25016 = ~n25014 & n25015;
  assign n25017 = n24711 & n25016;
  assign n25018 = n24711 | n25016;
  assign n25019 = ~n25017 & n25018;
  assign n25020 = n24710 & n25019;
  assign n25021 = n24710 | n25019;
  assign n25022 = ~n25020 & n25021;
  assign n25023 = n24709 | n25022;
  assign n25024 = n24709 & n25022;
  assign n25025 = n25023 & ~n25024;
  assign n25026 = n24702 | n24705;
  assign n25027 = n24701 & n25026;
  assign n25028 = n25025 & ~n25027;
  assign n25029 = ~n25025 & n25027;
  assign n25030 = n25028 | n25029;
  assign n25031 = x117 & x175;
  assign n25032 = n25017 | n25020;
  assign n25033 = x118 & x174;
  assign n25035 = x119 & x173;
  assign n25036 = n25002 | n25006;
  assign n25038 = n24730 & n24973;
  assign n25039 = n24730 | n24973;
  assign n25040 = ~n25038 & n25039;
  assign n32477 = n25038 | n25040;
  assign n32478 = (n24729 & n25038) | (n24729 & n32477) | (n25038 & n32477);
  assign n25043 = n24968 | n24971;
  assign n25045 = x127 & x165;
  assign n25047 = n24924 | n24932;
  assign n32479 = n24759 & n24897;
  assign n36062 = (n24897 & n32307) | (n24897 & n32479) | (n32307 & n32479);
  assign n36063 = (n24579 & n24897) | (n24579 & n32479) | (n24897 & n32479);
  assign n36064 = (n32169 & n36062) | (n32169 & n36063) | (n36062 & n36063);
  assign n36065 = n24759 & n24898;
  assign n36066 = (n24897 & n24898) | (n24897 & n36065) | (n24898 & n36065);
  assign n36067 = (n24898 & n32307) | (n24898 & n36066) | (n32307 & n36066);
  assign n36068 = (n24579 & n24898) | (n24579 & n36066) | (n24898 & n36066);
  assign n36069 = (n32169 & n36067) | (n32169 & n36068) | (n36067 & n36068);
  assign n25051 = ~n36064 & n36069;
  assign n25172 = n24574 | n24769;
  assign n32567 = n25172 | n32192;
  assign n32568 = n24421 | n25172;
  assign n32569 = (n31896 & n32567) | (n31896 & n32568) | (n32567 & n32568);
  assign n25068 = n24797 | n24862;
  assign n32503 = n25068 | n32354;
  assign n32504 = n24531 | n25068;
  assign n32505 = (n32213 & n32503) | (n32213 & n32504) | (n32503 & n32504);
  assign n36074 = n24794 & n32360;
  assign n36075 = n24791 & n24794;
  assign n36076 = (n32053 & n36074) | (n32053 & n36075) | (n36074 & n36075);
  assign n25072 = n36055 & ~n36076;
  assign n25073 = n24525 | n25072;
  assign n25074 = n24862 & n25073;
  assign n32506 = n25070 & n25074;
  assign n32507 = (n25074 & n32213) | (n25074 & n32506) | (n32213 & n32506);
  assign n25076 = n32505 & ~n32507;
  assign n25077 = n24863 & n25076;
  assign n32494 = n24787 & n24869;
  assign n32508 = n25077 | n32494;
  assign n32509 = n24869 | n25077;
  assign n32510 = (n32351 & n32508) | (n32351 & n32509) | (n32508 & n32509);
  assign n32512 = n24802 & n24855;
  assign n36077 = (n24794 & n24855) | (n24794 & n32512) | (n24855 & n32512);
  assign n36078 = (n32360 & n32512) | (n32360 & n36077) | (n32512 & n36077);
  assign n36079 = (n24791 & n32512) | (n24791 & n36077) | (n32512 & n36077);
  assign n36080 = (n32053 & n36078) | (n32053 & n36079) | (n36078 & n36079);
  assign n32514 = n24848 & n36050;
  assign n32515 = n24848 & n32382;
  assign n32516 = (n35950 & n32514) | (n35950 & n32515) | (n32514 & n32515);
  assign n37511 = (n24849 & n24851) | (n24849 & n32382) | (n24851 & n32382);
  assign n37512 = (n24849 & n24851) | (n24849 & n36050) | (n24851 & n36050);
  assign n36083 = (n35950 & n37511) | (n35950 & n37512) | (n37511 & n37512);
  assign n25083 = ~n32516 & n36083;
  assign n32520 = n24841 | n32394;
  assign n36084 = n24815 | n24841;
  assign n36085 = n32375 | n36084;
  assign n36086 = (n32520 & n35951) | (n32520 & n36085) | (n35951 & n36085);
  assign n36087 = (n32262 & n32520) | (n32262 & n36085) | (n32520 & n36085);
  assign n36088 = (n32071 & n36086) | (n32071 & n36087) | (n36086 & n36087);
  assign n25087 = n24495 | n24814;
  assign n25088 = n24841 & n25087;
  assign n32523 = n24509 | n24815;
  assign n32525 = n25088 & n32523;
  assign n36089 = (n25088 & n32525) | (n25088 & n35951) | (n32525 & n35951);
  assign n36090 = (n25088 & n32262) | (n25088 & n32525) | (n32262 & n32525);
  assign n36091 = (n32071 & n36089) | (n32071 & n36090) | (n36089 & n36090);
  assign n25090 = n36088 & ~n36091;
  assign n25091 = n24842 & n25090;
  assign n32398 = n24820 | n32390;
  assign n25099 = x142 & x150;
  assign n32528 = n24485 & n24828;
  assign n36092 = (n24487 & n24828) | (n24487 & n32528) | (n24828 & n32528);
  assign n32538 = n32407 | n36092;
  assign n36093 = n24828 | n32407;
  assign n36094 = (n24485 & n32407) | (n24485 & n36093) | (n32407 & n36093);
  assign n36095 = (n32253 & n32538) | (n32253 & n36094) | (n32538 & n36094);
  assign n36096 = (n32538 & n35966) | (n32538 & n36094) | (n35966 & n36094);
  assign n36097 = (n35760 & n36095) | (n35760 & n36096) | (n36095 & n36096);
  assign n25101 = x143 & x149;
  assign n25102 = n36097 & n25101;
  assign n25103 = n36097 | n25101;
  assign n25104 = ~n25102 & n25103;
  assign n25105 = n25099 & n25104;
  assign n25106 = n25099 | n25104;
  assign n25107 = ~n25105 & n25106;
  assign n36098 = (n32253 & n32528) | (n32253 & n36092) | (n32528 & n36092);
  assign n36099 = (n32528 & n35966) | (n32528 & n36092) | (n35966 & n36092);
  assign n36100 = (n35760 & n36098) | (n35760 & n36099) | (n36098 & n36099);
  assign n32531 = n24485 | n24828;
  assign n36101 = n24487 | n32531;
  assign n32533 = n24823 & n36101;
  assign n36102 = (n24485 & n24823) | (n24485 & n24829) | (n24823 & n24829);
  assign n36103 = (n32253 & n32533) | (n32253 & n36102) | (n32533 & n36102);
  assign n36104 = (n32533 & n35966) | (n32533 & n36102) | (n35966 & n36102);
  assign n36105 = (n35760 & n36103) | (n35760 & n36104) | (n36103 & n36104);
  assign n25097 = ~n36100 & n36105;
  assign n32536 = n24834 | n25097;
  assign n32541 = n25107 | n32536;
  assign n32542 = n25097 | n25107;
  assign n36106 = (n32398 & n32541) | (n32398 & n32542) | (n32541 & n32542);
  assign n32397 = n24820 | n32391;
  assign n36107 = (n32397 & n32541) | (n32397 & n32542) | (n32541 & n32542);
  assign n36108 = (n31943 & n36106) | (n31943 & n36107) | (n36106 & n36107);
  assign n32544 = n25107 & n32536;
  assign n32545 = n25097 & n25107;
  assign n36109 = (n32398 & n32544) | (n32398 & n32545) | (n32544 & n32545);
  assign n36110 = (n32397 & n32544) | (n32397 & n32545) | (n32544 & n32545);
  assign n36111 = (n31943 & n36109) | (n31943 & n36110) | (n36109 & n36110);
  assign n25110 = n36108 & ~n36111;
  assign n25111 = x141 & x151;
  assign n25112 = n25110 | n25111;
  assign n25113 = n25110 & n25111;
  assign n25114 = n25112 & ~n25113;
  assign n37513 = n24820 | n24834;
  assign n37514 = n32390 | n37513;
  assign n37515 = n32391 | n37513;
  assign n36114 = (n31943 & n37514) | (n31943 & n37515) | (n37514 & n37515);
  assign n32547 = ~n24834 & n24835;
  assign n37516 = (~n24820 & n24835) | (~n24820 & n32547) | (n24835 & n32547);
  assign n37518 = (~n32390 & n37516) | (~n32390 & n32547) | (n37516 & n32547);
  assign n37519 = (~n32391 & n37516) | (~n32391 & n32547) | (n37516 & n32547);
  assign n36117 = (~n31943 & n37518) | (~n31943 & n37519) | (n37518 & n37519);
  assign n25117 = n36114 & n36117;
  assign n32549 = n25117 | n32525;
  assign n36118 = ~n25114 & n32549;
  assign n32550 = n25088 | n25117;
  assign n36119 = ~n25114 & n32550;
  assign n36120 = (n32263 & n36118) | (n32263 & n36119) | (n36118 & n36119);
  assign n36121 = n25114 & ~n32549;
  assign n36122 = n25114 & ~n32550;
  assign n36123 = (~n32263 & n36121) | (~n32263 & n36122) | (n36121 & n36122);
  assign n25121 = n36120 | n36123;
  assign n25122 = x140 & x152;
  assign n25123 = n25121 & n25122;
  assign n25124 = n25121 | n25122;
  assign n25125 = ~n25123 & n25124;
  assign n32552 = n25091 | n25125;
  assign n32553 = n32516 | n32552;
  assign n32554 = n25091 & n25125;
  assign n32555 = (n25125 & n32516) | (n25125 & n32554) | (n32516 & n32554);
  assign n25128 = n32553 & ~n32555;
  assign n25129 = x139 & x153;
  assign n25130 = n25128 | n25129;
  assign n25131 = n25128 & n25129;
  assign n25132 = n25130 & ~n25131;
  assign n32556 = n25083 | n25132;
  assign n32557 = n36080 | n32556;
  assign n32558 = n25083 & n25132;
  assign n32559 = (n25132 & n36080) | (n25132 & n32558) | (n36080 & n32558);
  assign n25135 = n32557 & ~n32559;
  assign n25136 = x138 & x154;
  assign n25137 = n25135 | n25136;
  assign n25138 = n25135 & n25136;
  assign n25139 = n25137 & ~n25138;
  assign n32561 = n24802 | n24855;
  assign n36124 = n24794 | n32561;
  assign n36125 = (n32360 & n32561) | (n32360 & n36124) | (n32561 & n36124);
  assign n36126 = (n24791 & n32561) | (n24791 & n36124) | (n32561 & n36124);
  assign n36127 = (n32053 & n36125) | (n32053 & n36126) | (n36125 & n36126);
  assign n25141 = n24856 & ~n36080;
  assign n25142 = n36127 & n25141;
  assign n32563 = ~n25139 & n25142;
  assign n32564 = (~n25139 & n32507) | (~n25139 & n32563) | (n32507 & n32563);
  assign n32565 = n25139 & ~n25142;
  assign n32566 = ~n32507 & n32565;
  assign n25146 = n32564 | n32566;
  assign n25147 = x137 & x155;
  assign n25148 = n25146 & n25147;
  assign n25149 = n25146 | n25147;
  assign n25150 = ~n25148 & n25149;
  assign n25151 = x136 & x156;
  assign n25152 = n25150 & ~n25151;
  assign n25153 = ~n25150 & n25151;
  assign n25154 = n25152 | n25153;
  assign n25155 = n32510 | n25154;
  assign n25156 = n32510 & n25154;
  assign n25157 = n25155 & ~n25156;
  assign n25057 = n24543 | n24781;
  assign n25058 = n24876 & n25057;
  assign n32495 = (n24869 & n32351) | (n24869 & n32494) | (n32351 & n32494);
  assign n36070 = n24787 & n24870;
  assign n36071 = (n24869 & n24870) | (n24869 & n36070) | (n24870 & n36070);
  assign n32499 = (n24870 & n32351) | (n24870 & n36071) | (n32351 & n36071);
  assign n25066 = ~n32495 & n32499;
  assign n32501 = n25058 | n25066;
  assign n36128 = n25157 & ~n32501;
  assign n36072 = n24782 | n25066;
  assign n36073 = (n25058 & n25066) | (n25058 & n36072) | (n25066 & n36072);
  assign n36129 = n25157 & ~n36073;
  assign n36130 = (~n32299 & n36128) | (~n32299 & n36129) | (n36128 & n36129);
  assign n36131 = ~n25157 & n32501;
  assign n36132 = ~n25157 & n36073;
  assign n36133 = (n32299 & n36131) | (n32299 & n36132) | (n36131 & n36132);
  assign n25160 = n36130 | n36133;
  assign n25161 = x135 & x157;
  assign n25162 = n25160 & n25161;
  assign n25163 = n25160 | n25161;
  assign n25164 = ~n25162 & n25163;
  assign n25054 = n24782 | n24876;
  assign n32487 = n24549 | n25054;
  assign n32488 = (n25054 & n32299) | (n25054 & n32487) | (n32299 & n32487);
  assign n32489 = n24782 & n25058;
  assign n32490 = (n25058 & n32299) | (n25058 & n32489) | (n32299 & n32489);
  assign n25060 = n32488 & ~n32490;
  assign n25061 = n24877 & n25060;
  assign n32492 = n24883 | n25061;
  assign n36134 = n25164 | n32492;
  assign n32485 = n24774 & n24883;
  assign n32491 = n25061 | n32485;
  assign n36135 = n25164 | n32491;
  assign n36136 = (n32341 & n36134) | (n32341 & n36135) | (n36134 & n36135);
  assign n36137 = n25164 & n32492;
  assign n36138 = n25164 & n32491;
  assign n36139 = (n32341 & n36137) | (n32341 & n36138) | (n36137 & n36138);
  assign n25167 = n36136 & ~n36139;
  assign n25168 = x134 & x158;
  assign n25169 = n25167 | n25168;
  assign n25170 = n25167 & n25168;
  assign n25171 = n25169 & ~n25170;
  assign n25174 = n32339 & ~n32341;
  assign n25175 = n24561 | n25174;
  assign n25176 = n24890 & n25175;
  assign n32570 = n24774 | n24883;
  assign n32571 = n32341 | n32570;
  assign n32572 = n24884 & ~n32485;
  assign n32573 = (n24885 & ~n32341) | (n24885 & n32572) | (~n32341 & n32572);
  assign n25180 = n32571 & n32573;
  assign n32574 = n25176 | n25180;
  assign n36140 = ~n25171 & n32574;
  assign n36141 = ~n25171 & n25180;
  assign n36142 = (n32569 & n36140) | (n32569 & n36141) | (n36140 & n36141);
  assign n36143 = n25171 & ~n32574;
  assign n36144 = n25171 & ~n25180;
  assign n36145 = (~n32569 & n36143) | (~n32569 & n36144) | (n36143 & n36144);
  assign n25184 = n36142 | n36145;
  assign n32576 = n24890 | n32342;
  assign n32577 = n24769 | n24890;
  assign n32578 = (n32306 & n32576) | (n32306 & n32577) | (n32576 & n32577);
  assign n32579 = n24891 & ~n25176;
  assign n32580 = (n24891 & ~n32569) | (n24891 & n32579) | (~n32569 & n32579);
  assign n25187 = n32578 & n32580;
  assign n25188 = n25184 | n25187;
  assign n32581 = n25188 | n32479;
  assign n32582 = n24897 | n25188;
  assign n32583 = (n32308 & n32581) | (n32308 & n32582) | (n32581 & n32582);
  assign n25177 = n32569 & n25176;
  assign n36146 = n24891 | n32578;
  assign n36147 = (n24891 & ~n25177) | (n24891 & n36146) | (~n25177 & n36146);
  assign n25194 = n25184 & n36147;
  assign n25190 = n24759 | n25187;
  assign n32584 = n25190 & n25194;
  assign n32585 = (n25194 & n32308) | (n25194 & n32584) | (n32308 & n32584);
  assign n25196 = n32583 & ~n32585;
  assign n25197 = x133 & x159;
  assign n25198 = x132 & x160;
  assign n25199 = n25197 & n25198;
  assign n25200 = n25197 | n25198;
  assign n25201 = ~n25199 & n25200;
  assign n25202 = n25196 & n25201;
  assign n25203 = n25196 | n25201;
  assign n25204 = ~n25202 & n25203;
  assign n32586 = ~n25051 & n25204;
  assign n32587 = ~n32468 & n32586;
  assign n32588 = n25051 & ~n25204;
  assign n32589 = (~n25204 & n32468) | (~n25204 & n32588) | (n32468 & n32588);
  assign n25207 = n32587 | n32589;
  assign n25208 = n24915 | n25207;
  assign n32590 = n24916 | n25208;
  assign n32591 = (n25208 & n32472) | (n25208 & n32590) | (n32472 & n32590);
  assign n25212 = n24913 & n25207;
  assign n25210 = n24915 | n24919;
  assign n32592 = n25210 & n25212;
  assign n32593 = (n24599 & n25212) | (n24599 & n32592) | (n25212 & n32592);
  assign n25214 = n32591 & ~n32593;
  assign n25215 = x131 & x161;
  assign n25216 = n25214 & n25215;
  assign n25217 = n25214 | n25215;
  assign n25218 = ~n25216 & n25217;
  assign n25219 = x130 & x162;
  assign n25220 = n25218 & n25219;
  assign n25221 = n25218 | n25219;
  assign n25222 = ~n25220 & n25221;
  assign n25223 = ~n25047 & n25222;
  assign n25224 = n25047 & ~n25222;
  assign n25225 = n25223 | n25224;
  assign n25226 = n24935 | n25225;
  assign n25227 = n24942 | n25226;
  assign n32594 = n24935 | n24940;
  assign n32595 = n24617 | n32594;
  assign n25229 = n24936 & n25225;
  assign n25230 = n32595 & n25229;
  assign n25232 = x129 & x163;
  assign n25233 = x128 & x164;
  assign n25234 = n25232 & ~n25233;
  assign n25235 = ~n25232 & n25233;
  assign n25236 = n25234 | n25235;
  assign n32596 = n25230 | n25236;
  assign n32597 = n25227 & ~n32596;
  assign n32598 = n25230 & n25236;
  assign n32599 = (~n25227 & n25236) | (~n25227 & n32598) | (n25236 & n32598);
  assign n25239 = n32597 | n32599;
  assign n32600 = n24945 | n25239;
  assign n32601 = n24950 | n32600;
  assign n32602 = n24945 & n25239;
  assign n32603 = (n24950 & n25239) | (n24950 & n32602) | (n25239 & n32602);
  assign n25242 = n32601 & ~n32603;
  assign n25243 = n24954 | n25242;
  assign n32604 = n24956 | n25243;
  assign n32605 = (n24748 & n25243) | (n24748 & n32604) | (n25243 & n32604);
  assign n32606 = n24740 | n24954;
  assign n32607 = n24743 | n32606;
  assign n25246 = n24955 & n25242;
  assign n25247 = n32607 & n25246;
  assign n25248 = n32605 & ~n25247;
  assign n25249 = ~n25045 & n25248;
  assign n25250 = n25045 & ~n25248;
  assign n25251 = n25249 | n25250;
  assign n32608 = n24961 & n25251;
  assign n32609 = (n24964 & n25251) | (n24964 & n32608) | (n25251 & n32608);
  assign n32610 = n24961 | n25251;
  assign n32611 = n24964 | n32610;
  assign n25254 = ~n32609 & n32611;
  assign n25255 = x126 & x166;
  assign n25256 = n25254 & n25255;
  assign n25257 = n25254 | n25255;
  assign n25258 = ~n25256 & n25257;
  assign n25259 = n25043 | n25258;
  assign n25260 = n25043 & n25258;
  assign n25261 = n25259 & ~n25260;
  assign n25262 = x125 & x167;
  assign n25263 = x124 & x168;
  assign n25264 = n25262 & n25263;
  assign n25265 = n25262 | n25263;
  assign n25266 = ~n25264 & n25265;
  assign n25267 = n25261 & n25266;
  assign n25268 = n25261 | n25266;
  assign n25269 = ~n25267 & n25268;
  assign n25270 = n32478 | n25269;
  assign n25271 = n32478 & n25269;
  assign n25272 = n25270 & ~n25271;
  assign n25273 = x123 & x169;
  assign n25274 = ~n25272 & n25273;
  assign n25275 = n25272 & ~n25273;
  assign n25276 = n25274 | n25275;
  assign n25278 = n24729 | n25040;
  assign n32612 = n24731 & ~n25040;
  assign n32613 = (~n24729 & n24731) | (~n24729 & n32612) | (n24731 & n32612);
  assign n25280 = n25278 & n32613;
  assign n32614 = n24979 | n25280;
  assign n32615 = (n25280 & n32320) | (n25280 & n32614) | (n32320 & n32614);
  assign n25282 = n25276 & n32615;
  assign n25283 = n25276 | n32615;
  assign n25284 = ~n25282 & n25283;
  assign n25285 = x122 & x170;
  assign n25286 = ~n25284 & n25285;
  assign n25287 = n25284 & ~n25285;
  assign n25288 = n25286 | n25287;
  assign n32616 = n24984 | n24986;
  assign n32617 = (n24718 & n24984) | (n24718 & n32616) | (n24984 & n32616);
  assign n25290 = n25288 & n32617;
  assign n25291 = n25288 | n32617;
  assign n25292 = ~n25290 & n25291;
  assign n25293 = x121 & x171;
  assign n25294 = ~n25292 & n25293;
  assign n25295 = n25292 & ~n25293;
  assign n25296 = n25294 | n25295;
  assign n25297 = n24990 | n24993;
  assign n25298 = n25296 & n25297;
  assign n25299 = n25296 | n25297;
  assign n25300 = ~n25298 & n25299;
  assign n25301 = x120 & x172;
  assign n25302 = ~n25300 & n25301;
  assign n25303 = n25300 & ~n25301;
  assign n25304 = n25302 | n25303;
  assign n32618 = n24996 | n24998;
  assign n32619 = (n24714 & n24996) | (n24714 & n32618) | (n24996 & n32618);
  assign n25306 = n25304 & n32619;
  assign n25307 = n25304 | n32619;
  assign n25308 = ~n25306 & n25307;
  assign n32620 = n25003 & n25308;
  assign n32621 = n25036 & n32620;
  assign n32622 = n25003 | n25308;
  assign n32623 = (n25036 & n25308) | (n25036 & n32622) | (n25308 & n32622);
  assign n25311 = ~n32621 & n32623;
  assign n25312 = ~n25035 & n25311;
  assign n25313 = n25035 & ~n25311;
  assign n25314 = n25312 | n25313;
  assign n32624 = n25011 & n25314;
  assign n32625 = (n25014 & n25314) | (n25014 & n32624) | (n25314 & n32624);
  assign n32626 = n25011 | n25314;
  assign n32627 = n25014 | n32626;
  assign n25317 = ~n32625 & n32627;
  assign n25318 = n25033 & n25317;
  assign n25319 = n25033 | n25317;
  assign n25320 = ~n25318 & n25319;
  assign n25321 = n25032 & n25320;
  assign n25322 = n25032 | n25320;
  assign n25323 = ~n25321 & n25322;
  assign n25324 = n25031 | n25323;
  assign n25325 = n25031 & n25323;
  assign n25326 = n25324 & ~n25325;
  assign n25327 = n25024 | n25027;
  assign n25328 = n25023 & n25327;
  assign n25329 = n25326 & ~n25328;
  assign n25330 = ~n25326 & n25328;
  assign n25331 = n25329 | n25330;
  assign n25332 = x118 & x175;
  assign n32628 = n25318 | n25320;
  assign n32629 = (n25032 & n25318) | (n25032 & n32628) | (n25318 & n32628);
  assign n25334 = x119 & x174;
  assign n25337 = n25300 & n32619;
  assign n32630 = n25300 & n25301;
  assign n32631 = (n25301 & n32619) | (n25301 & n32630) | (n32619 & n32630);
  assign n25340 = ~n25337 & n32631;
  assign n25342 = n25261 & n25262;
  assign n25343 = n25261 | n25262;
  assign n25344 = ~n25342 & n25343;
  assign n25345 = n32478 & n25344;
  assign n25346 = n25342 | n25345;
  assign n32632 = n25256 | n25258;
  assign n32633 = (n25043 & n25256) | (n25043 & n32632) | (n25256 & n32632);
  assign n25348 = x127 & x166;
  assign n25349 = n25045 & n25248;
  assign n32634 = ~n25230 & n25232;
  assign n32635 = n25227 & n32634;
  assign n32636 = n25230 & ~n25232;
  assign n32637 = (n25227 & n25232) | (n25227 & ~n32636) | (n25232 & ~n32636);
  assign n25352 = ~n32635 & n32637;
  assign n32638 = n24945 | n25352;
  assign n32639 = n24950 | n32638;
  assign n32640 = n24945 & n25352;
  assign n32641 = (n24950 & n25352) | (n24950 & n32640) | (n25352 & n32640);
  assign n25355 = n25233 & ~n32641;
  assign n25356 = n32639 & n25355;
  assign n32642 = n25246 | n25356;
  assign n32643 = (n25356 & n32607) | (n25356 & n32642) | (n32607 & n32642);
  assign n25358 = n32635 | n32641;
  assign n25686 = n24924 | n25216;
  assign n36148 = (n25216 & n25218) | (n25216 & n25686) | (n25218 & n25686);
  assign n32651 = n25216 | n25218;
  assign n32652 = (n24932 & n36148) | (n24932 & n32651) | (n36148 & n32651);
  assign n25365 = x131 & x162;
  assign n25366 = x132 & x161;
  assign n25367 = n25196 | n25197;
  assign n36149 = n25197 & ~n32584;
  assign n36150 = ~n25194 & n25197;
  assign n36151 = (~n32308 & n36149) | (~n32308 & n36150) | (n36149 & n36150);
  assign n25369 = n32583 & n36151;
  assign n25370 = n25367 & ~n25369;
  assign n36152 = n25051 & ~n25369;
  assign n36153 = n25367 & n36152;
  assign n32654 = (n25370 & n32468) | (n25370 & n36153) | (n32468 & n36153);
  assign n32658 = n25167 & n25180;
  assign n36154 = (n25167 & n25176) | (n25167 & n32658) | (n25176 & n32658);
  assign n32659 = (n32569 & n36154) | (n32569 & n32658) | (n36154 & n32658);
  assign n32661 = n25167 | n25180;
  assign n36155 = n25176 | n32661;
  assign n36156 = n25168 & n36155;
  assign n36157 = n25168 & n32661;
  assign n36158 = (n32569 & n36156) | (n32569 & n36157) | (n36156 & n36157);
  assign n25380 = ~n32659 & n36158;
  assign n36159 = n24883 | n25160;
  assign n36160 = n25061 | n36159;
  assign n32664 = n25160 | n32491;
  assign n32665 = (n32341 & n36160) | (n32341 & n32664) | (n36160 & n32664);
  assign n25385 = n24877 | n25060;
  assign n25386 = n25160 & n25385;
  assign n25383 = n24774 | n25061;
  assign n32666 = n25383 & n25386;
  assign n32667 = (n25386 & n32341) | (n25386 & n32666) | (n32341 & n32666);
  assign n25388 = n32665 & ~n32667;
  assign n25389 = n25161 & n25388;
  assign n32764 = n25389 | n32574;
  assign n32765 = n25180 | n25389;
  assign n32766 = (n32569 & n32764) | (n32569 & n32765) | (n32764 & n32765);
  assign n32502 = (n32299 & n36073) | (n32299 & n32501) | (n36073 & n32501);
  assign n32679 = n25091 | n36050;
  assign n32680 = n25091 | n32382;
  assign n32681 = (n35950 & n32679) | (n35950 & n32680) | (n32679 & n32680);
  assign n25412 = x142 & x151;
  assign n25415 = x143 & x150;
  assign n36163 = n25097 | n25102;
  assign n36164 = (n25102 & n25104) | (n25102 & n36163) | (n25104 & n36163);
  assign n32692 = n25415 & n36164;
  assign n32685 = n25104 & n32536;
  assign n37520 = n25101 & n25415;
  assign n37521 = n36097 & n37520;
  assign n36162 = (n25415 & n32685) | (n25415 & n37521) | (n32685 & n37521);
  assign n36165 = (n32398 & n32692) | (n32398 & n36162) | (n32692 & n36162);
  assign n36166 = (n32397 & n32692) | (n32397 & n36162) | (n32692 & n36162);
  assign n36167 = (n31943 & n36165) | (n31943 & n36166) | (n36165 & n36166);
  assign n32695 = n25415 | n36164;
  assign n37522 = n25101 | n25415;
  assign n37523 = (n25415 & n36097) | (n25415 & n37522) | (n36097 & n37522);
  assign n36169 = n32685 | n37523;
  assign n36170 = (n32398 & n32695) | (n32398 & n36169) | (n32695 & n36169);
  assign n36171 = (n32397 & n32695) | (n32397 & n36169) | (n32695 & n36169);
  assign n36172 = (n31943 & n36170) | (n31943 & n36171) | (n36170 & n36171);
  assign n25418 = ~n36167 & n36172;
  assign n25419 = n25412 & n25418;
  assign n25420 = n25412 | n25418;
  assign n25421 = ~n25419 & n25420;
  assign n32697 = n25104 | n32536;
  assign n32698 = n25097 | n25104;
  assign n37524 = (n24820 & n32697) | (n24820 & n32698) | (n32697 & n32698);
  assign n37525 = n32697 | n32698;
  assign n37526 = (n32390 & n37524) | (n32390 & n37525) | (n37524 & n37525);
  assign n37527 = (n32391 & n37524) | (n32391 & n37525) | (n37524 & n37525);
  assign n36175 = (n31943 & n37526) | (n31943 & n37527) | (n37526 & n37527);
  assign n32701 = n25099 & ~n32685;
  assign n36176 = ~n25097 & n25099;
  assign n36177 = (n25099 & ~n25104) | (n25099 & n36176) | (~n25104 & n36176);
  assign n36178 = (~n32398 & n32701) | (~n32398 & n36177) | (n32701 & n36177);
  assign n36179 = (~n32397 & n32701) | (~n32397 & n36177) | (n32701 & n36177);
  assign n36180 = (~n31943 & n36178) | (~n31943 & n36179) | (n36178 & n36179);
  assign n25425 = n36175 & n36180;
  assign n32703 = n25110 | n25425;
  assign n32705 = n25421 | n32703;
  assign n32706 = n25421 | n25425;
  assign n36181 = (n32549 & n32705) | (n32549 & n32706) | (n32705 & n32706);
  assign n36182 = (n32550 & n32705) | (n32550 & n32706) | (n32705 & n32706);
  assign n36183 = (n32263 & n36181) | (n32263 & n36182) | (n36181 & n36182);
  assign n32708 = n25421 & n32703;
  assign n32709 = n25421 & n25425;
  assign n36184 = (n32549 & n32708) | (n32549 & n32709) | (n32708 & n32709);
  assign n36185 = (n32550 & n32708) | (n32550 & n32709) | (n32708 & n32709);
  assign n36186 = (n32263 & n36184) | (n32263 & n36185) | (n36184 & n36185);
  assign n25429 = n36183 & ~n36186;
  assign n25430 = x141 & x152;
  assign n25431 = n25429 | n25430;
  assign n25432 = n25429 & n25430;
  assign n25433 = n25431 & ~n25432;
  assign n25406 = n24842 | n25090;
  assign n25407 = n25121 & n25406;
  assign n37528 = n25110 | n25117;
  assign n37529 = n32525 | n37528;
  assign n37530 = n25088 | n37528;
  assign n36189 = (n32263 & n37529) | (n32263 & n37530) | (n37529 & n37530);
  assign n32711 = ~n25110 & n25111;
  assign n37531 = (n25111 & ~n25117) | (n25111 & n32711) | (~n25117 & n32711);
  assign n37533 = (~n32525 & n37531) | (~n32525 & n32711) | (n37531 & n32711);
  assign n36191 = (n25111 & ~n32550) | (n25111 & n32711) | (~n32550 & n32711);
  assign n36192 = (~n32263 & n37533) | (~n32263 & n36191) | (n37533 & n36191);
  assign n25436 = n36189 & n36192;
  assign n32713 = n25407 | n25436;
  assign n32715 = ~n25433 & n32713;
  assign n32716 = ~n25433 & n25436;
  assign n32717 = (n32681 & n32715) | (n32681 & n32716) | (n32715 & n32716);
  assign n32718 = n25433 & ~n32713;
  assign n32719 = n25433 & ~n25436;
  assign n32720 = (~n32681 & n32718) | (~n32681 & n32719) | (n32718 & n32719);
  assign n25440 = n32717 | n32720;
  assign n25441 = x140 & x153;
  assign n25442 = n25440 & n25441;
  assign n25443 = n25440 | n25441;
  assign n25444 = ~n25442 & n25443;
  assign n32677 = n25091 | n25121;
  assign n36193 = n32515 | n32677;
  assign n36194 = n32514 | n32677;
  assign n36195 = (n35950 & n36193) | (n35950 & n36194) | (n36193 & n36194);
  assign n36196 = n25407 & n32680;
  assign n36197 = n25407 & n32679;
  assign n36198 = (n35950 & n36196) | (n35950 & n36197) | (n36196 & n36197);
  assign n25409 = n36195 & ~n36198;
  assign n25410 = n25122 & n25409;
  assign n32683 = n25128 | n25410;
  assign n32721 = n25444 | n32683;
  assign n32675 = n25083 & n25128;
  assign n32682 = n25410 | n32675;
  assign n32722 = n25444 | n32682;
  assign n32723 = (n36080 & n32721) | (n36080 & n32722) | (n32721 & n32722);
  assign n32724 = n25444 & n32683;
  assign n32725 = n25444 & n32682;
  assign n32726 = (n36080 & n32724) | (n36080 & n32725) | (n32724 & n32725);
  assign n25447 = n32723 & ~n32726;
  assign n25448 = x139 & x154;
  assign n25449 = n25447 | n25448;
  assign n25450 = n25447 & n25448;
  assign n25451 = n25449 & ~n25450;
  assign n32729 = n25083 | n25128;
  assign n32730 = n36080 | n32729;
  assign n36199 = ~n25083 & n25129;
  assign n36200 = (~n25128 & n25129) | (~n25128 & n36199) | (n25129 & n36199);
  assign n32732 = ~n25128 & n25129;
  assign n32733 = (~n36080 & n36200) | (~n36080 & n32732) | (n36200 & n32732);
  assign n25455 = n32730 & n32733;
  assign n32727 = n25135 & n25142;
  assign n32734 = n25455 | n32727;
  assign n32737 = n25451 | n32734;
  assign n32735 = n25135 | n25455;
  assign n32738 = n25451 | n32735;
  assign n32739 = (n32507 & n32737) | (n32507 & n32738) | (n32737 & n32738);
  assign n32740 = n25451 & n32734;
  assign n32741 = n25451 & n32735;
  assign n32742 = (n32507 & n32740) | (n32507 & n32741) | (n32740 & n32741);
  assign n25459 = n32739 & ~n32742;
  assign n25460 = x138 & x155;
  assign n25461 = n25459 | n25460;
  assign n25462 = n25459 & n25460;
  assign n25463 = n25461 & ~n25462;
  assign n25397 = n24863 | n25076;
  assign n25398 = n25146 & n25397;
  assign n36201 = n24787 | n24863;
  assign n36202 = (n24787 & n25076) | (n24787 & n36201) | (n25076 & n36201);
  assign n32671 = n36202 & n25398;
  assign n32672 = (n25398 & n32351) | (n25398 & n32671) | (n32351 & n32671);
  assign n32743 = n25135 | n25142;
  assign n36203 = n32506 | n32743;
  assign n36204 = n25074 | n32743;
  assign n36205 = (n32213 & n36203) | (n32213 & n36204) | (n36203 & n36204);
  assign n32745 = n25136 & ~n32727;
  assign n32746 = ~n25135 & n25136;
  assign n36206 = (~n32506 & n32745) | (~n32506 & n32746) | (n32745 & n32746);
  assign n36207 = (~n25074 & n32745) | (~n25074 & n32746) | (n32745 & n32746);
  assign n36208 = (~n32213 & n36206) | (~n32213 & n36207) | (n36206 & n36207);
  assign n25466 = n36205 & n36208;
  assign n32748 = ~n25463 & n25466;
  assign n32749 = (~n25463 & n32672) | (~n25463 & n32748) | (n32672 & n32748);
  assign n32750 = n25463 & ~n25466;
  assign n32751 = ~n32672 & n32750;
  assign n25470 = n32749 | n32751;
  assign n25471 = x137 & x156;
  assign n25472 = n25470 & n25471;
  assign n25473 = n25470 | n25471;
  assign n25474 = ~n25472 & n25473;
  assign n25390 = n32510 | n25150;
  assign n25391 = n32510 & n25150;
  assign n25392 = n25390 & ~n25391;
  assign n32668 = n25146 | n32509;
  assign n32669 = n25146 | n32508;
  assign n32670 = (n32351 & n32668) | (n32351 & n32669) | (n32668 & n32669);
  assign n25400 = n32670 & ~n32672;
  assign n25401 = n25147 & n25400;
  assign n32673 = n25392 | n25401;
  assign n32752 = n25474 | n32673;
  assign n32753 = n25401 | n25474;
  assign n32754 = (n32502 & n32752) | (n32502 & n32753) | (n32752 & n32753);
  assign n32755 = n25474 & n32673;
  assign n32756 = n25401 & n25474;
  assign n32757 = (n32502 & n32755) | (n32502 & n32756) | (n32755 & n32756);
  assign n25477 = n32754 & ~n32757;
  assign n25478 = x136 & x157;
  assign n25479 = n25477 | n25478;
  assign n25480 = n25477 & n25478;
  assign n25481 = n25479 & ~n25480;
  assign n36209 = n25392 | n32501;
  assign n36210 = n25392 | n36073;
  assign n36211 = (n32299 & n36209) | (n32299 & n36210) | (n36209 & n36210);
  assign n32758 = n25151 & ~n25392;
  assign n36212 = (n25151 & ~n32501) | (n25151 & n32758) | (~n32501 & n32758);
  assign n36213 = (n25151 & n32758) | (n25151 & ~n36073) | (n32758 & ~n36073);
  assign n36214 = (~n32299 & n36212) | (~n32299 & n36213) | (n36212 & n36213);
  assign n25484 = n36211 & n36214;
  assign n32760 = ~n25481 & n25484;
  assign n32761 = (~n25481 & n32667) | (~n25481 & n32760) | (n32667 & n32760);
  assign n32762 = n25481 & ~n25484;
  assign n32763 = ~n32667 & n32762;
  assign n25488 = n32761 | n32763;
  assign n25492 = n25161 | n25388;
  assign n25493 = n25488 & n25492;
  assign n25494 = n32766 & n25493;
  assign n25496 = x135 & x158;
  assign n25497 = x134 & x159;
  assign n25498 = n25496 & n25497;
  assign n25499 = n25496 | n25497;
  assign n25500 = ~n25498 & n25499;
  assign n25489 = n25389 | n25488;
  assign n36215 = n25489 | n36154;
  assign n36216 = n25489 | n32658;
  assign n36217 = (n32569 & n36215) | (n32569 & n36216) | (n36215 & n36216);
  assign n36218 = n25500 & n36217;
  assign n36219 = ~n25494 & n36218;
  assign n36220 = n25500 | n36217;
  assign n36221 = (~n25494 & n25500) | (~n25494 & n36220) | (n25500 & n36220);
  assign n25503 = ~n36219 & n36221;
  assign n32767 = ~n25380 & n25503;
  assign n32768 = ~n32585 & n32767;
  assign n32769 = n25380 & ~n25503;
  assign n32770 = (~n25503 & n32585) | (~n25503 & n32769) | (n32585 & n32769);
  assign n25506 = n32768 | n32770;
  assign n25507 = x133 & x160;
  assign n25508 = n25506 & n25507;
  assign n25509 = n25506 | n25507;
  assign n25510 = ~n25508 & n25509;
  assign n32771 = n25369 | n25510;
  assign n32772 = n32654 | n32771;
  assign n32773 = n25369 & n25510;
  assign n32774 = (n25510 & n32654) | (n25510 & n32773) | (n32654 & n32773);
  assign n25513 = n32772 & ~n32774;
  assign n36222 = ~n25051 & n25369;
  assign n36223 = (n25051 & n25367) | (n25051 & ~n36222) | (n25367 & ~n36222);
  assign n36224 = n25198 & n36223;
  assign n36225 = (n25198 & n32468) | (n25198 & n36224) | (n32468 & n36224);
  assign n25374 = ~n32654 & n36225;
  assign n32775 = n25374 & n25513;
  assign n32776 = (n25513 & n32593) | (n25513 & n32775) | (n32593 & n32775);
  assign n32777 = n25374 | n25513;
  assign n32778 = n32593 | n32777;
  assign n25516 = ~n32776 & n32778;
  assign n25517 = n25366 & n25516;
  assign n25518 = n25366 | n25516;
  assign n25519 = ~n25517 & n25518;
  assign n25520 = n25365 & n25519;
  assign n25521 = n25365 | n25519;
  assign n25522 = ~n25520 & n25521;
  assign n25523 = n32652 | n25522;
  assign n25524 = n32652 & n25522;
  assign n25525 = n25523 & ~n25524;
  assign n32644 = n24924 & n25218;
  assign n32645 = (n24932 & n25218) | (n24932 & n32644) | (n25218 & n32644);
  assign n37534 = n24751 & n25219;
  assign n37535 = n24923 & n37534;
  assign n36227 = (n25218 & n25219) | (n25218 & n37535) | (n25219 & n37535);
  assign n32649 = (n24932 & n25219) | (n24932 & n36227) | (n25219 & n36227);
  assign n25362 = ~n32645 & n32649;
  assign n32779 = n25362 & n25525;
  assign n32780 = (n25230 & n25525) | (n25230 & n32779) | (n25525 & n32779);
  assign n32781 = n25362 | n25525;
  assign n32782 = n25230 | n32781;
  assign n25528 = ~n32780 & n32782;
  assign n25529 = x130 & x163;
  assign n25530 = n25528 & n25529;
  assign n25531 = n25528 | n25529;
  assign n25532 = ~n25530 & n25531;
  assign n25533 = x129 & x164;
  assign n25534 = n25532 & n25533;
  assign n25535 = n25532 | n25533;
  assign n25536 = ~n25534 & n25535;
  assign n25537 = n25358 | n25536;
  assign n25538 = n25358 & n25536;
  assign n25539 = n25537 & ~n25538;
  assign n25540 = x128 & x165;
  assign n25541 = ~n25539 & n25540;
  assign n25542 = n25539 & ~n25540;
  assign n25543 = n25541 | n25542;
  assign n25544 = n32643 | n25543;
  assign n25545 = n32643 & n25543;
  assign n25546 = n25544 & ~n25545;
  assign n25547 = n25349 | n25546;
  assign n25548 = n32609 | n25547;
  assign n32783 = n24961 | n25349;
  assign n32784 = n24964 | n32783;
  assign n25550 = n25045 | n25248;
  assign n25551 = n25546 & n25550;
  assign n25552 = n32784 & n25551;
  assign n25553 = n25548 & ~n25552;
  assign n25554 = ~n25348 & n25553;
  assign n25555 = n25348 & ~n25553;
  assign n25556 = n25554 | n25555;
  assign n25557 = n32633 | n25556;
  assign n25558 = n32633 & n25556;
  assign n25559 = n25557 & ~n25558;
  assign n25560 = x126 & x167;
  assign n25561 = x125 & x168;
  assign n25562 = n25560 & n25561;
  assign n25563 = n25560 | n25561;
  assign n25564 = ~n25562 & n25563;
  assign n25565 = n25559 & n25564;
  assign n25566 = n25559 | n25564;
  assign n25567 = ~n25565 & n25566;
  assign n25568 = n25346 | n25567;
  assign n25569 = n25346 & n25567;
  assign n25570 = n25568 & ~n25569;
  assign n25571 = x124 & x169;
  assign n25572 = ~n25570 & n25571;
  assign n25573 = n25570 & ~n25571;
  assign n25574 = n25572 | n25573;
  assign n25575 = n25272 & n32615;
  assign n25576 = n32478 | n25344;
  assign n25577 = n25263 & ~n25345;
  assign n25578 = n25576 & n25577;
  assign n25579 = n25575 | n25578;
  assign n25580 = n25574 & n25579;
  assign n25581 = n25574 | n25579;
  assign n25582 = ~n25580 & n25581;
  assign n25583 = x123 & x170;
  assign n25584 = ~n25582 & n25583;
  assign n25585 = n25582 & ~n25583;
  assign n25586 = n25584 | n25585;
  assign n25588 = n25272 | n32615;
  assign n32785 = (n25273 & n25274) | (n25273 & ~n32615) | (n25274 & ~n32615);
  assign n25590 = n25588 & n32785;
  assign n32786 = n25284 | n25590;
  assign n32787 = (n25590 & n32617) | (n25590 & n32786) | (n32617 & n32786);
  assign n25592 = n25586 & n32787;
  assign n25593 = n25586 | n32787;
  assign n25594 = ~n25592 & n25593;
  assign n25595 = x122 & x171;
  assign n25596 = ~n25594 & n25595;
  assign n25597 = n25594 & ~n25595;
  assign n25598 = n25596 | n25597;
  assign n25600 = n25284 | n32617;
  assign n32790 = (n25285 & n25286) | (n25285 & ~n32617) | (n25286 & ~n32617);
  assign n25602 = n25600 & n32790;
  assign n32788 = n24990 & n25292;
  assign n32791 = n25602 | n32788;
  assign n32792 = n25292 | n25602;
  assign n32793 = (n24993 & n32791) | (n24993 & n32792) | (n32791 & n32792);
  assign n25604 = n25598 & n32793;
  assign n25605 = n25598 | n32793;
  assign n25606 = ~n25604 & n25605;
  assign n25607 = x121 & x172;
  assign n25608 = ~n25606 & n25607;
  assign n25609 = n25606 & ~n25607;
  assign n25610 = n25608 | n25609;
  assign n32794 = n24990 | n25292;
  assign n32795 = n24993 | n32794;
  assign n32796 = n25293 & ~n32788;
  assign n32797 = (~n24993 & n25294) | (~n24993 & n32796) | (n25294 & n32796);
  assign n25613 = n32795 & n32797;
  assign n32798 = n25300 | n25613;
  assign n32799 = (n25613 & n32619) | (n25613 & n32798) | (n32619 & n32798);
  assign n25615 = n25610 & n32799;
  assign n25616 = n25610 | n32799;
  assign n25617 = ~n25615 & n25616;
  assign n32800 = ~n25340 & n25617;
  assign n32801 = ~n32621 & n32800;
  assign n32802 = n25340 & ~n25617;
  assign n32803 = (~n25617 & n32621) | (~n25617 & n32802) | (n32621 & n32802);
  assign n25620 = n32801 | n32803;
  assign n25621 = x120 & x173;
  assign n25622 = n25620 & n25621;
  assign n25623 = n25620 | n25621;
  assign n25624 = ~n25622 & n25623;
  assign n25335 = n25035 & n25311;
  assign n32804 = n25335 & n25624;
  assign n32805 = (n25624 & n32625) | (n25624 & n32804) | (n32625 & n32804);
  assign n32806 = n25335 | n25624;
  assign n32807 = n32625 | n32806;
  assign n25627 = ~n32805 & n32807;
  assign n25628 = n25334 & n25627;
  assign n25629 = n25334 | n25627;
  assign n25630 = ~n25628 & n25629;
  assign n25631 = n32629 & n25630;
  assign n25632 = n32629 | n25630;
  assign n25633 = ~n25631 & n25632;
  assign n25634 = n25332 | n25633;
  assign n25635 = n25332 & n25633;
  assign n25636 = n25634 & ~n25635;
  assign n25637 = n25325 | n25328;
  assign n25638 = n25324 & n25637;
  assign n25639 = n25636 & ~n25638;
  assign n25640 = ~n25636 & n25638;
  assign n25641 = n25639 | n25640;
  assign n25642 = x119 & x175;
  assign n32808 = n25628 | n25630;
  assign n32809 = (n25628 & n32629) | (n25628 & n32808) | (n32629 & n32808);
  assign n25644 = x120 & x174;
  assign n32810 = n25340 & n25617;
  assign n32811 = (n25617 & n32621) | (n25617 & n32810) | (n32621 & n32810);
  assign n32812 = n25606 & n32798;
  assign n32813 = n25606 & n25613;
  assign n32814 = (n32619 & n32812) | (n32619 & n32813) | (n32812 & n32813);
  assign n32815 = n25606 | n32798;
  assign n32816 = n25606 | n25613;
  assign n32817 = (n32619 & n32815) | (n32619 & n32816) | (n32815 & n32816);
  assign n25649 = n25607 & n32817;
  assign n25650 = ~n32814 & n25649;
  assign n25652 = n25559 & n25560;
  assign n25653 = n25559 | n25560;
  assign n25654 = ~n25652 & n25653;
  assign n32818 = n25652 | n25654;
  assign n32819 = (n25346 & n25652) | (n25346 & n32818) | (n25652 & n32818);
  assign n25657 = n25348 & n25553;
  assign n32820 = n25556 | n25657;
  assign n32821 = (n25657 & n32633) | (n25657 & n32820) | (n32633 & n32820);
  assign n25659 = x126 & x168;
  assign n25660 = ~n32821 & n25659;
  assign n25661 = n32821 & ~n25659;
  assign n25662 = n25660 | n25661;
  assign n25668 = n32635 | n25532;
  assign n25669 = n32641 | n25668;
  assign n25670 = n24945 | n32635;
  assign n25671 = n24950 | n25670;
  assign n25363 = n25230 | n25362;
  assign n25672 = ~n25525 & n25529;
  assign n25673 = n25525 & ~n25529;
  assign n25674 = n25672 | n25673;
  assign n25675 = ~n25363 & n25674;
  assign n25676 = n25363 & ~n25674;
  assign n25677 = n25675 | n25676;
  assign n36230 = n25533 & ~n32637;
  assign n36231 = (n25533 & ~n25677) | (n25533 & n36230) | (~n25677 & n36230);
  assign n32827 = (n25533 & ~n25671) | (n25533 & n36231) | (~n25671 & n36231);
  assign n25681 = n25669 & n32827;
  assign n32828 = n25539 | n25681;
  assign n32829 = (n25681 & n32643) | (n25681 & n32828) | (n32643 & n32828);
  assign n25678 = n32637 & n25677;
  assign n32830 = n25530 | n25678;
  assign n32831 = (n25530 & n25671) | (n25530 & n32830) | (n25671 & n32830);
  assign n25684 = n25216 | n25519;
  assign n25685 = n32645 | n25684;
  assign n25687 = n24932 | n25686;
  assign n25688 = n25217 & n25519;
  assign n25689 = n25687 & n25688;
  assign n25690 = n25685 & ~n25689;
  assign n25691 = n25365 & n25690;
  assign n32832 = n25691 | n32779;
  assign n32833 = n25525 | n25691;
  assign n32834 = (n25230 & n32832) | (n25230 & n32833) | (n32832 & n32833);
  assign n25693 = x131 & x163;
  assign n36232 = n25217 | n25517;
  assign n36233 = (n25517 & n25519) | (n25517 & n36232) | (n25519 & n36232);
  assign n32836 = (n25517 & n25687) | (n25517 & n36233) | (n25687 & n36233);
  assign n25695 = x132 & x162;
  assign n25696 = x133 & x161;
  assign n32839 = n25369 | n25506;
  assign n36234 = n32839 | n36153;
  assign n36235 = n25370 | n32839;
  assign n36236 = (n32468 & n36234) | (n32468 & n36235) | (n36234 & n36235);
  assign n25699 = n25367 & n25506;
  assign n25697 = n25051 | n25369;
  assign n32837 = n25697 & n25699;
  assign n32838 = (n25699 & n32468) | (n25699 & n32837) | (n32468 & n32837);
  assign n32841 = n25507 & ~n32838;
  assign n32842 = n36236 & n32841;
  assign n32843 = n32775 | n32842;
  assign n32844 = n25513 | n32842;
  assign n32845 = (n32593 & n32843) | (n32593 & n32844) | (n32843 & n32844);
  assign n36237 = n25496 & n36217;
  assign n36238 = ~n25494 & n36237;
  assign n36239 = n25496 | n36217;
  assign n36240 = (~n25494 & n25496) | (~n25494 & n36239) | (n25496 & n36239);
  assign n25707 = ~n36238 & n36240;
  assign n32846 = n25380 & n25707;
  assign n32847 = (n25707 & n32585) | (n25707 & n32846) | (n32585 & n32846);
  assign n37536 = n25380 & n25497;
  assign n37537 = (n25497 & n25707) | (n25497 & n37536) | (n25707 & n37536);
  assign n36242 = (n25497 & n32585) | (n25497 & n37537) | (n32585 & n37537);
  assign n25711 = ~n32847 & n36242;
  assign n25712 = n32838 | n25711;
  assign n32858 = n25470 | n32673;
  assign n32859 = n25401 | n25470;
  assign n32860 = (n32502 & n32858) | (n32502 & n32859) | (n32858 & n32859);
  assign n25721 = n25147 | n25400;
  assign n25722 = n25470 & n25721;
  assign n32861 = n25401 & n25722;
  assign n32862 = (n25722 & n32502) | (n25722 & n32861) | (n32502 & n32861);
  assign n25724 = n32860 & ~n32862;
  assign n25727 = n25471 | n25724;
  assign n32875 = n25447 & n32735;
  assign n36247 = n25447 & n25455;
  assign n36248 = (n25447 & n32727) | (n25447 & n36247) | (n32727 & n36247);
  assign n36249 = (n32506 & n32875) | (n32506 & n36248) | (n32875 & n36248);
  assign n36250 = (n25074 & n32875) | (n25074 & n36248) | (n32875 & n36248);
  assign n36251 = (n32213 & n36249) | (n32213 & n36250) | (n36249 & n36250);
  assign n32883 = n25440 | n32683;
  assign n36257 = n25410 | n25440;
  assign n36258 = n32675 | n36257;
  assign n32885 = (n36080 & n32883) | (n36080 & n36258) | (n32883 & n36258);
  assign n25740 = n25122 | n25409;
  assign n25741 = n25440 & n25740;
  assign n32886 = n25083 | n25410;
  assign n32888 = n25741 & n32886;
  assign n36259 = n25441 & ~n32888;
  assign n36260 = n25441 & ~n25741;
  assign n36261 = (~n36080 & n36259) | (~n36080 & n36260) | (n36259 & n36260);
  assign n25744 = n32885 & n36261;
  assign n32889 = (n25741 & n36080) | (n25741 & n32888) | (n36080 & n32888);
  assign n32891 = n25429 & n25436;
  assign n36262 = (n25407 & n25429) | (n25407 & n32891) | (n25429 & n32891);
  assign n36263 = (n32680 & n32891) | (n32680 & n36262) | (n32891 & n36262);
  assign n36264 = (n32679 & n32891) | (n32679 & n36262) | (n32891 & n36262);
  assign n36265 = (n35950 & n36263) | (n35950 & n36264) | (n36263 & n36264);
  assign n32894 = n25429 | n25436;
  assign n36266 = n25407 | n32894;
  assign n36267 = (n32680 & n32894) | (n32680 & n36266) | (n32894 & n36266);
  assign n36268 = (n32679 & n32894) | (n32679 & n36266) | (n32894 & n36266);
  assign n36269 = (n35950 & n36267) | (n35950 & n36268) | (n36267 & n36268);
  assign n25748 = n25430 & n36269;
  assign n25749 = ~n36265 & n25748;
  assign n32896 = n25418 & n32703;
  assign n32897 = n25418 & n25425;
  assign n36270 = (n32549 & n32896) | (n32549 & n32897) | (n32896 & n32897);
  assign n36271 = (n32550 & n32896) | (n32550 & n32897) | (n32896 & n32897);
  assign n36272 = (n32263 & n36270) | (n32263 & n36271) | (n36270 & n36271);
  assign n32900 = n25418 | n25425;
  assign n32903 = n25412 & n32900;
  assign n36273 = (n25412 & n25419) | (n25412 & n32703) | (n25419 & n32703);
  assign n36274 = (n32549 & n32903) | (n32549 & n36273) | (n32903 & n36273);
  assign n36275 = (n32550 & n32903) | (n32550 & n36273) | (n32903 & n36273);
  assign n36276 = (n32263 & n36274) | (n32263 & n36275) | (n36274 & n36275);
  assign n25754 = ~n36272 & n36276;
  assign n25756 = x142 & x152;
  assign n25758 = x143 & x151;
  assign n36277 = n25418 | n36167;
  assign n36278 = (n32703 & n36167) | (n32703 & n36277) | (n36167 & n36277);
  assign n32908 = n25758 & n36278;
  assign n36279 = n25758 & n36167;
  assign n36280 = (n25758 & n32897) | (n25758 & n36279) | (n32897 & n36279);
  assign n36281 = (n32549 & n32908) | (n32549 & n36280) | (n32908 & n36280);
  assign n36282 = (n32550 & n32908) | (n32550 & n36280) | (n32908 & n36280);
  assign n36283 = (n32263 & n36281) | (n32263 & n36282) | (n36281 & n36282);
  assign n32911 = n25758 | n36278;
  assign n36284 = n25758 | n36167;
  assign n36285 = n32897 | n36284;
  assign n36286 = (n32549 & n32911) | (n32549 & n36285) | (n32911 & n36285);
  assign n36287 = (n32550 & n32911) | (n32550 & n36285) | (n32911 & n36285);
  assign n36288 = (n32263 & n36286) | (n32263 & n36287) | (n36286 & n36287);
  assign n25761 = ~n36283 & n36288;
  assign n25762 = n25756 & n25761;
  assign n25763 = n25756 | n25761;
  assign n25764 = ~n25762 & n25763;
  assign n32914 = n25754 | n25764;
  assign n32915 = n36265 | n32914;
  assign n32916 = n25754 & n25764;
  assign n32917 = (n25764 & n36265) | (n25764 & n32916) | (n36265 & n32916);
  assign n25767 = n32915 & ~n32917;
  assign n25768 = x141 & x153;
  assign n25769 = n25767 | n25768;
  assign n25770 = n25767 & n25768;
  assign n25771 = n25769 & ~n25770;
  assign n32918 = n25749 | n25771;
  assign n32919 = n32889 | n32918;
  assign n32920 = n25749 & n25771;
  assign n32921 = (n25771 & n32889) | (n25771 & n32920) | (n32889 & n32920);
  assign n25774 = n32919 & ~n32921;
  assign n25775 = x140 & x154;
  assign n25776 = n25774 | n25775;
  assign n25777 = n25774 & n25775;
  assign n25778 = n25776 & ~n25777;
  assign n32922 = n25744 | n25778;
  assign n32923 = n36251 | n32922;
  assign n32924 = n25744 & n25778;
  assign n32925 = (n25778 & n36251) | (n25778 & n32924) | (n36251 & n32924);
  assign n25781 = n32923 & ~n32925;
  assign n25782 = x139 & x155;
  assign n25783 = n25781 | n25782;
  assign n25784 = n25781 & n25782;
  assign n25785 = n25783 & ~n25784;
  assign n32878 = n25447 | n32735;
  assign n36252 = n25447 | n25455;
  assign n36253 = n32727 | n36252;
  assign n36254 = (n32506 & n32878) | (n32506 & n36253) | (n32878 & n36253);
  assign n36255 = (n25074 & n32878) | (n25074 & n36253) | (n32878 & n36253);
  assign n36256 = (n32213 & n36254) | (n32213 & n36255) | (n36254 & n36255);
  assign n25735 = n25448 & n36256;
  assign n25736 = ~n36251 & n25735;
  assign n32865 = n25459 & n25466;
  assign n32880 = n25736 | n32865;
  assign n36289 = n25785 | n32880;
  assign n32881 = n25459 | n25736;
  assign n36290 = n25785 | n32881;
  assign n36291 = (n32672 & n36289) | (n32672 & n36290) | (n36289 & n36290);
  assign n36292 = n25785 & n32880;
  assign n36293 = n25785 & n32881;
  assign n36294 = (n32672 & n36292) | (n32672 & n36293) | (n36292 & n36293);
  assign n25788 = n36291 & ~n36294;
  assign n25789 = x138 & x156;
  assign n25790 = ~n25788 & n25789;
  assign n25791 = n25788 & ~n25789;
  assign n25792 = n25790 | n25791;
  assign n32866 = (n25459 & n32672) | (n25459 & n32865) | (n32672 & n32865);
  assign n36243 = n25460 & n25466;
  assign n36244 = (n25459 & n25460) | (n25459 & n36243) | (n25460 & n36243);
  assign n32870 = (n25460 & n32672) | (n25460 & n36244) | (n32672 & n36244);
  assign n25731 = ~n32866 & n32870;
  assign n32872 = n25722 | n25731;
  assign n36295 = n25792 | n32872;
  assign n36245 = n25401 | n25731;
  assign n36246 = (n25722 & n25731) | (n25722 & n36245) | (n25731 & n36245);
  assign n36296 = n25792 | n36246;
  assign n36297 = (n32502 & n36295) | (n32502 & n36296) | (n36295 & n36296);
  assign n36298 = n25792 & n32872;
  assign n36299 = n25792 & n36246;
  assign n36300 = (n32502 & n36298) | (n32502 & n36299) | (n36298 & n36299);
  assign n25795 = n36297 & ~n36300;
  assign n25796 = n25727 & n25795;
  assign n36301 = n25471 | n25484;
  assign n36302 = (n25484 & n25724) | (n25484 & n36301) | (n25724 & n36301);
  assign n32926 = n25796 & n36302;
  assign n32927 = (n25796 & n32667) | (n25796 & n32926) | (n32667 & n32926);
  assign n25725 = n25471 & n25724;
  assign n25798 = n25725 | n25795;
  assign n32850 = n25477 & n25484;
  assign n32928 = n25798 | n32850;
  assign n36303 = n25477 | n25795;
  assign n36304 = n25725 | n36303;
  assign n32930 = (n32667 & n32928) | (n32667 & n36304) | (n32928 & n36304);
  assign n25800 = ~n32927 & n32930;
  assign n25801 = x137 & x157;
  assign n25802 = n25800 & n25801;
  assign n25803 = n25800 | n25801;
  assign n25804 = ~n25802 & n25803;
  assign n32851 = (n25477 & n32667) | (n25477 & n32850) | (n32667 & n32850);
  assign n36305 = n25478 & n25484;
  assign n36306 = (n25477 & n25478) | (n25477 & n36305) | (n25478 & n36305);
  assign n32855 = (n25478 & n32667) | (n25478 & n36306) | (n32667 & n36306);
  assign n25717 = ~n32851 & n32855;
  assign n32856 = n25493 | n25717;
  assign n32931 = n25804 & n32856;
  assign n32932 = n25717 & n25804;
  assign n32933 = (n32766 & n32931) | (n32766 & n32932) | (n32931 & n32932);
  assign n32934 = n25804 | n32856;
  assign n32935 = n25717 | n25804;
  assign n32936 = (n32766 & n32934) | (n32766 & n32935) | (n32934 & n32935);
  assign n25807 = ~n32933 & n32936;
  assign n25808 = x136 & x158;
  assign n25809 = x135 & x159;
  assign n25810 = n25808 | n25809;
  assign n25811 = n25808 & n25809;
  assign n25812 = n25810 & ~n25811;
  assign n25813 = n25807 | n25812;
  assign n25814 = n25807 & n25812;
  assign n25815 = n25813 & ~n25814;
  assign n32937 = n36238 | n25815;
  assign n32938 = n32847 | n32937;
  assign n32939 = n36238 & n25815;
  assign n32940 = (n25815 & n32847) | (n25815 & n32939) | (n32847 & n32939);
  assign n25818 = n32938 & ~n32940;
  assign n25819 = x134 & x160;
  assign n25820 = ~n25818 & n25819;
  assign n25821 = n25818 & ~n25819;
  assign n25822 = n25820 | n25821;
  assign n25823 = n25712 | n25822;
  assign n25824 = n25712 & n25822;
  assign n25825 = n25823 & ~n25824;
  assign n25826 = n32845 | n25825;
  assign n25827 = n32845 & n25825;
  assign n25828 = n25826 & ~n25827;
  assign n25829 = n25696 & n25828;
  assign n25830 = n25696 | n25828;
  assign n25831 = ~n25829 & n25830;
  assign n25832 = n25695 & ~n25831;
  assign n25833 = ~n25695 & n25831;
  assign n25834 = n25832 | n25833;
  assign n25835 = n32836 | n25834;
  assign n25836 = n32836 & n25834;
  assign n25837 = n25835 & ~n25836;
  assign n25838 = n25693 & n25837;
  assign n25839 = n25693 | n25837;
  assign n25840 = ~n25838 & n25839;
  assign n25841 = n32834 | n25840;
  assign n25842 = n32834 & n25840;
  assign n25843 = n25841 & ~n25842;
  assign n25844 = n32831 & n25843;
  assign n25845 = n32831 | n25843;
  assign n25846 = ~n25844 & n25845;
  assign n25847 = x130 & x164;
  assign n25848 = x129 & x165;
  assign n25849 = n25847 & n25848;
  assign n25850 = n25847 | n25848;
  assign n25851 = ~n25849 & n25850;
  assign n25852 = n25846 & n25851;
  assign n25853 = n25846 | n25851;
  assign n25854 = ~n25852 & n25853;
  assign n25855 = n32829 | n25854;
  assign n25856 = n32829 & n25854;
  assign n25857 = n25855 & ~n25856;
  assign n25663 = n32643 & n25539;
  assign n32822 = n25539 & n25540;
  assign n32823 = (n25540 & n32643) | (n25540 & n32822) | (n32643 & n32822);
  assign n25666 = ~n25663 & n32823;
  assign n36228 = n25550 | n25666;
  assign n36229 = (n25546 & n25666) | (n25546 & n36228) | (n25666 & n36228);
  assign n36307 = n25857 & n36229;
  assign n36308 = n25666 & n25857;
  assign n36309 = (n32784 & n36307) | (n32784 & n36308) | (n36307 & n36308);
  assign n36310 = n25857 | n36229;
  assign n36311 = n25666 | n25857;
  assign n36312 = (n32784 & n36310) | (n32784 & n36311) | (n36310 & n36311);
  assign n25860 = ~n36309 & n36312;
  assign n25861 = x128 & x166;
  assign n25862 = n25860 & n25861;
  assign n25863 = n25860 | n25861;
  assign n25864 = ~n25862 & n25863;
  assign n25865 = x127 & x167;
  assign n25866 = n25864 & n25865;
  assign n25867 = n25864 | n25865;
  assign n25868 = ~n25866 & n25867;
  assign n25869 = n25662 & ~n25868;
  assign n25870 = ~n25662 & n25868;
  assign n25871 = n25869 | n25870;
  assign n25872 = n32819 | n25871;
  assign n25873 = n32819 & n25871;
  assign n25874 = n25872 & ~n25873;
  assign n25875 = x125 & x169;
  assign n25876 = n25874 | n25875;
  assign n25877 = n25874 & n25875;
  assign n25878 = n25876 & ~n25877;
  assign n25880 = n25346 | n25654;
  assign n32941 = n25561 & ~n25654;
  assign n32942 = (~n25346 & n25561) | (~n25346 & n32941) | (n25561 & n32941);
  assign n25882 = n25880 & n32942;
  assign n32943 = n25570 | n25882;
  assign n32944 = (n25579 & n25882) | (n25579 & n32943) | (n25882 & n32943);
  assign n25884 = ~n25878 & n32944;
  assign n25885 = n25878 & ~n32944;
  assign n25886 = n25884 | n25885;
  assign n25887 = x124 & x170;
  assign n25888 = n25886 & n25887;
  assign n25889 = n25886 | n25887;
  assign n25890 = ~n25888 & n25889;
  assign n25892 = n25570 | n25579;
  assign n32945 = (n25571 & n25572) | (n25571 & ~n25579) | (n25572 & ~n25579);
  assign n25894 = n25892 & n32945;
  assign n32946 = n25582 | n25894;
  assign n32947 = (n25894 & n32787) | (n25894 & n32946) | (n32787 & n32946);
  assign n25896 = ~n25890 & n32947;
  assign n25897 = n25890 & ~n32947;
  assign n25898 = n25896 | n25897;
  assign n25899 = x123 & x171;
  assign n25900 = n25898 & ~n25899;
  assign n25901 = ~n25898 & n25899;
  assign n25902 = n25900 | n25901;
  assign n25904 = n25582 | n32787;
  assign n32948 = (n25583 & n25584) | (n25583 & ~n32787) | (n25584 & ~n32787);
  assign n25906 = n25904 & n32948;
  assign n32949 = n25594 | n25906;
  assign n32950 = (n25906 & n32793) | (n25906 & n32949) | (n32793 & n32949);
  assign n25908 = n25902 & n32950;
  assign n25909 = n25902 | n32950;
  assign n25910 = ~n25908 & n25909;
  assign n25911 = x122 & x172;
  assign n25912 = ~n25910 & n25911;
  assign n25913 = n25910 & ~n25911;
  assign n25914 = n25912 | n25913;
  assign n25915 = n25594 | n32793;
  assign n32951 = (n25595 & n25596) | (n25595 & ~n32793) | (n25596 & ~n32793);
  assign n25917 = n25915 & n32951;
  assign n25918 = n32814 | n25917;
  assign n25919 = n25914 & n25918;
  assign n25920 = n25914 | n25918;
  assign n25921 = ~n25919 & n25920;
  assign n32952 = ~n25650 & n25921;
  assign n32953 = ~n32811 & n32952;
  assign n32954 = n25650 & ~n25921;
  assign n32955 = (~n25921 & n32811) | (~n25921 & n32954) | (n32811 & n32954);
  assign n25924 = n32953 | n32955;
  assign n25925 = x121 & x173;
  assign n25926 = n25924 & n25925;
  assign n25927 = n25924 | n25925;
  assign n25928 = ~n25926 & n25927;
  assign n32956 = n25622 & n25928;
  assign n32957 = (n25928 & n32805) | (n25928 & n32956) | (n32805 & n32956);
  assign n32958 = n25622 | n25928;
  assign n32959 = n32805 | n32958;
  assign n25931 = ~n32957 & n32959;
  assign n25932 = n25644 & n25931;
  assign n25933 = n25644 | n25931;
  assign n25934 = ~n25932 & n25933;
  assign n25935 = n32809 & n25934;
  assign n25936 = n32809 | n25934;
  assign n25937 = ~n25935 & n25936;
  assign n25938 = n25642 & n25937;
  assign n25939 = n25642 | n25937;
  assign n25940 = ~n25938 & n25939;
  assign n32960 = n25634 & n25635;
  assign n32961 = (n25634 & n25638) | (n25634 & n32960) | (n25638 & n32960);
  assign n25943 = n25940 & ~n32961;
  assign n25944 = ~n25940 & n32961;
  assign n25945 = n25943 | n25944;
  assign n32962 = n25932 | n25934;
  assign n32963 = (n25932 & n32809) | (n25932 & n32962) | (n32809 & n32962);
  assign n25947 = x121 & x174;
  assign n25948 = n25926 | n32957;
  assign n32964 = n25910 & n25917;
  assign n32965 = (n25910 & n32814) | (n25910 & n32964) | (n32814 & n32964);
  assign n25950 = n25898 | n32950;
  assign n32966 = (n25899 & n25901) | (n25899 & ~n32950) | (n25901 & ~n32950);
  assign n25953 = n25950 & n32966;
  assign n25954 = n32965 | n25953;
  assign n25955 = n25886 | n32947;
  assign n32967 = ~n25886 & n25887;
  assign n32968 = (n25887 & ~n32947) | (n25887 & n32967) | (~n32947 & n32967);
  assign n25958 = n25955 & n32968;
  assign n32969 = n25898 | n25958;
  assign n32970 = (n25958 & n32950) | (n25958 & n32969) | (n32950 & n32969);
  assign n25960 = x125 & x170;
  assign n25961 = n25874 & n32944;
  assign n32971 = (n25875 & n25877) | (n25875 & n32944) | (n25877 & n32944);
  assign n25964 = ~n25961 & n32971;
  assign n32972 = n25886 | n25964;
  assign n32973 = (n25964 & n32947) | (n25964 & n32972) | (n32947 & n32972);
  assign n25966 = n32821 | n25868;
  assign n25967 = n32821 & n25868;
  assign n25968 = n25966 & ~n25967;
  assign n25969 = n32819 & n25968;
  assign n32974 = n25659 & n25968;
  assign n32975 = (n25659 & n32819) | (n25659 & n32974) | (n32819 & n32974);
  assign n25972 = ~n25969 & n32975;
  assign n32976 = n25874 | n25972;
  assign n32977 = (n25972 & n32944) | (n25972 & n32976) | (n32944 & n32976);
  assign n25974 = n32821 | n25864;
  assign n25977 = n25348 | n25553;
  assign n32825 = (n25666 & n32784) | (n25666 & n36229) | (n32784 & n36229);
  assign n25978 = ~n25857 & n25861;
  assign n25979 = n25857 & ~n25861;
  assign n25980 = n25978 | n25979;
  assign n25981 = ~n32825 & n25980;
  assign n25982 = n32825 & ~n25980;
  assign n25983 = n25981 | n25982;
  assign n25984 = n25977 & n25983;
  assign n25975 = n25256 | n25657;
  assign n32978 = n25975 & n25984;
  assign n32979 = (n25260 & n25984) | (n25260 & n32978) | (n25984 & n32978);
  assign n32980 = n25865 & ~n32979;
  assign n32981 = n25974 & n32980;
  assign n25988 = n32819 | n32981;
  assign n25990 = ~n25843 & n25847;
  assign n25991 = n25843 & ~n25847;
  assign n25992 = n25990 | n25991;
  assign n25993 = ~n32831 & n25992;
  assign n25994 = n32831 & ~n25992;
  assign n25995 = n25993 | n25994;
  assign n25996 = n25681 | n25995;
  assign n25997 = n25663 | n25996;
  assign n25998 = n25356 | n25681;
  assign n25999 = n25247 | n25998;
  assign n25679 = n25671 & n25678;
  assign n26000 = n25669 & ~n25679;
  assign n26001 = n25533 | n26000;
  assign n26002 = n25995 & n26001;
  assign n26003 = n25999 & n26002;
  assign n26004 = n25997 & ~n26003;
  assign n26005 = n25848 & n26004;
  assign n26006 = n25846 & n25847;
  assign n32982 = n26002 | n26006;
  assign n32983 = (n25999 & n26006) | (n25999 & n32982) | (n26006 & n32982);
  assign n26009 = n25807 & n25808;
  assign n26010 = n25807 | n25808;
  assign n26011 = ~n26009 & n26010;
  assign n32984 = n36238 | n26011;
  assign n32985 = n32847 | n32984;
  assign n26014 = n25801 & n25808;
  assign n26015 = n25801 | n25808;
  assign n26016 = ~n26014 & n26015;
  assign n26017 = n25800 & n26016;
  assign n26018 = n25800 | n26016;
  assign n26019 = ~n26017 & n26018;
  assign n32988 = n26019 | n32856;
  assign n32989 = n25717 | n26019;
  assign n32990 = (n32766 & n32988) | (n32766 & n32989) | (n32988 & n32989);
  assign n25495 = n36217 & ~n25494;
  assign n32991 = n26019 & n32856;
  assign n32992 = n25717 & n26019;
  assign n32993 = (n32766 & n32991) | (n32766 & n32992) | (n32991 & n32992);
  assign n32994 = n25496 & ~n32993;
  assign n32995 = (n25495 & ~n32993) | (n25495 & n32994) | (~n32993 & n32994);
  assign n26023 = n32990 & n32995;
  assign n32986 = n25380 | n36238;
  assign n32996 = n26023 & n32986;
  assign n32997 = (n26023 & n32585) | (n26023 & n32996) | (n32585 & n32996);
  assign n33002 = ~n25809 & n32997;
  assign n33003 = (n25809 & n32985) | (n25809 & ~n33002) | (n32985 & ~n33002);
  assign n33004 = n25802 | n32856;
  assign n33005 = n25717 | n25802;
  assign n33006 = (n32766 & n33004) | (n32766 & n33005) | (n33004 & n33005);
  assign n32873 = (n32502 & n36246) | (n32502 & n32872) | (n36246 & n32872);
  assign n33007 = n25781 & n32881;
  assign n36313 = n25736 & n25781;
  assign n36314 = (n25781 & n32865) | (n25781 & n36313) | (n32865 & n36313);
  assign n33009 = (n32672 & n33007) | (n32672 & n36314) | (n33007 & n36314);
  assign n33015 = n25744 & n25774;
  assign n33016 = (n25774 & n36251) | (n25774 & n33015) | (n36251 & n33015);
  assign n36315 = n25744 & n25775;
  assign n36316 = (n25774 & n25775) | (n25774 & n36315) | (n25775 & n36315);
  assign n33020 = (n25775 & n36251) | (n25775 & n36316) | (n36251 & n36316);
  assign n26039 = ~n33016 & n33020;
  assign n26051 = x142 & x153;
  assign n26053 = x143 & x152;
  assign n33030 = n25754 & n25761;
  assign n36317 = n26053 & n36283;
  assign n36318 = (n26053 & n33030) | (n26053 & n36317) | (n33030 & n36317);
  assign n36319 = (n25761 & n26053) | (n25761 & n36317) | (n26053 & n36317);
  assign n33044 = (n36265 & n36318) | (n36265 & n36319) | (n36318 & n36319);
  assign n36320 = n26053 | n36283;
  assign n36321 = n33030 | n36320;
  assign n36322 = n25761 | n36320;
  assign n33047 = (n36265 & n36321) | (n36265 & n36322) | (n36321 & n36322);
  assign n26056 = ~n33044 & n33047;
  assign n26057 = n26051 & n26056;
  assign n26058 = n26051 | n26056;
  assign n26059 = ~n26057 & n26058;
  assign n33031 = (n25761 & n36265) | (n25761 & n33030) | (n36265 & n33030);
  assign n33032 = n25754 | n25761;
  assign n33034 = n25756 & n33032;
  assign n33035 = (n25756 & n36265) | (n25756 & n33034) | (n36265 & n33034);
  assign n26049 = ~n33031 & n33035;
  assign n33021 = n25749 & n25767;
  assign n33036 = n26049 | n33021;
  assign n33048 = n26059 | n33036;
  assign n33037 = n25767 | n26049;
  assign n33049 = n26059 | n33037;
  assign n33050 = (n32889 & n33048) | (n32889 & n33049) | (n33048 & n33049);
  assign n33051 = n26059 & n33036;
  assign n33052 = n26059 & n33037;
  assign n33053 = (n32889 & n33051) | (n32889 & n33052) | (n33051 & n33052);
  assign n26062 = n33050 & ~n33053;
  assign n26063 = x141 & x154;
  assign n26064 = n26062 | n26063;
  assign n26065 = n26062 & n26063;
  assign n26066 = n26064 & ~n26065;
  assign n36323 = (n25767 & n32888) | (n25767 & n33021) | (n32888 & n33021);
  assign n36324 = (n25741 & n25767) | (n25741 & n33021) | (n25767 & n33021);
  assign n36325 = (n36080 & n36323) | (n36080 & n36324) | (n36323 & n36324);
  assign n33023 = n25749 | n25767;
  assign n33025 = n25768 & n33023;
  assign n36326 = (n25768 & n32888) | (n25768 & n33025) | (n32888 & n33025);
  assign n36327 = (n25741 & n25768) | (n25741 & n33025) | (n25768 & n33025);
  assign n36328 = (n36080 & n36326) | (n36080 & n36327) | (n36326 & n36327);
  assign n26044 = ~n36325 & n36328;
  assign n36329 = n25744 | n26044;
  assign n36330 = (n25774 & n26044) | (n25774 & n36329) | (n26044 & n36329);
  assign n33054 = n26066 | n36330;
  assign n33028 = n25774 | n26044;
  assign n33055 = n26066 | n33028;
  assign n33056 = (n36251 & n33054) | (n36251 & n33055) | (n33054 & n33055);
  assign n33057 = n26066 & n36330;
  assign n33058 = n26066 & n33028;
  assign n33059 = (n36251 & n33057) | (n36251 & n33058) | (n33057 & n33058);
  assign n26069 = n33056 & ~n33059;
  assign n26070 = x140 & x155;
  assign n26071 = n26069 | n26070;
  assign n26072 = n26069 & n26070;
  assign n26073 = n26071 & ~n26072;
  assign n33060 = n26039 | n26073;
  assign n33061 = n33009 | n33060;
  assign n33062 = n26039 & n26073;
  assign n33063 = (n26073 & n33009) | (n26073 & n33062) | (n33009 & n33062);
  assign n26076 = n33061 & ~n33063;
  assign n26077 = x139 & x156;
  assign n26078 = n26076 | n26077;
  assign n26079 = n26076 & n26077;
  assign n26080 = n26078 & ~n26079;
  assign n36331 = n25736 | n25781;
  assign n36332 = n32865 | n36331;
  assign n36333 = n25782 & n36332;
  assign n37538 = (n25782 & n25784) | (n25782 & n32881) | (n25784 & n32881);
  assign n36335 = (n32672 & n36333) | (n32672 & n37538) | (n36333 & n37538);
  assign n26034 = ~n33009 & n36335;
  assign n33013 = n25788 | n26034;
  assign n33064 = n26080 | n33013;
  assign n33065 = n26034 | n26080;
  assign n33066 = (n32873 & n33064) | (n32873 & n33065) | (n33064 & n33065);
  assign n33067 = n26080 & n33013;
  assign n33068 = n26034 & n26080;
  assign n33069 = (n32873 & n33067) | (n32873 & n33068) | (n33067 & n33068);
  assign n26083 = n33066 & ~n33069;
  assign n26084 = x138 & x157;
  assign n26085 = ~n26083 & n26084;
  assign n26086 = n26083 & ~n26084;
  assign n26087 = n26085 | n26086;
  assign n37539 = n25731 | n25788;
  assign n37540 = n25722 | n37539;
  assign n36337 = n25788 | n36246;
  assign n36338 = (n32502 & n37540) | (n32502 & n36337) | (n37540 & n36337);
  assign n36339 = (n25789 & n25790) | (n25789 & ~n32872) | (n25790 & ~n32872);
  assign n36340 = (n25789 & n25790) | (n25789 & ~n36246) | (n25790 & ~n36246);
  assign n36341 = (~n32502 & n36339) | (~n32502 & n36340) | (n36339 & n36340);
  assign n26090 = n36338 & n36341;
  assign n33071 = n26087 & n26090;
  assign n33072 = (n26087 & n32927) | (n26087 & n33071) | (n32927 & n33071);
  assign n33073 = n26087 | n26090;
  assign n33074 = n32927 | n33073;
  assign n26094 = ~n33072 & n33074;
  assign n26095 = n25803 & n26094;
  assign n26096 = n33006 & n26095;
  assign n26097 = n25802 | n26094;
  assign n26098 = n32933 | n26097;
  assign n26099 = ~n26096 & n26098;
  assign n26100 = x137 & x158;
  assign n26101 = x136 & x159;
  assign n26102 = n26100 | n26101;
  assign n26103 = n26100 & n26101;
  assign n26104 = n26102 & ~n26103;
  assign n26105 = n26099 | n26104;
  assign n26106 = n26099 & n26104;
  assign n26107 = n26105 & ~n26106;
  assign n33075 = n26009 | n26107;
  assign n33076 = n32997 | n33075;
  assign n33077 = n26009 & n26107;
  assign n33078 = (n26107 & n32997) | (n26107 & n33077) | (n32997 & n33077);
  assign n26111 = n33076 & ~n33078;
  assign n26112 = n33003 & n26111;
  assign n32998 = n25809 & ~n32997;
  assign n32999 = n32985 & n32998;
  assign n33000 = n25711 | n32999;
  assign n33079 = n26112 & n33000;
  assign n33080 = (n26112 & n32838) | (n26112 & n33079) | (n32838 & n33079);
  assign n26115 = n32999 | n26111;
  assign n33081 = n25711 & n25818;
  assign n33083 = n26115 | n33081;
  assign n33084 = n25818 | n26115;
  assign n33085 = (n32838 & n33083) | (n32838 & n33084) | (n33083 & n33084);
  assign n26117 = ~n33080 & n33085;
  assign n26118 = x135 & x160;
  assign n26119 = n26117 & n26118;
  assign n26120 = n26117 | n26118;
  assign n26121 = ~n26119 & n26120;
  assign n26122 = x134 & x161;
  assign n26123 = n26121 & n26122;
  assign n26124 = n26121 | n26122;
  assign n26125 = ~n26123 & n26124;
  assign n33086 = n25711 | n25818;
  assign n33087 = n32838 | n33086;
  assign n36342 = ~n25711 & n25819;
  assign n36343 = (~n25818 & n25819) | (~n25818 & n36342) | (n25819 & n36342);
  assign n33089 = (n25820 & ~n32838) | (n25820 & n36343) | (~n32838 & n36343);
  assign n26128 = n33087 & n33089;
  assign n33090 = n25374 | n32842;
  assign n33091 = n32593 | n33090;
  assign n33092 = ~n25507 & n32838;
  assign n33093 = (n25507 & n36236) | (n25507 & ~n33092) | (n36236 & ~n33092);
  assign n36344 = n26128 | n33093;
  assign n36345 = (n25825 & n26128) | (n25825 & n36344) | (n26128 & n36344);
  assign n33095 = (n26128 & n33091) | (n26128 & n36345) | (n33091 & n36345);
  assign n26134 = ~n26125 & n33095;
  assign n26135 = n26125 & ~n33095;
  assign n26136 = n26134 | n26135;
  assign n26131 = n25825 & n33093;
  assign n26132 = n33091 & n26131;
  assign n26137 = n25826 & ~n26132;
  assign n26138 = n25696 & n26137;
  assign n26139 = n26136 | n26138;
  assign n33096 = n25831 | n26139;
  assign n33097 = (n26139 & n32836) | (n26139 & n33096) | (n32836 & n33096);
  assign n26141 = n25517 | n26138;
  assign n33098 = n25688 | n26141;
  assign n33099 = (n25687 & n26141) | (n25687 & n33098) | (n26141 & n33098);
  assign n26143 = n25696 | n26137;
  assign n26144 = n26136 & n26143;
  assign n26145 = n33099 & n26144;
  assign n26146 = n33097 & ~n26145;
  assign n26147 = x133 & x162;
  assign n26148 = n26146 & n26147;
  assign n26149 = n26146 | n26147;
  assign n26150 = ~n26148 & n26149;
  assign n26151 = x132 & x163;
  assign n26152 = n26150 & n26151;
  assign n26153 = n26150 | n26151;
  assign n26154 = ~n26152 & n26153;
  assign n36346 = n25831 | n36233;
  assign n36347 = n25517 | n25831;
  assign n36348 = (n25687 & n36346) | (n25687 & n36347) | (n36346 & n36347);
  assign n33100 = (n25695 & n25832) | (n25695 & ~n32836) | (n25832 & ~n32836);
  assign n26157 = n36348 & n33100;
  assign n33101 = n25362 | n25365;
  assign n33102 = (n25362 & n25690) | (n25362 & n33101) | (n25690 & n33101);
  assign n26159 = n25230 | n33102;
  assign n26160 = n25365 | n25690;
  assign n26161 = n25837 & n26160;
  assign n33103 = n26157 | n26161;
  assign n33104 = (n26157 & n26159) | (n26157 & n33103) | (n26159 & n33103);
  assign n26164 = ~n26154 & n33104;
  assign n26165 = n26154 & ~n33104;
  assign n26166 = n26164 | n26165;
  assign n26162 = n26159 & n26161;
  assign n26167 = n25691 | n25837;
  assign n26168 = n32780 | n26167;
  assign n26169 = ~n26162 & n26168;
  assign n26170 = n25693 & n26169;
  assign n26171 = n26166 | n26170;
  assign n26172 = n25844 | n26171;
  assign n26173 = n25530 | n26170;
  assign n26174 = n25679 | n26173;
  assign n26175 = n25693 | n26169;
  assign n26176 = n26166 & n26175;
  assign n26177 = n26174 & n26176;
  assign n26178 = n26172 & ~n26177;
  assign n26179 = x131 & x164;
  assign n26180 = x130 & x165;
  assign n26181 = n26179 & n26180;
  assign n26182 = n26179 | n26180;
  assign n26183 = ~n26181 & n26182;
  assign n26184 = n26178 & n26183;
  assign n26185 = n26178 | n26183;
  assign n26186 = ~n26184 & n26185;
  assign n26187 = ~n32983 & n26186;
  assign n26188 = n32983 & ~n26186;
  assign n26189 = n26187 | n26188;
  assign n26190 = n26005 | n26189;
  assign n33105 = n25857 | n26190;
  assign n33106 = (n26190 & n32825) | (n26190 & n33105) | (n32825 & n33105);
  assign n33107 = n25666 | n25848;
  assign n33108 = (n25666 & n26004) | (n25666 & n33107) | (n26004 & n33107);
  assign n33109 = n25551 | n33108;
  assign n33110 = (n32784 & n33108) | (n32784 & n33109) | (n33108 & n33109);
  assign n26194 = n25848 | n26004;
  assign n26195 = n26189 & n26194;
  assign n26196 = n33110 & n26195;
  assign n26197 = n33106 & ~n26196;
  assign n26198 = x129 & x166;
  assign n26199 = n26197 | n26198;
  assign n26200 = n26197 & n26198;
  assign n26201 = n26199 & ~n26200;
  assign n33111 = n25862 | n26201;
  assign n33112 = n32979 | n33111;
  assign n33113 = n25862 & n26201;
  assign n33114 = (n26201 & n32979) | (n26201 & n33113) | (n32979 & n33113);
  assign n26204 = n33112 & ~n33114;
  assign n26205 = x128 & x167;
  assign n26206 = n26204 & n26205;
  assign n26207 = n26204 | n26205;
  assign n26208 = ~n26206 & n26207;
  assign n33115 = ~n25865 & n32979;
  assign n33116 = (n25865 & n25974) | (n25865 & ~n33115) | (n25974 & ~n33115);
  assign n26210 = n26208 & n33116;
  assign n26211 = n25988 & n26210;
  assign n26212 = n32981 | n26208;
  assign n26213 = n25969 | n26212;
  assign n26214 = ~n26211 & n26213;
  assign n26215 = x127 & x168;
  assign n26216 = n26214 & n26215;
  assign n26217 = n26214 | n26215;
  assign n26218 = ~n26216 & n26217;
  assign n26219 = n32977 | n26218;
  assign n26220 = n32977 & n26218;
  assign n26221 = n26219 & ~n26220;
  assign n26222 = x126 & x169;
  assign n26223 = n26221 & n26222;
  assign n26224 = n26221 | n26222;
  assign n26225 = ~n26223 & n26224;
  assign n26226 = n32973 & n26225;
  assign n26227 = n32973 | n26225;
  assign n26228 = ~n26226 & n26227;
  assign n26229 = n25960 | n26228;
  assign n26230 = n25960 & n26228;
  assign n26231 = n26229 & ~n26230;
  assign n26232 = n32970 | n26231;
  assign n26233 = n32970 & n26231;
  assign n26234 = n26232 & ~n26233;
  assign n26235 = x124 & x171;
  assign n26236 = n26234 | n26235;
  assign n26237 = n26234 & n26235;
  assign n26238 = n26236 & ~n26237;
  assign n26239 = n25954 | n26238;
  assign n26240 = n25954 & n26238;
  assign n26241 = n26239 & ~n26240;
  assign n26242 = x123 & x172;
  assign n26243 = n26241 | n26242;
  assign n26244 = n26241 & n26242;
  assign n26245 = n26243 & ~n26244;
  assign n33117 = n25650 & n25921;
  assign n33118 = (n25921 & n32811) | (n25921 & n33117) | (n32811 & n33117);
  assign n33119 = n25910 | n25917;
  assign n33120 = n32814 | n33119;
  assign n26248 = n25911 & ~n32965;
  assign n26249 = n33120 & n26248;
  assign n26250 = n33118 | n26249;
  assign n26251 = n26245 & n26250;
  assign n26252 = n26245 | n26250;
  assign n26253 = ~n26251 & n26252;
  assign n26254 = x122 & x173;
  assign n26255 = n26253 & n26254;
  assign n26256 = n26253 | n26254;
  assign n26257 = ~n26255 & n26256;
  assign n26258 = n25948 & n26257;
  assign n26259 = n25948 | n26257;
  assign n26260 = ~n26258 & n26259;
  assign n26261 = n25947 & n26260;
  assign n26262 = n25947 | n26260;
  assign n26263 = ~n26261 & n26262;
  assign n26264 = n32963 & n26263;
  assign n26265 = n32963 | n26263;
  assign n26266 = ~n26264 & n26265;
  assign n26267 = x120 & x175;
  assign n26268 = n26266 & n26267;
  assign n26269 = n26266 | n26267;
  assign n26270 = ~n26268 & n26269;
  assign n33121 = n25938 & n25939;
  assign n33122 = (n25939 & n32961) | (n25939 & n33121) | (n32961 & n33121);
  assign n26273 = n26270 & ~n33122;
  assign n26274 = ~n26270 & n33122;
  assign n26275 = n26273 | n26274;
  assign n33123 = n26268 & n26269;
  assign n33124 = (n26269 & n33122) | (n26269 & n33123) | (n33122 & n33123);
  assign n26278 = x121 & x175;
  assign n33125 = n26255 | n26257;
  assign n33126 = (n25948 & n26255) | (n25948 & n33125) | (n26255 & n33125);
  assign n26280 = n26237 | n26240;
  assign n33127 = n26230 | n32970;
  assign n33128 = (n26230 & n26231) | (n26230 & n33127) | (n26231 & n33127);
  assign n33129 = n26223 | n32973;
  assign n33130 = (n26223 & n26225) | (n26223 & n33129) | (n26225 & n33129);
  assign n33131 = n26216 | n32977;
  assign n33132 = (n26216 & n26218) | (n26216 & n33131) | (n26218 & n33131);
  assign n36349 = n26206 | n33116;
  assign n36350 = (n26206 & n26208) | (n26206 & n36349) | (n26208 & n36349);
  assign n33134 = (n25988 & n26206) | (n25988 & n36350) | (n26206 & n36350);
  assign n26285 = n26200 | n33114;
  assign n26286 = n26178 | n26179;
  assign n26287 = n26178 & n26179;
  assign n26288 = n26286 & ~n26287;
  assign n26289 = n32983 & n26288;
  assign n26290 = n32983 | n26288;
  assign n26291 = n26180 & n26290;
  assign n26292 = ~n26289 & n26291;
  assign n33135 = n26195 | n26292;
  assign n33136 = (n26292 & n33110) | (n26292 & n33135) | (n33110 & n33135);
  assign n33140 = n26148 | n26150;
  assign n33141 = (n26148 & n33104) | (n26148 & n33140) | (n33104 & n33140);
  assign n33145 = n26119 | n26121;
  assign n33146 = (n26119 & n33095) | (n26119 & n33145) | (n33095 & n33145);
  assign n26306 = n26099 & n26100;
  assign n26307 = n26099 | n26100;
  assign n26308 = ~n26306 & n26307;
  assign n33147 = n26009 & n26308;
  assign n33148 = (n26308 & n32997) | (n26308 & n33147) | (n32997 & n33147);
  assign n33149 = n26009 | n26308;
  assign n33150 = n32997 | n33149;
  assign n26311 = n26101 & n33150;
  assign n26312 = ~n33148 & n26311;
  assign n26313 = n33080 | n26312;
  assign n33161 = n26062 & n36330;
  assign n33162 = n26062 & n33028;
  assign n33163 = (n36251 & n33161) | (n36251 & n33162) | (n33161 & n33162);
  assign n37541 = (n26063 & n26065) | (n26063 & n33028) | (n26065 & n33028);
  assign n37542 = (n26063 & n26065) | (n26063 & n36330) | (n26065 & n36330);
  assign n36361 = (n36251 & n37541) | (n36251 & n37542) | (n37541 & n37542);
  assign n26323 = ~n33163 & n36361;
  assign n33154 = n26039 & n26069;
  assign n33167 = n26323 | n33154;
  assign n33168 = n26069 | n26323;
  assign n36362 = (n33167 & n33168) | (n33167 & n36314) | (n33168 & n36314);
  assign n36363 = (n33007 & n33167) | (n33007 & n33168) | (n33167 & n33168);
  assign n36364 = (n32672 & n36362) | (n32672 & n36363) | (n36362 & n36363);
  assign n33171 = n26056 & n33037;
  assign n36365 = n26049 & n26056;
  assign n36366 = (n26056 & n33021) | (n26056 & n36365) | (n33021 & n36365);
  assign n36367 = (n32888 & n33171) | (n32888 & n36366) | (n33171 & n36366);
  assign n36368 = (n25741 & n33171) | (n25741 & n36366) | (n33171 & n36366);
  assign n36369 = (n36080 & n36367) | (n36080 & n36368) | (n36367 & n36368);
  assign n33174 = n26056 | n33037;
  assign n36370 = n26049 | n26056;
  assign n36371 = n33021 | n36370;
  assign n36372 = (n32888 & n33174) | (n32888 & n36371) | (n33174 & n36371);
  assign n36373 = (n25741 & n33174) | (n25741 & n36371) | (n33174 & n36371);
  assign n36374 = (n36080 & n36372) | (n36080 & n36373) | (n36372 & n36373);
  assign n26327 = n26051 & n36374;
  assign n26328 = ~n36369 & n26327;
  assign n26330 = x142 & x154;
  assign n26332 = x143 & x153;
  assign n37544 = n26053 & n26332;
  assign n37782 = n36283 & n37544;
  assign n37545 = (n33030 & n37782) | (n33030 & n37544) | (n37782 & n37544);
  assign n36376 = n26332 & n36319;
  assign n36377 = (n36265 & n37545) | (n36265 & n36376) | (n37545 & n36376);
  assign n33177 = (n26332 & n36369) | (n26332 & n36377) | (n36369 & n36377);
  assign n37547 = n26053 | n26332;
  assign n37783 = (n26332 & n36283) | (n26332 & n37547) | (n36283 & n37547);
  assign n37548 = (n33030 & n37783) | (n33030 & n37547) | (n37783 & n37547);
  assign n36379 = n26332 | n36319;
  assign n36380 = (n36265 & n37548) | (n36265 & n36379) | (n37548 & n36379);
  assign n33179 = n36369 | n36380;
  assign n26335 = ~n33177 & n33179;
  assign n26336 = n26330 & n26335;
  assign n26337 = n26330 | n26335;
  assign n26338 = ~n26336 & n26337;
  assign n33180 = n26328 | n26338;
  assign n33181 = n33163 | n33180;
  assign n33182 = n26328 & n26338;
  assign n33183 = (n26338 & n33163) | (n26338 & n33182) | (n33163 & n33182);
  assign n26341 = n33181 & ~n33183;
  assign n26342 = x141 & x155;
  assign n26343 = n26341 | n26342;
  assign n26344 = n26341 & n26342;
  assign n26345 = n26343 & ~n26344;
  assign n26346 = ~n36364 & n26345;
  assign n26347 = n36364 & ~n26345;
  assign n26348 = n26346 | n26347;
  assign n26349 = x140 & x156;
  assign n26350 = n26348 & n26349;
  assign n26351 = n26348 | n26349;
  assign n26352 = ~n26350 & n26351;
  assign n36353 = (n26069 & n33154) | (n26069 & n36314) | (n33154 & n36314);
  assign n36354 = (n26069 & n33007) | (n26069 & n33154) | (n33007 & n33154);
  assign n36355 = (n32672 & n36353) | (n32672 & n36354) | (n36353 & n36354);
  assign n33156 = n26039 | n26069;
  assign n36356 = n33156 | n36314;
  assign n36357 = n33007 | n33156;
  assign n36358 = (n32672 & n36356) | (n32672 & n36357) | (n36356 & n36357);
  assign n26317 = ~n36355 & n36358;
  assign n26318 = n26070 & n26317;
  assign n33152 = n26034 & n26076;
  assign n33159 = n26318 | n33152;
  assign n36381 = n26352 | n33159;
  assign n33151 = n26076 & n33013;
  assign n33158 = n26318 | n33151;
  assign n36382 = n26352 | n33158;
  assign n36383 = (n32873 & n36381) | (n32873 & n36382) | (n36381 & n36382);
  assign n36384 = n26352 & n33159;
  assign n36385 = n26352 & n33158;
  assign n36386 = (n32873 & n36384) | (n32873 & n36385) | (n36384 & n36385);
  assign n26355 = n36383 & ~n36386;
  assign n26356 = x139 & x157;
  assign n26357 = n26355 | n26356;
  assign n26358 = n26355 & n26356;
  assign n26359 = n26357 & ~n26358;
  assign n33186 = n26076 | n33013;
  assign n33187 = n26034 | n26076;
  assign n36387 = (n32872 & n33186) | (n32872 & n33187) | (n33186 & n33187);
  assign n36388 = (n33186 & n33187) | (n33186 & n36246) | (n33187 & n36246);
  assign n36389 = (n32502 & n36387) | (n32502 & n36388) | (n36387 & n36388);
  assign n33189 = n26077 & ~n33151;
  assign n36390 = ~n26034 & n26077;
  assign n36391 = (~n26076 & n26077) | (~n26076 & n36390) | (n26077 & n36390);
  assign n33191 = (~n32873 & n33189) | (~n32873 & n36391) | (n33189 & n36391);
  assign n26363 = n36389 & n33191;
  assign n33184 = n26083 & n26090;
  assign n33192 = n26363 | n33184;
  assign n36392 = n26359 | n33192;
  assign n33193 = n26083 | n26363;
  assign n36393 = n26359 | n33193;
  assign n36394 = (n32927 & n36392) | (n32927 & n36393) | (n36392 & n36393);
  assign n36395 = n26359 & n33192;
  assign n36396 = n26359 & n33193;
  assign n36397 = (n32927 & n36395) | (n32927 & n36396) | (n36395 & n36396);
  assign n26367 = n36394 & ~n36397;
  assign n26368 = x138 & x158;
  assign n26369 = n26367 | n26368;
  assign n26370 = n26367 & n26368;
  assign n26371 = n26369 & ~n26370;
  assign n33195 = n26083 | n26090;
  assign n33196 = n32927 | n33195;
  assign n36398 = n26084 & ~n26090;
  assign n36399 = (~n26083 & n26084) | (~n26083 & n36398) | (n26084 & n36398);
  assign n33198 = (n26085 & ~n32927) | (n26085 & n36399) | (~n32927 & n36399);
  assign n26374 = n33196 & n33198;
  assign n33199 = n26095 | n26374;
  assign n36400 = ~n26371 & n33199;
  assign n36401 = ~n26371 & n26374;
  assign n36402 = (n33006 & n36400) | (n33006 & n36401) | (n36400 & n36401);
  assign n36403 = n26371 & ~n33199;
  assign n36404 = n26371 & ~n26374;
  assign n36405 = (~n33006 & n36403) | (~n33006 & n36404) | (n36403 & n36404);
  assign n26378 = n36402 | n36405;
  assign n26379 = x137 & x159;
  assign n26380 = n26378 & n26379;
  assign n26381 = n26378 | n26379;
  assign n26382 = ~n26380 & n26381;
  assign n33201 = n26306 | n26382;
  assign n33202 = n33148 | n33201;
  assign n33203 = n26306 & n26382;
  assign n33204 = (n26382 & n33148) | (n26382 & n33203) | (n33148 & n33203);
  assign n26386 = n33202 & ~n33204;
  assign n26387 = x136 & x160;
  assign n26388 = n26386 & n26387;
  assign n26389 = n26386 | n26387;
  assign n26390 = ~n26388 & n26389;
  assign n26391 = ~n26313 & n26390;
  assign n26392 = n26313 & ~n26390;
  assign n26393 = n26391 | n26392;
  assign n26394 = x135 & x161;
  assign n26395 = n26393 & n26394;
  assign n26396 = n26393 | n26394;
  assign n26397 = ~n26395 & n26396;
  assign n26398 = ~n33146 & n26397;
  assign n26399 = n33146 & ~n26397;
  assign n26400 = n26398 | n26399;
  assign n36406 = n26121 & n36345;
  assign n36407 = n26121 & n26128;
  assign n36408 = (n33091 & n36406) | (n33091 & n36407) | (n36406 & n36407);
  assign n33142 = (n26122 & n26123) | (n26122 & n33095) | (n26123 & n33095);
  assign n26303 = ~n36408 & n33142;
  assign n33143 = n26144 | n26303;
  assign n33205 = n26400 & n33143;
  assign n33206 = n26303 & n26400;
  assign n33207 = (n33099 & n33205) | (n33099 & n33206) | (n33205 & n33206);
  assign n33208 = n26400 | n33143;
  assign n33209 = n26303 | n26400;
  assign n33210 = (n33099 & n33208) | (n33099 & n33209) | (n33208 & n33209);
  assign n26403 = ~n33207 & n33210;
  assign n26404 = x134 & x162;
  assign n26405 = n26403 & n26404;
  assign n26406 = n26403 | n26404;
  assign n26407 = ~n26405 & n26406;
  assign n26408 = x133 & x163;
  assign n26409 = n26407 & n26408;
  assign n26410 = n26407 | n26408;
  assign n26411 = ~n26409 & n26410;
  assign n26412 = n33141 | n26411;
  assign n26413 = n33141 & n26411;
  assign n26414 = n26412 & ~n26413;
  assign n26294 = n26150 & n33104;
  assign n33137 = (n26151 & n26152) | (n26151 & n33104) | (n26152 & n33104);
  assign n26297 = ~n26294 & n33137;
  assign n36351 = n26175 | n26297;
  assign n36352 = (n26166 & n26297) | (n26166 & n36351) | (n26297 & n36351);
  assign n36409 = n26414 & n36352;
  assign n36410 = n26297 & n26414;
  assign n36411 = (n26174 & n36409) | (n26174 & n36410) | (n36409 & n36410);
  assign n36412 = n26414 | n36352;
  assign n36413 = n26297 | n26414;
  assign n36414 = (n26174 & n36412) | (n26174 & n36413) | (n36412 & n36413);
  assign n26417 = ~n36411 & n36414;
  assign n26418 = x132 & x164;
  assign n26419 = n26417 & n26418;
  assign n26420 = n26417 | n26418;
  assign n26421 = ~n26419 & n26420;
  assign n26422 = x131 & x165;
  assign n26423 = n26421 & n26422;
  assign n26424 = n26421 | n26422;
  assign n26425 = ~n26423 & n26424;
  assign n26426 = n26287 | n26289;
  assign n26427 = n26425 | n26426;
  assign n26428 = n26425 & n26426;
  assign n26429 = n26427 & ~n26428;
  assign n26430 = n33136 & n26429;
  assign n26431 = n33136 | n26429;
  assign n26432 = ~n26430 & n26431;
  assign n26433 = x130 & x166;
  assign n26434 = n26432 & n26433;
  assign n26435 = n26432 | n26433;
  assign n26436 = ~n26434 & n26435;
  assign n26437 = x129 & x167;
  assign n26438 = n26436 & n26437;
  assign n26439 = n26436 | n26437;
  assign n26440 = ~n26438 & n26439;
  assign n26441 = n26285 | n26440;
  assign n26442 = n26285 & n26440;
  assign n26443 = n26441 & ~n26442;
  assign n26444 = x128 & x168;
  assign n26445 = n26443 | n26444;
  assign n26446 = n26443 & n26444;
  assign n26447 = n26445 & ~n26446;
  assign n26448 = n33134 | n26447;
  assign n26449 = n33134 & n26447;
  assign n26450 = n26448 & ~n26449;
  assign n26451 = x127 & x169;
  assign n26452 = n26450 | n26451;
  assign n26453 = n26450 & n26451;
  assign n26454 = n26452 & ~n26453;
  assign n26455 = n33132 | n26454;
  assign n26456 = n33132 & n26454;
  assign n26457 = n26455 & ~n26456;
  assign n26458 = x126 & x170;
  assign n26459 = n26457 | n26458;
  assign n26460 = n26457 & n26458;
  assign n26461 = n26459 & ~n26460;
  assign n26462 = n33130 | n26461;
  assign n26463 = n33130 & n26461;
  assign n26464 = n26462 & ~n26463;
  assign n26465 = x125 & x171;
  assign n26466 = n26464 | n26465;
  assign n26467 = n26464 & n26465;
  assign n26468 = n26466 & ~n26467;
  assign n26469 = n33128 | n26468;
  assign n26470 = n33128 & n26468;
  assign n26471 = n26469 & ~n26470;
  assign n26472 = x124 & x172;
  assign n26473 = n26471 | n26472;
  assign n26474 = n26471 & n26472;
  assign n26475 = n26473 & ~n26474;
  assign n26476 = n26280 | n26475;
  assign n26477 = n26280 & n26475;
  assign n26478 = n26476 & ~n26477;
  assign n26479 = x123 & x173;
  assign n26480 = n26478 | n26479;
  assign n26481 = n26478 & n26479;
  assign n26482 = n26480 & ~n26481;
  assign n33211 = n26243 & n26244;
  assign n33212 = (n26243 & n26250) | (n26243 & n33211) | (n26250 & n33211);
  assign n26485 = n26482 | n33212;
  assign n26486 = n26482 & n33212;
  assign n26487 = n26485 & ~n26486;
  assign n26488 = x122 & x174;
  assign n26489 = n26487 | n26488;
  assign n26490 = n26487 & n26488;
  assign n26491 = n26489 & ~n26490;
  assign n26492 = n33126 | n26491;
  assign n26493 = n33126 & n26491;
  assign n26494 = n26492 & ~n26493;
  assign n26495 = n26261 | n26494;
  assign n26496 = n26264 | n26495;
  assign n26497 = n32963 | n26261;
  assign n26498 = n26262 & n26494;
  assign n26499 = n26497 & n26498;
  assign n26500 = n26496 & ~n26499;
  assign n26501 = n26278 | n26500;
  assign n26502 = n26278 & n26500;
  assign n26503 = n26501 & ~n26502;
  assign n26504 = n33124 & n26503;
  assign n26505 = n33124 | n26503;
  assign n26506 = ~n26504 & n26505;
  assign n26507 = n26502 | n26504;
  assign n26508 = x122 & x175;
  assign n26509 = n33126 | n26487;
  assign n33213 = ~n26487 & n26488;
  assign n33214 = (n26488 & ~n33126) | (n26488 & n33213) | (~n33126 & n33213);
  assign n26512 = n26509 & n33214;
  assign n33215 = n26498 | n26512;
  assign n33216 = (n26497 & n26512) | (n26497 & n33215) | (n26512 & n33215);
  assign n26514 = x123 & x174;
  assign n26515 = n26478 | n33212;
  assign n33217 = ~n26478 & n26479;
  assign n33218 = (n26479 & ~n33212) | (n26479 & n33217) | (~n33212 & n33217);
  assign n26518 = n26515 & n33218;
  assign n33219 = n26487 | n26518;
  assign n33220 = (n26518 & n33126) | (n26518 & n33219) | (n33126 & n33219);
  assign n26520 = x124 & x173;
  assign n33221 = n26237 | n26471;
  assign n33222 = n26240 | n33221;
  assign n26522 = n25954 | n26237;
  assign n26523 = n26236 & n26471;
  assign n33223 = n26472 & ~n26523;
  assign n33224 = (n26472 & ~n26522) | (n26472 & n33223) | (~n26522 & n33223);
  assign n26526 = n33222 & n33224;
  assign n33225 = n26478 | n26526;
  assign n33226 = (n26526 & n33212) | (n26526 & n33225) | (n33212 & n33225);
  assign n26528 = x125 & x172;
  assign n26529 = n33128 | n26464;
  assign n26530 = n32970 | n26230;
  assign n26531 = n26229 & n26464;
  assign n26532 = n26530 & n26531;
  assign n26533 = n26465 & ~n26532;
  assign n26534 = n26529 & n26533;
  assign n33227 = n26523 | n26534;
  assign n33228 = (n26522 & n26534) | (n26522 & n33227) | (n26534 & n33227);
  assign n26536 = n33130 | n26457;
  assign n33229 = ~n26457 & n26458;
  assign n33230 = (n26458 & ~n33130) | (n26458 & n33229) | (~n33130 & n33229);
  assign n26539 = n26536 & n33230;
  assign n26541 = n33132 & n26450;
  assign n33231 = (n26451 & n26453) | (n26451 & n33132) | (n26453 & n33132);
  assign n26544 = ~n26541 & n33231;
  assign n33232 = n26457 | n26544;
  assign n33233 = (n26544 & n33130) | (n26544 & n33232) | (n33130 & n33232);
  assign n36415 = n26443 & n36350;
  assign n36416 = n26206 & n26443;
  assign n36417 = (n25988 & n36415) | (n25988 & n36416) | (n36415 & n36416);
  assign n36418 = (n26444 & n26446) | (n26444 & n36350) | (n26446 & n36350);
  assign n37784 = n26205 & n26444;
  assign n37785 = n26204 & n37784;
  assign n37550 = (n26443 & n26444) | (n26443 & n37785) | (n26444 & n37785);
  assign n36420 = (n25988 & n36418) | (n25988 & n37550) | (n36418 & n37550);
  assign n26549 = ~n36417 & n36420;
  assign n33235 = n26450 | n26549;
  assign n33236 = (n26549 & n33132) | (n26549 & n33235) | (n33132 & n33235);
  assign n33237 = n26200 | n26436;
  assign n33238 = n33114 | n33237;
  assign n33239 = n25862 | n26200;
  assign n33240 = n32979 | n33239;
  assign n26553 = n26429 | n26433;
  assign n26554 = n26429 & n26433;
  assign n26555 = n26553 & ~n26554;
  assign n26556 = n33136 | n26555;
  assign n26557 = n33136 & n26555;
  assign n26558 = n26199 & ~n26557;
  assign n26559 = n26556 & n26558;
  assign n26560 = n33240 & n26559;
  assign n26561 = n33238 & ~n26560;
  assign n26562 = n26437 & n26561;
  assign n33241 = n26443 | n26562;
  assign n36421 = (n26562 & n33241) | (n26562 & n36350) | (n33241 & n36350);
  assign n36422 = (n26206 & n26562) | (n26206 & n33241) | (n26562 & n33241);
  assign n36423 = (n25988 & n36421) | (n25988 & n36422) | (n36421 & n36422);
  assign n26564 = x129 & x168;
  assign n36424 = n26434 | n26559;
  assign n36425 = (n26434 & n33240) | (n26434 & n36424) | (n33240 & n36424);
  assign n26566 = x131 & x166;
  assign n26567 = n32983 | n26287;
  assign n33139 = (n26174 & n26297) | (n26174 & n36352) | (n26297 & n36352);
  assign n26568 = ~n26414 & n26418;
  assign n26569 = n26414 & ~n26418;
  assign n26570 = n26568 | n26569;
  assign n26571 = ~n33139 & n26570;
  assign n26572 = n33139 & ~n26570;
  assign n26573 = n26571 | n26572;
  assign n26574 = n26286 & n26573;
  assign n33243 = n26419 | n26574;
  assign n33244 = (n26419 & n26567) | (n26419 & n33243) | (n26567 & n33243);
  assign n26591 = x135 & x162;
  assign n26600 = x137 & x160;
  assign n33255 = n26312 & n26386;
  assign n33264 = n26306 | n26378;
  assign n33265 = n33148 | n33264;
  assign n26602 = n26307 & n26378;
  assign n33260 = n26009 | n26306;
  assign n33262 = n26602 & n33260;
  assign n33263 = (n26602 & n32997) | (n26602 & n33262) | (n32997 & n33262);
  assign n33266 = n26379 & ~n33263;
  assign n33267 = n33265 & n33266;
  assign n33268 = n33255 | n33267;
  assign n33269 = n26386 | n33267;
  assign n33270 = (n33080 & n33268) | (n33080 & n33269) | (n33268 & n33269);
  assign n33272 = n26367 | n26374;
  assign n36426 = n26095 | n33272;
  assign n33273 = (n33006 & n36426) | (n33006 & n33272) | (n36426 & n33272);
  assign n33275 = n26367 & n26374;
  assign n36427 = (n26095 & n26367) | (n26095 & n33275) | (n26367 & n33275);
  assign n36428 = n26368 & ~n36427;
  assign n36429 = n26368 & ~n33275;
  assign n36430 = (~n33006 & n36428) | (~n33006 & n36429) | (n36428 & n36429);
  assign n26611 = n33273 & n36430;
  assign n33276 = (n33006 & n36427) | (n33006 & n33275) | (n36427 & n33275);
  assign n36431 = n26355 & n26363;
  assign n36432 = (n26355 & n33184) | (n26355 & n36431) | (n33184 & n36431);
  assign n33313 = n26355 & n33193;
  assign n33314 = (n32927 & n36432) | (n32927 & n33313) | (n36432 & n33313);
  assign n26636 = n26070 | n26317;
  assign n26637 = n26348 & n26636;
  assign n33300 = n26034 | n26318;
  assign n33302 = n26637 & n33300;
  assign n33299 = n26318 | n33013;
  assign n33303 = n26637 & n33299;
  assign n33304 = (n32873 & n33302) | (n32873 & n33303) | (n33302 & n33303);
  assign n33278 = n26341 & n33167;
  assign n33280 = n26328 & n26335;
  assign n36433 = (n26335 & n33162) | (n26335 & n33280) | (n33162 & n33280);
  assign n36434 = (n26335 & n33161) | (n26335 & n33280) | (n33161 & n33280);
  assign n36435 = (n36251 & n36433) | (n36251 & n36434) | (n36433 & n36434);
  assign n33282 = n26328 | n26335;
  assign n33284 = n26330 & n33282;
  assign n36436 = (n26330 & n33162) | (n26330 & n33284) | (n33162 & n33284);
  assign n36437 = (n26330 & n33161) | (n26330 & n33284) | (n33161 & n33284);
  assign n36438 = (n36251 & n36436) | (n36251 & n36437) | (n36436 & n36437);
  assign n26617 = ~n36435 & n36438;
  assign n26619 = x142 & x155;
  assign n26621 = x143 & x154;
  assign n37552 = n26332 & n26621;
  assign n37885 = n36319 & n37552;
  assign n37887 = n26621 & n37544;
  assign n37920 = n36283 & n37887;
  assign n37888 = (n33030 & n37920) | (n33030 & n37887) | (n37920 & n37887);
  assign n37788 = (n36265 & n37885) | (n36265 & n37888) | (n37885 & n37888);
  assign n37553 = (n36369 & n37788) | (n36369 & n37552) | (n37788 & n37552);
  assign n36440 = (n26621 & n33280) | (n26621 & n37553) | (n33280 & n37553);
  assign n36441 = (n26335 & n26621) | (n26335 & n37553) | (n26621 & n37553);
  assign n36442 = (n33162 & n36440) | (n33162 & n36441) | (n36440 & n36441);
  assign n36443 = (n33161 & n36440) | (n33161 & n36441) | (n36440 & n36441);
  assign n36444 = (n36251 & n36442) | (n36251 & n36443) | (n36442 & n36443);
  assign n37555 = n26332 | n26621;
  assign n37889 = (n26621 & n36319) | (n26621 & n37555) | (n36319 & n37555);
  assign n37891 = n26621 | n37544;
  assign n37921 = (n26621 & n36283) | (n26621 & n37891) | (n36283 & n37891);
  assign n37892 = (n33030 & n37921) | (n33030 & n37891) | (n37921 & n37891);
  assign n37791 = (n36265 & n37889) | (n36265 & n37892) | (n37889 & n37892);
  assign n37556 = (n36369 & n37791) | (n36369 & n37555) | (n37791 & n37555);
  assign n36446 = n33280 | n37556;
  assign n36447 = n26335 | n37556;
  assign n36448 = (n33162 & n36446) | (n33162 & n36447) | (n36446 & n36447);
  assign n36449 = (n33161 & n36446) | (n33161 & n36447) | (n36446 & n36447);
  assign n36450 = (n36251 & n36448) | (n36251 & n36449) | (n36448 & n36449);
  assign n26624 = ~n36444 & n36450;
  assign n26625 = n26619 & n26624;
  assign n26626 = n26619 | n26624;
  assign n26627 = ~n26625 & n26626;
  assign n33295 = n26617 | n26627;
  assign n36451 = n33278 | n33295;
  assign n33277 = n26341 & n33168;
  assign n36452 = n33277 | n33295;
  assign n36453 = (n33009 & n36451) | (n33009 & n36452) | (n36451 & n36452);
  assign n33297 = n26617 & n26627;
  assign n36454 = (n26627 & n33278) | (n26627 & n33297) | (n33278 & n33297);
  assign n36455 = (n26627 & n33277) | (n26627 & n33297) | (n33277 & n33297);
  assign n36456 = (n33009 & n36454) | (n33009 & n36455) | (n36454 & n36455);
  assign n26630 = n36453 & ~n36456;
  assign n26631 = x141 & x156;
  assign n26632 = n26630 | n26631;
  assign n26633 = n26630 & n26631;
  assign n26634 = n26632 & ~n26633;
  assign n33305 = n26341 | n33168;
  assign n33306 = n26341 | n33167;
  assign n33307 = (n33009 & n33305) | (n33009 & n33306) | (n33305 & n33306);
  assign n37557 = ~n26341 & n26342;
  assign n37558 = (n26342 & ~n33167) | (n26342 & n37557) | (~n33167 & n37557);
  assign n36458 = n26342 & ~n33277;
  assign n36459 = (~n33009 & n37558) | (~n33009 & n36458) | (n37558 & n36458);
  assign n26641 = n33307 & n36459;
  assign n33308 = n26634 | n26641;
  assign n33309 = n33304 | n33308;
  assign n33310 = n26634 & n26641;
  assign n33311 = (n26634 & n33304) | (n26634 & n33310) | (n33304 & n33310);
  assign n26645 = n33309 & ~n33311;
  assign n26646 = x140 & x157;
  assign n26647 = n26645 | n26646;
  assign n26648 = n26645 & n26646;
  assign n26649 = n26647 & ~n26648;
  assign n37559 = n26318 | n26348;
  assign n37560 = n33152 | n37559;
  assign n37561 = n33151 | n37559;
  assign n36462 = (n32873 & n37560) | (n32873 & n37561) | (n37560 & n37561);
  assign n36463 = n26349 & ~n33303;
  assign n36464 = n26349 & ~n33302;
  assign n36465 = (~n32873 & n36463) | (~n32873 & n36464) | (n36463 & n36464);
  assign n26653 = n36462 & n36465;
  assign n33315 = n26649 | n26653;
  assign n33316 = n33314 | n33315;
  assign n33317 = n26649 & n26653;
  assign n33318 = (n26649 & n33314) | (n26649 & n33317) | (n33314 & n33317);
  assign n26657 = n33316 & ~n33318;
  assign n26658 = x139 & x158;
  assign n26659 = n26657 | n26658;
  assign n26660 = n26657 & n26658;
  assign n26661 = n26659 & ~n26660;
  assign n36466 = n26355 | n26363;
  assign n36467 = n33184 | n36466;
  assign n33320 = n26355 | n33193;
  assign n33321 = (n32927 & n36467) | (n32927 & n33320) | (n36467 & n33320);
  assign n37562 = ~n26355 & n26356;
  assign n37563 = (n26356 & ~n33193) | (n26356 & n37562) | (~n33193 & n37562);
  assign n36469 = n26356 & ~n36432;
  assign n36470 = (~n32927 & n37563) | (~n32927 & n36469) | (n37563 & n36469);
  assign n26664 = n33321 & n36470;
  assign n33322 = n26661 | n26664;
  assign n33323 = n33276 | n33322;
  assign n33324 = n26661 & n26664;
  assign n33325 = (n26661 & n33276) | (n26661 & n33324) | (n33276 & n33324);
  assign n26668 = n33323 & ~n33325;
  assign n26669 = x138 & x159;
  assign n26670 = ~n26668 & n26669;
  assign n26671 = n26668 & ~n26669;
  assign n26672 = n26670 | n26671;
  assign n33326 = n26611 | n26672;
  assign n33327 = n33263 | n33326;
  assign n33328 = n26611 & n26672;
  assign n33329 = (n26672 & n33263) | (n26672 & n33328) | (n33263 & n33328);
  assign n26675 = n33327 & ~n33329;
  assign n26676 = n33270 | n26675;
  assign n26677 = n33270 & n26675;
  assign n26678 = n26676 & ~n26677;
  assign n26679 = n26600 & n26678;
  assign n26680 = n26600 | n26678;
  assign n26681 = ~n26679 & n26680;
  assign n26593 = n26120 & n26393;
  assign n36471 = n26119 & n26120;
  assign n36472 = n26393 & n36471;
  assign n33252 = (n26593 & n33095) | (n26593 & n36472) | (n33095 & n36472);
  assign n33253 = n26312 | n26386;
  assign n33254 = n33080 | n33253;
  assign n33257 = n26387 & ~n33255;
  assign n33258 = ~n26386 & n26387;
  assign n33259 = (~n33080 & n33257) | (~n33080 & n33258) | (n33257 & n33258);
  assign n26598 = n33254 & n33259;
  assign n33330 = n26598 & n26681;
  assign n33331 = (n26681 & n33252) | (n26681 & n33330) | (n33252 & n33330);
  assign n33332 = n26598 | n26681;
  assign n33333 = n33252 | n33332;
  assign n26684 = ~n33331 & n33333;
  assign n26685 = x136 & x161;
  assign n26686 = n26684 & n26685;
  assign n26687 = n26684 | n26685;
  assign n26688 = ~n26686 & n26687;
  assign n26689 = n26119 | n26393;
  assign n33334 = n26121 | n26689;
  assign n33335 = (n26689 & n33095) | (n26689 & n33334) | (n33095 & n33334);
  assign n26691 = ~n33252 & n33335;
  assign n26692 = n26394 & n26691;
  assign n33336 = n26688 | n26692;
  assign n33337 = n33207 | n33336;
  assign n33338 = n26688 & n26692;
  assign n33339 = (n26688 & n33207) | (n26688 & n33338) | (n33207 & n33338);
  assign n26696 = n33337 & ~n33339;
  assign n26697 = n26591 & n26696;
  assign n26698 = n26591 | n26696;
  assign n26699 = ~n26697 & n26698;
  assign n33144 = (n26303 & n33099) | (n26303 & n33143) | (n33099 & n33143);
  assign n26579 = ~n26400 & n26404;
  assign n26580 = n26400 & ~n26404;
  assign n26581 = n26579 | n26580;
  assign n26582 = n33144 | n26581;
  assign n26583 = n33144 & n26581;
  assign n26584 = n26582 & ~n26583;
  assign n26585 = n26149 & n26584;
  assign n33245 = n26148 & n26585;
  assign n33246 = (n26585 & n33104) | (n26585 & n33245) | (n33104 & n33245);
  assign n33340 = n26405 & n26699;
  assign n33341 = (n26699 & n33246) | (n26699 & n33340) | (n33246 & n33340);
  assign n33342 = n26405 | n26699;
  assign n33343 = n33246 | n33342;
  assign n26702 = ~n33341 & n33343;
  assign n26703 = x134 & x163;
  assign n26704 = x133 & x164;
  assign n26705 = n26703 | n26704;
  assign n26706 = n26703 & n26704;
  assign n26707 = n26705 & ~n26706;
  assign n26708 = n26702 | n26707;
  assign n26709 = n26702 & n26707;
  assign n26710 = n26708 & ~n26709;
  assign n26577 = n33141 | n26407;
  assign n33247 = n26408 & ~n33246;
  assign n33248 = n26577 & n33247;
  assign n33249 = n26414 | n33248;
  assign n33344 = n26710 | n33249;
  assign n33345 = n26710 | n33248;
  assign n33346 = (n33139 & n33344) | (n33139 & n33345) | (n33344 & n33345);
  assign n33347 = n26710 & n33249;
  assign n33348 = n26710 & n33248;
  assign n33349 = (n33139 & n33347) | (n33139 & n33348) | (n33347 & n33348);
  assign n26713 = n33346 & ~n33349;
  assign n26714 = x132 & x165;
  assign n26715 = ~n26713 & n26714;
  assign n26716 = n26713 & ~n26714;
  assign n26717 = n26715 | n26716;
  assign n26718 = n33244 | n26717;
  assign n26719 = n33244 & n26717;
  assign n26720 = n26718 & ~n26719;
  assign n26721 = n26566 & n26720;
  assign n26722 = n26566 | n26720;
  assign n26723 = ~n26721 & n26722;
  assign n26575 = n26567 & n26574;
  assign n26724 = n26287 | n26573;
  assign n26725 = n26289 | n26724;
  assign n26726 = ~n26575 & n26725;
  assign n26727 = n26422 & n26726;
  assign n36473 = n26429 | n26727;
  assign n36474 = (n26727 & n33136) | (n26727 & n36473) | (n33136 & n36473);
  assign n26729 = n26723 | n36474;
  assign n26730 = n26723 & n36474;
  assign n26731 = n26729 & ~n26730;
  assign n26732 = x130 & x167;
  assign n26733 = ~n26731 & n26732;
  assign n26734 = n26731 & ~n26732;
  assign n26735 = n26733 | n26734;
  assign n26736 = n36425 | n26735;
  assign n26737 = n36425 & n26735;
  assign n26738 = n26736 & ~n26737;
  assign n26739 = n26564 & n26738;
  assign n26740 = n26564 | n26738;
  assign n26741 = ~n26739 & n26740;
  assign n26742 = n36423 | n26741;
  assign n26743 = n36423 & n26741;
  assign n26744 = n26742 & ~n26743;
  assign n26745 = x128 & x169;
  assign n26746 = n26744 | n26745;
  assign n26747 = n26744 & n26745;
  assign n26748 = n26746 & ~n26747;
  assign n26749 = n33236 | n26748;
  assign n26750 = n33236 & n26748;
  assign n26751 = n26749 & ~n26750;
  assign n26752 = x127 & x170;
  assign n26753 = n26751 | n26752;
  assign n26754 = n26751 & n26752;
  assign n26755 = n26753 & ~n26754;
  assign n26756 = n33233 | n26755;
  assign n26757 = n33233 & n26755;
  assign n26758 = n26756 & ~n26757;
  assign n33350 = ~n26539 & n26758;
  assign n33351 = ~n26532 & n33350;
  assign n33352 = n26539 & ~n26758;
  assign n33353 = (n26532 & ~n26758) | (n26532 & n33352) | (~n26758 & n33352);
  assign n26761 = n33351 | n33353;
  assign n26762 = x126 & x171;
  assign n26763 = n26761 & n26762;
  assign n26764 = n26761 | n26762;
  assign n26765 = ~n26763 & n26764;
  assign n26766 = n33228 & n26765;
  assign n26767 = n33228 | n26765;
  assign n26768 = ~n26766 & n26767;
  assign n26769 = n26528 & n26768;
  assign n26770 = n26528 | n26768;
  assign n26771 = ~n26769 & n26770;
  assign n26772 = n33226 & n26771;
  assign n26773 = n33226 | n26771;
  assign n26774 = ~n26772 & n26773;
  assign n26775 = n26520 & n26774;
  assign n26776 = n26520 | n26774;
  assign n26777 = ~n26775 & n26776;
  assign n26778 = n33220 & n26777;
  assign n26779 = n33220 | n26777;
  assign n26780 = ~n26778 & n26779;
  assign n26781 = n26514 & n26780;
  assign n26782 = n26514 | n26780;
  assign n26783 = ~n26781 & n26782;
  assign n26784 = n33216 & n26783;
  assign n26785 = n33216 | n26783;
  assign n26786 = ~n26784 & n26785;
  assign n26787 = n26508 & n26786;
  assign n26788 = n26508 | n26786;
  assign n26789 = ~n26787 & n26788;
  assign n26790 = n26507 & n26789;
  assign n26791 = n26507 | n26789;
  assign n26792 = ~n26790 & n26791;
  assign n33354 = n26787 | n26789;
  assign n33355 = (n26507 & n26787) | (n26507 & n33354) | (n26787 & n33354);
  assign n26794 = x123 & x175;
  assign n26795 = n26781 | n26784;
  assign n26796 = x124 & x174;
  assign n33356 = n26775 | n26777;
  assign n33357 = (n26775 & n33220) | (n26775 & n33356) | (n33220 & n33356);
  assign n26798 = x125 & x173;
  assign n26799 = n26769 | n26772;
  assign n26800 = x126 & x172;
  assign n33358 = n26763 | n26765;
  assign n33359 = (n26763 & n33228) | (n26763 & n33358) | (n33228 & n33358);
  assign n33365 = n26751 & n33232;
  assign n33366 = n26544 & n26751;
  assign n33367 = (n33130 & n33365) | (n33130 & n33366) | (n33365 & n33366);
  assign n33368 = n26744 & n33235;
  assign n33369 = n26549 & n26744;
  assign n33370 = (n33132 & n33368) | (n33132 & n33369) | (n33368 & n33369);
  assign n33371 = n26744 | n33235;
  assign n33372 = n26549 | n26744;
  assign n33373 = (n33132 & n33371) | (n33132 & n33372) | (n33371 & n33372);
  assign n26810 = n26745 & n33373;
  assign n26811 = ~n33370 & n26810;
  assign n26812 = n33367 | n26811;
  assign n26813 = n26562 | n26738;
  assign n33374 = n26443 | n26813;
  assign n33375 = (n26813 & n33134) | (n26813 & n33374) | (n33134 & n33374);
  assign n26815 = n26206 | n26562;
  assign n33376 = n26210 | n26815;
  assign n33377 = (n25988 & n26815) | (n25988 & n33376) | (n26815 & n33376);
  assign n26817 = n26437 | n26561;
  assign n26818 = n26738 & n26817;
  assign n26819 = n33377 & n26818;
  assign n26820 = n33375 & ~n26819;
  assign n26821 = n26564 & n26820;
  assign n26822 = n33370 | n26821;
  assign n26823 = x129 & x169;
  assign n33378 = n26434 & n26731;
  assign n36475 = (n26559 & n26731) | (n26559 & n33378) | (n26731 & n33378);
  assign n36476 = n26731 & n33378;
  assign n36477 = (n33240 & n36475) | (n33240 & n36476) | (n36475 & n36476);
  assign n33380 = n26434 | n26731;
  assign n33382 = n26732 & n33380;
  assign n33383 = (n26560 & n26732) | (n26560 & n33382) | (n26732 & n33382);
  assign n26827 = ~n36477 & n33383;
  assign n33384 = n26818 | n26827;
  assign n33385 = (n26827 & n33377) | (n26827 & n33384) | (n33377 & n33384);
  assign n33386 = n26720 | n26727;
  assign n33387 = n26430 | n33386;
  assign n26830 = n26292 | n26727;
  assign n26831 = n26196 | n26830;
  assign n26832 = n26422 | n26726;
  assign n26833 = n26720 & n26832;
  assign n26834 = n26831 & n26833;
  assign n26835 = n33387 & ~n26834;
  assign n26836 = n26566 & n26835;
  assign n33388 = n26836 | n33378;
  assign n33389 = n26731 | n26836;
  assign n33390 = (n26560 & n33388) | (n26560 & n33389) | (n33388 & n33389);
  assign n26838 = n33244 & n26713;
  assign n33391 = n26713 & n26714;
  assign n33392 = (n26714 & n33244) | (n26714 & n33391) | (n33244 & n33391);
  assign n26841 = ~n26838 & n33392;
  assign n33393 = n26833 | n26841;
  assign n33394 = (n26831 & n26841) | (n26831 & n33393) | (n26841 & n33393);
  assign n26843 = n26702 | n26703;
  assign n26844 = n26702 & n26703;
  assign n26845 = n26843 & ~n26844;
  assign n33395 = n26845 | n33249;
  assign n33396 = n26845 | n33248;
  assign n33397 = (n33139 & n33395) | (n33139 & n33396) | (n33395 & n33396);
  assign n26590 = n26405 | n33246;
  assign n26849 = ~n26699 & n26703;
  assign n26850 = n26699 & ~n26703;
  assign n26851 = n26849 | n26850;
  assign n26852 = ~n26590 & n26851;
  assign n26853 = n26590 & ~n26851;
  assign n26854 = n26852 | n26853;
  assign n33398 = ~n26408 & n33246;
  assign n33399 = (n26408 & n26577) | (n26408 & ~n33398) | (n26577 & ~n33398);
  assign n36478 = n33248 & n33399;
  assign n36479 = n26854 & n36478;
  assign n36480 = n26704 & ~n36479;
  assign n37564 = n26704 & ~n33399;
  assign n37565 = (n26704 & ~n26854) | (n26704 & n37564) | (~n26854 & n37564);
  assign n36482 = (~n33139 & n36480) | (~n33139 & n37565) | (n36480 & n37565);
  assign n26858 = n33397 & n36482;
  assign n33402 = n26713 | n26858;
  assign n33403 = (n26858 & n33244) | (n26858 & n33402) | (n33244 & n33402);
  assign n36483 = n26844 | n36479;
  assign n26855 = n33399 & n26854;
  assign n36484 = n26844 | n26855;
  assign n36485 = (n33139 & n36483) | (n33139 & n36484) | (n36483 & n36484);
  assign n26861 = n26303 | n26692;
  assign n33404 = n26144 | n26861;
  assign n33405 = (n26861 & n33099) | (n26861 & n33404) | (n33099 & n33404);
  assign n26863 = n26394 | n26691;
  assign n33406 = n26688 & n26863;
  assign n33407 = n33405 & n33406;
  assign n26866 = n33337 & ~n33407;
  assign n26867 = n26591 & n26866;
  assign n26868 = n33341 | n26867;
  assign n26869 = x135 & x163;
  assign n26870 = n26686 | n33407;
  assign n33410 = ~n26379 & n33263;
  assign n33411 = (n26379 & n33265) | (n26379 & ~n33410) | (n33265 & ~n33410);
  assign n26873 = n26675 & n33411;
  assign n33408 = n26312 | n33267;
  assign n33412 = n26873 & n33408;
  assign n33413 = (n26873 & n33080) | (n26873 & n33412) | (n33080 & n33412);
  assign n33414 = n26600 & ~n33413;
  assign n33415 = n26676 & n33414;
  assign n33418 = n26611 & n26668;
  assign n33419 = (n26668 & n33263) | (n26668 & n33418) | (n33263 & n33418);
  assign n36486 = n26611 & n26669;
  assign n36487 = (n26668 & n26669) | (n26668 & n36486) | (n26669 & n36486);
  assign n33423 = (n26669 & n33263) | (n26669 & n36487) | (n33263 & n36487);
  assign n26881 = ~n33419 & n33423;
  assign n26888 = x140 & x158;
  assign n26894 = x141 & x157;
  assign n26900 = x142 & x156;
  assign n26907 = x143 & x155;
  assign n33451 = n26617 & n26624;
  assign n36488 = n26907 & n36444;
  assign n36489 = (n26907 & n33451) | (n26907 & n36488) | (n33451 & n36488);
  assign n36490 = (n26624 & n26907) | (n26624 & n36488) | (n26907 & n36488);
  assign n36491 = (n33278 & n36489) | (n33278 & n36490) | (n36489 & n36490);
  assign n36492 = (n33277 & n36489) | (n33277 & n36490) | (n36489 & n36490);
  assign n36493 = (n33009 & n36491) | (n33009 & n36492) | (n36491 & n36492);
  assign n36494 = n26907 | n36444;
  assign n36495 = n33451 | n36494;
  assign n36496 = n26624 | n36494;
  assign n36497 = (n33278 & n36495) | (n33278 & n36496) | (n36495 & n36496);
  assign n36498 = (n33277 & n36495) | (n33277 & n36496) | (n36495 & n36496);
  assign n36499 = (n33009 & n36497) | (n33009 & n36498) | (n36497 & n36498);
  assign n26910 = ~n36493 & n36499;
  assign n37566 = (n26341 & n26624) | (n26341 & n33451) | (n26624 & n33451);
  assign n37567 = n26624 & n33451;
  assign n37568 = (n33167 & n37566) | (n33167 & n37567) | (n37566 & n37567);
  assign n36501 = (n26624 & n33277) | (n26624 & n33451) | (n33277 & n33451);
  assign n36502 = (n33009 & n37568) | (n33009 & n36501) | (n37568 & n36501);
  assign n33453 = n26617 | n26624;
  assign n33455 = n26619 & n33453;
  assign n36503 = (n26619 & n33278) | (n26619 & n33455) | (n33278 & n33455);
  assign n36504 = (n26619 & n33277) | (n26619 & n33455) | (n33277 & n33455);
  assign n36505 = (n33009 & n36503) | (n33009 & n36504) | (n36503 & n36504);
  assign n26904 = ~n36502 & n36505;
  assign n33458 = n26630 | n26904;
  assign n33470 = n26910 & n33458;
  assign n33442 = n26630 & n26641;
  assign n36506 = n26904 & n26910;
  assign n36507 = (n26910 & n33442) | (n26910 & n36506) | (n33442 & n36506);
  assign n36508 = (n33303 & n33470) | (n33303 & n36507) | (n33470 & n36507);
  assign n36509 = (n33302 & n33470) | (n33302 & n36507) | (n33470 & n36507);
  assign n36510 = (n32873 & n36508) | (n32873 & n36509) | (n36508 & n36509);
  assign n33473 = n26910 | n33458;
  assign n36511 = n26904 | n26910;
  assign n36512 = n33442 | n36511;
  assign n36513 = (n33303 & n33473) | (n33303 & n36512) | (n33473 & n36512);
  assign n36514 = (n33302 & n33473) | (n33302 & n36512) | (n33473 & n36512);
  assign n36515 = (n32873 & n36513) | (n32873 & n36514) | (n36513 & n36514);
  assign n26913 = ~n36510 & n36515;
  assign n26914 = n26900 & n26913;
  assign n26915 = n26900 | n26913;
  assign n26916 = ~n26914 & n26915;
  assign n36516 = (n26630 & n33303) | (n26630 & n33442) | (n33303 & n33442);
  assign n36517 = (n26630 & n33302) | (n26630 & n33442) | (n33302 & n33442);
  assign n36518 = (n32873 & n36516) | (n32873 & n36517) | (n36516 & n36517);
  assign n33444 = n26630 | n26641;
  assign n33446 = n26631 & n33444;
  assign n36519 = (n26631 & n33303) | (n26631 & n33446) | (n33303 & n33446);
  assign n36520 = (n26631 & n33302) | (n26631 & n33446) | (n33302 & n33446);
  assign n36521 = (n32873 & n36519) | (n32873 & n36520) | (n36519 & n36520);
  assign n26898 = ~n36518 & n36521;
  assign n36522 = n26653 | n26898;
  assign n36523 = (n26645 & n26898) | (n26645 & n36522) | (n26898 & n36522);
  assign n33475 = n26916 & n36523;
  assign n33449 = n26645 | n26898;
  assign n33476 = n26916 & n33449;
  assign n33477 = (n33314 & n33475) | (n33314 & n33476) | (n33475 & n33476);
  assign n33478 = n26916 | n36523;
  assign n33479 = n26916 | n33449;
  assign n33480 = (n33314 & n33478) | (n33314 & n33479) | (n33478 & n33479);
  assign n26919 = ~n33477 & n33480;
  assign n26920 = n26894 & n26919;
  assign n26921 = n26894 | n26919;
  assign n26922 = ~n26920 & n26921;
  assign n33433 = n26645 & n26653;
  assign n36524 = (n26645 & n33313) | (n26645 & n33433) | (n33313 & n33433);
  assign n36525 = (n26645 & n33433) | (n26645 & n36432) | (n33433 & n36432);
  assign n36526 = (n32927 & n36524) | (n32927 & n36525) | (n36524 & n36525);
  assign n36527 = n26646 & n26653;
  assign n36528 = (n26645 & n26646) | (n26645 & n36527) | (n26646 & n36527);
  assign n36529 = (n26646 & n33313) | (n26646 & n36528) | (n33313 & n36528);
  assign n36530 = (n26646 & n36432) | (n26646 & n36528) | (n36432 & n36528);
  assign n36531 = (n32927 & n36529) | (n32927 & n36530) | (n36529 & n36530);
  assign n26892 = ~n36526 & n36531;
  assign n36532 = n26664 | n26892;
  assign n36533 = (n26657 & n26892) | (n26657 & n36532) | (n26892 & n36532);
  assign n33481 = n26922 & n36533;
  assign n33440 = n26657 | n26892;
  assign n33482 = n26922 & n33440;
  assign n33483 = (n33276 & n33481) | (n33276 & n33482) | (n33481 & n33482);
  assign n33484 = n26922 | n36533;
  assign n33485 = n26922 | n33440;
  assign n33486 = (n33276 & n33484) | (n33276 & n33485) | (n33484 & n33485);
  assign n26925 = ~n33483 & n33486;
  assign n26926 = n26888 | n26925;
  assign n26927 = n26888 & n26925;
  assign n26928 = n26926 & ~n26927;
  assign n33424 = n26657 & n26664;
  assign n36534 = (n26657 & n33424) | (n26657 & n36427) | (n33424 & n36427);
  assign n36535 = (n26657 & n33275) | (n26657 & n33424) | (n33275 & n33424);
  assign n36536 = (n33006 & n36534) | (n33006 & n36535) | (n36534 & n36535);
  assign n36537 = n26658 & n26664;
  assign n36538 = (n26657 & n26658) | (n26657 & n36537) | (n26658 & n36537);
  assign n36539 = (n26658 & n36427) | (n26658 & n36538) | (n36427 & n36538);
  assign n36540 = (n26658 & n33275) | (n26658 & n36538) | (n33275 & n36538);
  assign n36541 = (n33006 & n36539) | (n33006 & n36540) | (n36539 & n36540);
  assign n26886 = ~n36536 & n36541;
  assign n36542 = n26611 | n26886;
  assign n36543 = (n26668 & n26886) | (n26668 & n36542) | (n26886 & n36542);
  assign n33487 = n26928 | n36543;
  assign n33431 = n26668 | n26886;
  assign n33488 = n26928 | n33431;
  assign n33489 = (n33263 & n33487) | (n33263 & n33488) | (n33487 & n33488);
  assign n33490 = n26928 & n36543;
  assign n33491 = n26928 & n33431;
  assign n33492 = (n33263 & n33490) | (n33263 & n33491) | (n33490 & n33491);
  assign n26931 = n33489 & ~n33492;
  assign n26932 = x139 & x159;
  assign n26933 = x138 & x160;
  assign n26934 = n26932 & n26933;
  assign n26935 = n26932 | n26933;
  assign n26936 = ~n26934 & n26935;
  assign n26937 = n26931 & ~n26936;
  assign n26938 = ~n26931 & n26936;
  assign n26939 = n26937 | n26938;
  assign n33493 = n26881 | n26939;
  assign n33494 = n33413 | n33493;
  assign n33495 = n26881 & n26939;
  assign n33496 = (n26939 & n33413) | (n26939 & n33495) | (n33413 & n33495);
  assign n26942 = n33494 & ~n33496;
  assign n26946 = n33415 | n26942;
  assign n26947 = n33331 | n26946;
  assign n26949 = x137 & x161;
  assign n33497 = ~n26600 & n33413;
  assign n33498 = (n26600 & n26676) | (n26600 & ~n33497) | (n26676 & ~n33497);
  assign n26944 = n26942 & n33498;
  assign n33416 = n26598 | n33415;
  assign n33499 = n26944 & n33416;
  assign n36544 = n26949 & ~n33499;
  assign n36545 = ~n26944 & n26949;
  assign n36546 = (~n33252 & n36544) | (~n33252 & n36545) | (n36544 & n36545);
  assign n33502 = n26947 & n36546;
  assign n36547 = ~n26949 & n33499;
  assign n36548 = n26944 & ~n26949;
  assign n36549 = (n33252 & n36547) | (n33252 & n36548) | (n36547 & n36548);
  assign n33504 = (n26947 & n26949) | (n26947 & ~n36549) | (n26949 & ~n36549);
  assign n26952 = ~n33502 & n33504;
  assign n26953 = x136 & x162;
  assign n26954 = n26952 & ~n26953;
  assign n26955 = ~n26952 & n26953;
  assign n26956 = n26954 | n26955;
  assign n26957 = n26870 & n26956;
  assign n26958 = n26870 | n26956;
  assign n26959 = ~n26957 & n26958;
  assign n26960 = n26869 & n26959;
  assign n26961 = n26869 | n26959;
  assign n26962 = ~n26960 & n26961;
  assign n26963 = n26868 | n26962;
  assign n26964 = n26868 & n26962;
  assign n26965 = n26963 & ~n26964;
  assign n26966 = x134 & x164;
  assign n26967 = n26965 | n26966;
  assign n26968 = n26965 & n26966;
  assign n26969 = n26967 & ~n26968;
  assign n26970 = ~n36485 & n26969;
  assign n26971 = n36485 & ~n26969;
  assign n26972 = n26970 | n26971;
  assign n26973 = x133 & x165;
  assign n26974 = n26972 & n26973;
  assign n26975 = n26972 | n26973;
  assign n26976 = ~n26974 & n26975;
  assign n26977 = n33403 | n26976;
  assign n26978 = n33403 & n26976;
  assign n26979 = n26977 & ~n26978;
  assign n26980 = n33394 & n26979;
  assign n26981 = n33394 | n26979;
  assign n26982 = ~n26980 & n26981;
  assign n26983 = x132 & x166;
  assign n26984 = n26982 & n26983;
  assign n26985 = n26982 | n26983;
  assign n26986 = ~n26984 & n26985;
  assign n26987 = x131 & x167;
  assign n26988 = n26986 & n26987;
  assign n26989 = n26986 | n26987;
  assign n26990 = ~n26988 & n26989;
  assign n26991 = n33390 | n26990;
  assign n26992 = n33390 & n26990;
  assign n26993 = n26991 & ~n26992;
  assign n26994 = x130 & x168;
  assign n26995 = ~n26993 & n26994;
  assign n26996 = n26993 & ~n26994;
  assign n26997 = n26995 | n26996;
  assign n26998 = n33385 | n26997;
  assign n26999 = n33385 & n26997;
  assign n27000 = n26998 & ~n26999;
  assign n27001 = n26823 & n27000;
  assign n27002 = n26823 | n27000;
  assign n27003 = ~n27001 & n27002;
  assign n27004 = n26822 | n27003;
  assign n27005 = n26822 & n27003;
  assign n27006 = n27004 & ~n27005;
  assign n27007 = x128 & x170;
  assign n27008 = n27006 | n27007;
  assign n27009 = n27006 & n27007;
  assign n27010 = n27008 & ~n27009;
  assign n27011 = n26812 | n27010;
  assign n27012 = n26812 & n27010;
  assign n27013 = n27011 & ~n27012;
  assign n33360 = n26539 & n26758;
  assign n33361 = (n26532 & n26758) | (n26532 & n33360) | (n26758 & n33360);
  assign n33362 = n26751 | n33232;
  assign n33363 = n26544 | n26751;
  assign n33364 = (n33130 & n33362) | (n33130 & n33363) | (n33362 & n33363);
  assign n26805 = n26752 & ~n33367;
  assign n26806 = n33364 & n26805;
  assign n33505 = n26806 & n27013;
  assign n33506 = (n27013 & n33361) | (n27013 & n33505) | (n33361 & n33505);
  assign n33507 = n26806 | n27013;
  assign n33508 = n33361 | n33507;
  assign n27016 = ~n33506 & n33508;
  assign n27017 = x127 & x171;
  assign n27018 = n27016 & n27017;
  assign n27019 = n27016 | n27017;
  assign n27020 = ~n27018 & n27019;
  assign n27021 = n33359 & n27020;
  assign n27022 = n33359 | n27020;
  assign n27023 = ~n27021 & n27022;
  assign n27024 = n26800 & n27023;
  assign n27025 = n26800 | n27023;
  assign n27026 = ~n27024 & n27025;
  assign n27027 = n26799 & n27026;
  assign n27028 = n26799 | n27026;
  assign n27029 = ~n27027 & n27028;
  assign n27030 = n26798 & n27029;
  assign n27031 = n26798 | n27029;
  assign n27032 = ~n27030 & n27031;
  assign n27033 = n33357 & n27032;
  assign n27034 = n33357 | n27032;
  assign n27035 = ~n27033 & n27034;
  assign n27036 = n26796 & n27035;
  assign n27037 = n26796 | n27035;
  assign n27038 = ~n27036 & n27037;
  assign n27039 = n26795 & n27038;
  assign n27040 = n26795 | n27038;
  assign n27041 = ~n27039 & n27040;
  assign n27042 = n26794 & n27041;
  assign n27043 = n26794 | n27041;
  assign n27044 = ~n27042 & n27043;
  assign n27045 = n33355 & n27044;
  assign n27046 = n33355 | n27044;
  assign n27047 = ~n27045 & n27046;
  assign n27048 = n27042 | n27045;
  assign n27049 = x124 & x175;
  assign n33509 = n27036 | n27038;
  assign n33510 = (n26795 & n27036) | (n26795 & n33509) | (n27036 & n33509);
  assign n27051 = x125 & x174;
  assign n27052 = n27030 | n27033;
  assign n27053 = x126 & x173;
  assign n33511 = n27024 | n27026;
  assign n33512 = (n26799 & n27024) | (n26799 & n33511) | (n27024 & n33511);
  assign n33513 = n27018 | n27020;
  assign n33514 = (n27018 & n33359) | (n27018 & n33513) | (n33359 & n33513);
  assign n33517 = n26811 & n27006;
  assign n33518 = (n27006 & n33367) | (n27006 & n33517) | (n33367 & n33517);
  assign n27061 = n26821 | n27000;
  assign n27062 = n33370 | n27061;
  assign n27065 = n26564 | n26820;
  assign n27066 = n27000 & n27065;
  assign n36550 = n26549 | n26564;
  assign n36551 = (n26549 & n26820) | (n26549 & n36550) | (n26820 & n36550);
  assign n33519 = n36551 & n27066;
  assign n33520 = (n26541 & n27066) | (n26541 & n33519) | (n27066 & n33519);
  assign n27068 = n27062 & ~n33520;
  assign n27069 = n26823 & n27068;
  assign n27070 = n33518 | n27069;
  assign n27071 = x129 & x170;
  assign n36552 = n26993 & n33384;
  assign n36553 = n26827 & n26993;
  assign n36554 = (n33377 & n36552) | (n33377 & n36553) | (n36552 & n36553);
  assign n33521 = n26993 & n26994;
  assign n33522 = (n26994 & n33385) | (n26994 & n33521) | (n33385 & n33521);
  assign n27075 = ~n36554 & n33522;
  assign n27076 = n33520 | n27075;
  assign n27077 = n33390 | n26986;
  assign n33523 = n26434 | n26836;
  assign n33524 = n26560 | n33523;
  assign n27079 = n26566 | n26835;
  assign n27080 = n26986 & n27079;
  assign n27081 = n33524 & n27080;
  assign n27082 = n27077 & ~n27081;
  assign n27083 = n26987 & n27082;
  assign n27084 = n26984 | n27081;
  assign n27085 = x132 & x167;
  assign n27086 = x133 & x166;
  assign n27087 = n26419 | n26858;
  assign n36555 = n26574 | n27087;
  assign n36556 = (n26567 & n27087) | (n26567 & n36555) | (n27087 & n36555);
  assign n33401 = (n26855 & n33139) | (n26855 & n36479) | (n33139 & n36479);
  assign n33525 = n26844 & n26965;
  assign n33526 = (n26965 & n33401) | (n26965 & n33525) | (n33401 & n33525);
  assign n37569 = n26703 & n26966;
  assign n37570 = n26702 & n37569;
  assign n36558 = (n26965 & n26966) | (n26965 & n37570) | (n26966 & n37570);
  assign n33530 = (n26966 & n33401) | (n26966 & n36558) | (n33401 & n36558);
  assign n27096 = ~n33526 & n33530;
  assign n27089 = n33397 & ~n33401;
  assign n27090 = n26704 | n27089;
  assign n27091 = n26972 & n27090;
  assign n33531 = n27091 | n27096;
  assign n33532 = (n36556 & n27096) | (n36556 & n33531) | (n27096 & n33531);
  assign n33533 = n26867 | n26959;
  assign n33534 = n33341 | n33533;
  assign n27099 = n26405 | n26867;
  assign n27100 = n33246 | n27099;
  assign n27101 = n26591 | n26866;
  assign n27102 = n26959 & n27101;
  assign n27103 = n27100 & n27102;
  assign n27104 = n33534 & ~n27103;
  assign n27105 = n26869 & n27104;
  assign n33535 = n26844 | n27105;
  assign n33536 = n33401 | n33535;
  assign n27107 = n26931 & n26932;
  assign n27108 = n26931 | n26932;
  assign n27109 = ~n27107 & n27108;
  assign n33537 = n26881 & n27109;
  assign n33538 = (n27109 & n33413) | (n27109 & n33537) | (n33413 & n33537);
  assign n33539 = n26881 | n27109;
  assign n33540 = n33413 | n33539;
  assign n27112 = n26933 & n33540;
  assign n27113 = ~n33538 & n27112;
  assign n33541 = n27113 | n33499;
  assign n33542 = n26944 | n27113;
  assign n33543 = (n33252 & n33541) | (n33252 & n33542) | (n33541 & n33542);
  assign n27119 = x142 & x157;
  assign n27121 = x143 & x156;
  assign n33547 = n27121 & n36493;
  assign n33548 = (n27121 & n36510) | (n27121 & n33547) | (n36510 & n33547);
  assign n33549 = n27121 | n36493;
  assign n33550 = n36510 | n33549;
  assign n27124 = ~n33548 & n33550;
  assign n27125 = n27119 & n27124;
  assign n27126 = n27119 | n27124;
  assign n27127 = ~n27125 & n27126;
  assign n33551 = n26914 | n27127;
  assign n33552 = n33477 | n33551;
  assign n33553 = n26914 & n27127;
  assign n33554 = (n27127 & n33477) | (n27127 & n33553) | (n33477 & n33553);
  assign n27130 = n33552 & ~n33554;
  assign n27131 = x141 & x158;
  assign n27132 = ~n27130 & n27131;
  assign n27133 = n27130 & ~n27131;
  assign n27134 = n27132 | n27133;
  assign n33555 = n26920 | n27134;
  assign n33556 = n33483 | n33555;
  assign n33557 = n26920 & n27134;
  assign n33558 = (n27134 & n33483) | (n27134 & n33557) | (n33483 & n33557);
  assign n27137 = n33556 & ~n33558;
  assign n27140 = n26927 | n27137;
  assign n27141 = n33492 | n27140;
  assign n27143 = x140 & x159;
  assign n27144 = x139 & x160;
  assign n27145 = n27143 & n27144;
  assign n27146 = n27143 | n27144;
  assign n27147 = ~n27145 & n27146;
  assign n27138 = n26926 & n27137;
  assign n33545 = n26927 | n33431;
  assign n36559 = n27138 & n33545;
  assign n33544 = n26927 | n36543;
  assign n36560 = n27138 & n33544;
  assign n36561 = (n33263 & n36559) | (n33263 & n36560) | (n36559 & n36560);
  assign n36562 = n27147 & ~n36561;
  assign n36563 = n27141 & n36562;
  assign n36564 = ~n27147 & n36561;
  assign n36565 = (n27141 & n27147) | (n27141 & ~n36564) | (n27147 & ~n36564);
  assign n27150 = ~n36563 & n36565;
  assign n33559 = n27107 | n27150;
  assign n33560 = n33538 | n33559;
  assign n33561 = n27107 & n27150;
  assign n33562 = (n27150 & n33538) | (n27150 & n33561) | (n33538 & n33561);
  assign n27153 = n33560 & ~n33562;
  assign n27154 = n33543 | n27153;
  assign n27155 = n33543 & n27153;
  assign n27156 = n27154 & ~n27155;
  assign n27157 = x138 & x161;
  assign n27158 = n27156 & n27157;
  assign n27159 = n27156 | n27157;
  assign n27160 = ~n27158 & n27159;
  assign n33563 = n26686 | n33502;
  assign n33565 = n33504 & n33563;
  assign n33567 = n27160 & n33565;
  assign n33568 = n27160 & n33504;
  assign n33569 = (n33407 & n33567) | (n33407 & n33568) | (n33567 & n33568);
  assign n33570 = n27160 | n33565;
  assign n33571 = n27160 | n33504;
  assign n33572 = (n33407 & n33570) | (n33407 & n33571) | (n33570 & n33571);
  assign n27165 = ~n33569 & n33572;
  assign n27166 = x137 & x162;
  assign n27167 = n27165 & n27166;
  assign n27168 = n27165 | n27166;
  assign n27169 = ~n27167 & n27168;
  assign n33573 = n26686 & n26952;
  assign n33574 = (n26952 & n33407) | (n26952 & n33573) | (n33407 & n33573);
  assign n37571 = n26685 & n26953;
  assign n37572 = n26684 & n37571;
  assign n36567 = (n26952 & n26953) | (n26952 & n37572) | (n26953 & n37572);
  assign n33578 = (n26953 & n33407) | (n26953 & n36567) | (n33407 & n36567);
  assign n27173 = ~n33574 & n33578;
  assign n36568 = n27101 | n27173;
  assign n36569 = (n26959 & n27173) | (n26959 & n36568) | (n27173 & n36568);
  assign n36570 = n27169 & ~n36569;
  assign n36571 = n27169 & ~n27173;
  assign n36572 = (~n27100 & n36570) | (~n27100 & n36571) | (n36570 & n36571);
  assign n36573 = ~n27169 & n36569;
  assign n36574 = ~n27169 & n27173;
  assign n36575 = (n27100 & n36573) | (n27100 & n36574) | (n36573 & n36574);
  assign n27177 = n36572 | n36575;
  assign n27178 = x136 & x163;
  assign n27179 = n27177 & n27178;
  assign n27180 = n27177 | n27178;
  assign n27181 = ~n27179 & n27180;
  assign n27182 = n26869 | n27104;
  assign n27183 = n27181 & n27182;
  assign n27184 = n33536 & n27183;
  assign n27185 = n27105 | n27181;
  assign n27186 = n33526 | n27185;
  assign n27187 = ~n27184 & n27186;
  assign n27188 = x135 & x164;
  assign n27189 = n27187 & n27188;
  assign n27190 = n27187 | n27188;
  assign n27191 = ~n27189 & n27190;
  assign n27192 = n33532 & n27191;
  assign n27193 = n33532 | n27191;
  assign n27194 = ~n27192 & n27193;
  assign n27195 = x134 & x165;
  assign n27196 = n27194 & n27195;
  assign n27197 = n27194 | n27195;
  assign n27198 = ~n27196 & n27197;
  assign n27092 = n36556 & n27091;
  assign n37573 = n26858 & n26973;
  assign n37574 = (n26972 & n26973) | (n26972 & n37573) | (n26973 & n37573);
  assign n33581 = n26972 | n33402;
  assign n36577 = n26973 & n33581;
  assign n36578 = (n33244 & n37574) | (n33244 & n36577) | (n37574 & n36577);
  assign n33585 = ~n27092 & n36578;
  assign n33586 = n26979 | n33585;
  assign n33587 = (n33394 & n33585) | (n33394 & n33586) | (n33585 & n33586);
  assign n27203 = n27198 | n33587;
  assign n27204 = n27198 & n33587;
  assign n27205 = n27203 & ~n27204;
  assign n27206 = n27086 & n27205;
  assign n27207 = n27086 | n27205;
  assign n27208 = ~n27206 & n27207;
  assign n27209 = n27085 | n27208;
  assign n27210 = n27085 & n27208;
  assign n27211 = n27209 & ~n27210;
  assign n27212 = ~n27084 & n27211;
  assign n27213 = n27084 & ~n27211;
  assign n27214 = n27212 | n27213;
  assign n27215 = n27083 | n27214;
  assign n27216 = n36554 | n27215;
  assign n36579 = n27083 | n33384;
  assign n37792 = ~n26987 & n36477;
  assign n37793 = (n26987 & n33383) | (n26987 & ~n37792) | (n33383 & ~n37792);
  assign n37576 = (n26827 & n27082) | (n26827 & n37793) | (n27082 & n37793);
  assign n36581 = (n33377 & n36579) | (n33377 & n37576) | (n36579 & n37576);
  assign n27218 = n26987 | n27082;
  assign n27219 = n27214 & n27218;
  assign n27220 = n36581 & n27219;
  assign n27221 = n27216 & ~n27220;
  assign n27222 = x131 & x168;
  assign n27223 = n27221 & n27222;
  assign n27224 = n27221 | n27222;
  assign n27225 = ~n27223 & n27224;
  assign n27226 = x130 & x169;
  assign n27227 = n27225 & ~n27226;
  assign n27228 = ~n27225 & n27226;
  assign n27229 = n27227 | n27228;
  assign n27230 = n27076 | n27229;
  assign n27231 = n27076 & n27229;
  assign n27232 = n27230 & ~n27231;
  assign n27233 = n27071 & n27232;
  assign n27234 = n27071 | n27232;
  assign n27235 = ~n27233 & n27234;
  assign n27236 = n27070 | n27235;
  assign n27237 = n27070 & n27235;
  assign n27238 = n27236 & ~n27237;
  assign n33515 = n26811 | n27006;
  assign n33516 = n33367 | n33515;
  assign n27058 = n27007 & ~n33518;
  assign n27059 = n33516 & n27058;
  assign n36582 = n27059 & n27238;
  assign n36583 = (n27238 & n33506) | (n27238 & n36582) | (n33506 & n36582);
  assign n36584 = n27059 | n27238;
  assign n36585 = n33506 | n36584;
  assign n27241 = ~n36583 & n36585;
  assign n27242 = x128 & x171;
  assign n27243 = n27241 & n27242;
  assign n27244 = n27241 | n27242;
  assign n27245 = ~n27243 & n27244;
  assign n27246 = n33514 & n27245;
  assign n27247 = n33514 | n27245;
  assign n27248 = ~n27246 & n27247;
  assign n27249 = x127 & x172;
  assign n27250 = n27248 & n27249;
  assign n27251 = n27248 | n27249;
  assign n27252 = ~n27250 & n27251;
  assign n27253 = n33512 & n27252;
  assign n27254 = n33512 | n27252;
  assign n27255 = ~n27253 & n27254;
  assign n27256 = n27053 & n27255;
  assign n27257 = n27053 | n27255;
  assign n27258 = ~n27256 & n27257;
  assign n27259 = n27052 & n27258;
  assign n27260 = n27052 | n27258;
  assign n27261 = ~n27259 & n27260;
  assign n27262 = n27051 & n27261;
  assign n27263 = n27051 | n27261;
  assign n27264 = ~n27262 & n27263;
  assign n27265 = n33510 & n27264;
  assign n27266 = n33510 | n27264;
  assign n27267 = ~n27265 & n27266;
  assign n27268 = n27049 & n27267;
  assign n27269 = n27049 | n27267;
  assign n27270 = ~n27268 & n27269;
  assign n27271 = n27048 & n27270;
  assign n27272 = n27048 | n27270;
  assign n27273 = ~n27271 & n27272;
  assign n33588 = n27268 | n27270;
  assign n33589 = (n27048 & n27268) | (n27048 & n33588) | (n27268 & n33588);
  assign n27275 = x125 & x175;
  assign n27276 = n27262 | n27265;
  assign n27277 = x126 & x174;
  assign n33590 = n27256 | n27258;
  assign n33591 = (n27052 & n27256) | (n27052 & n33590) | (n27256 & n33590);
  assign n27279 = x127 & x173;
  assign n33592 = n27250 | n27252;
  assign n33593 = (n27250 & n33512) | (n27250 & n33592) | (n33512 & n33592);
  assign n27281 = x128 & x172;
  assign n36586 = n27243 | n27245;
  assign n36587 = (n27243 & n33514) | (n27243 & n36586) | (n33514 & n36586);
  assign n27060 = n33506 | n27059;
  assign n27287 = n26823 | n27068;
  assign n27288 = n27232 & n27287;
  assign n36588 = n27075 & n27225;
  assign n36589 = (n27225 & n33520) | (n27225 & n36588) | (n33520 & n36588);
  assign n33598 = n27225 & n27226;
  assign n33599 = (n27076 & n27226) | (n27076 & n33598) | (n27226 & n33598);
  assign n27296 = ~n36589 & n33599;
  assign n27285 = n26811 | n27069;
  assign n27286 = n33367 | n27285;
  assign n33600 = n27286 | n27296;
  assign n33601 = (n27288 & n27296) | (n27288 & n33600) | (n27296 & n33600);
  assign n33602 = n26984 & n27208;
  assign n33603 = (n27081 & n27208) | (n27081 & n33602) | (n27208 & n33602);
  assign n33604 = n26984 | n27208;
  assign n33605 = n27081 | n33604;
  assign n27300 = n27085 & n33605;
  assign n27301 = ~n33603 & n27300;
  assign n33606 = n27219 | n27301;
  assign n33607 = (n36581 & n27301) | (n36581 & n33606) | (n27301 & n33606);
  assign n27303 = n33532 | n27189;
  assign n37577 = n27179 | n27182;
  assign n37578 = (n27179 & n27181) | (n27179 & n37577) | (n27181 & n37577);
  assign n36591 = (n27179 & n33536) | (n27179 & n37578) | (n33536 & n37578);
  assign n36592 = n27143 & ~n36561;
  assign n36593 = n27141 & n36592;
  assign n33608 = n27107 | n36593;
  assign n33609 = n33538 | n33608;
  assign n33546 = (n33263 & n33544) | (n33263 & n33545) | (n33544 & n33545);
  assign n33610 = n26920 & n27130;
  assign n33611 = (n27130 & n33483) | (n27130 & n33610) | (n33483 & n33610);
  assign n33612 = n26920 | n27130;
  assign n33614 = n27131 & n33612;
  assign n33615 = (n27131 & n33483) | (n27131 & n33614) | (n33483 & n33614);
  assign n27311 = ~n33611 & n33615;
  assign n27318 = x142 & x158;
  assign n27320 = x143 & x157;
  assign n33618 = n26914 & n27124;
  assign n37580 = n27121 & n27320;
  assign n37794 = n36493 & n37580;
  assign n37581 = (n36510 & n37794) | (n36510 & n37580) | (n37794 & n37580);
  assign n36595 = (n27320 & n33618) | (n27320 & n37581) | (n33618 & n37581);
  assign n36596 = (n27124 & n27320) | (n27124 & n37581) | (n27320 & n37581);
  assign n36597 = (n33476 & n36595) | (n33476 & n36596) | (n36595 & n36596);
  assign n36598 = (n33475 & n36595) | (n33475 & n36596) | (n36595 & n36596);
  assign n36599 = (n33314 & n36597) | (n33314 & n36598) | (n36597 & n36598);
  assign n37583 = n27121 | n27320;
  assign n37795 = (n27320 & n36493) | (n27320 & n37583) | (n36493 & n37583);
  assign n37584 = (n36510 & n37795) | (n36510 & n37583) | (n37795 & n37583);
  assign n36601 = n33618 | n37584;
  assign n36602 = n27124 | n37584;
  assign n36603 = (n33476 & n36601) | (n33476 & n36602) | (n36601 & n36602);
  assign n36604 = (n33475 & n36601) | (n33475 & n36602) | (n36601 & n36602);
  assign n36605 = (n33314 & n36603) | (n33314 & n36604) | (n36603 & n36604);
  assign n27323 = ~n36599 & n36605;
  assign n27324 = n27318 & n27323;
  assign n27325 = n27318 | n27323;
  assign n27326 = ~n27324 & n27325;
  assign n36606 = (n27124 & n33476) | (n27124 & n33618) | (n33476 & n33618);
  assign n36607 = (n27124 & n33475) | (n27124 & n33618) | (n33475 & n33618);
  assign n36608 = (n33314 & n36606) | (n33314 & n36607) | (n36606 & n36607);
  assign n33620 = n26914 | n27124;
  assign n33622 = n27119 & n33620;
  assign n36609 = (n27119 & n33476) | (n27119 & n33622) | (n33476 & n33622);
  assign n36610 = (n27119 & n33475) | (n27119 & n33622) | (n33475 & n33622);
  assign n36611 = (n33314 & n36609) | (n33314 & n36610) | (n36609 & n36610);
  assign n27316 = ~n36608 & n36611;
  assign n33624 = n27316 | n33610;
  assign n33636 = n27326 | n33624;
  assign n33625 = n27130 | n27316;
  assign n33637 = n27326 | n33625;
  assign n33638 = (n33483 & n33636) | (n33483 & n33637) | (n33636 & n33637);
  assign n33639 = n27326 & n33624;
  assign n33640 = n27326 & n33625;
  assign n33641 = (n33483 & n33639) | (n33483 & n33640) | (n33639 & n33640);
  assign n27329 = n33638 & ~n33641;
  assign n33643 = ~n27311 & n27329;
  assign n36612 = ~n27138 & n33643;
  assign n33644 = (~n33546 & n36612) | (~n33546 & n33643) | (n36612 & n33643);
  assign n33646 = n27311 & ~n27329;
  assign n36613 = (n27138 & ~n27329) | (n27138 & n33646) | (~n27329 & n33646);
  assign n33647 = (n33546 & n36613) | (n33546 & n33646) | (n36613 & n33646);
  assign n27332 = n33644 | n33647;
  assign n27333 = x141 & x159;
  assign n27334 = n27332 & n27333;
  assign n27335 = n27332 | n27333;
  assign n27336 = ~n27334 & n27335;
  assign n36614 = ~n27143 & n36561;
  assign n36615 = (n27141 & n27143) | (n27141 & ~n36614) | (n27143 & ~n36614);
  assign n27338 = n27336 & n36615;
  assign n27339 = n33609 & n27338;
  assign n27340 = ~n36593 & n36615;
  assign n33648 = n27107 & n27340;
  assign n33649 = (n27340 & n33538) | (n27340 & n33648) | (n33538 & n33648);
  assign n27342 = n36593 | n27336;
  assign n27343 = n33649 | n27342;
  assign n27344 = ~n27339 & n27343;
  assign n27345 = x140 & x160;
  assign n27346 = x139 & x161;
  assign n27347 = n27345 & n27346;
  assign n27348 = n27345 | n27346;
  assign n27349 = ~n27347 & n27348;
  assign n27350 = n27344 & n27349;
  assign n27351 = n27344 | n27349;
  assign n27352 = ~n27350 & n27351;
  assign n33650 = n27107 | n27340;
  assign n33651 = n33538 | n33650;
  assign n37796 = ~n26932 & n27144;
  assign n37797 = (~n26931 & n27144) | (~n26931 & n37796) | (n27144 & n37796);
  assign n37586 = (n27144 & ~n27340) | (n27144 & n37797) | (~n27340 & n37797);
  assign n36617 = n27144 & ~n27340;
  assign n36618 = (~n33538 & n37586) | (~n33538 & n36617) | (n37586 & n36617);
  assign n27355 = n33651 & n36618;
  assign n33652 = n27153 | n27355;
  assign n33653 = (n27355 & n33543) | (n27355 & n33652) | (n33543 & n33652);
  assign n27357 = n27352 | n33653;
  assign n27358 = n27352 & n33653;
  assign n27359 = n27357 & ~n27358;
  assign n27360 = x138 & x162;
  assign n27361 = ~n27359 & n27360;
  assign n27362 = n27359 & ~n27360;
  assign n27363 = n27361 | n27362;
  assign n33654 = n27159 & n33565;
  assign n33655 = n27159 & n33504;
  assign n33656 = (n33407 & n33654) | (n33407 & n33655) | (n33654 & n33655);
  assign n33657 = n27158 & n27363;
  assign n33658 = (n27363 & n33656) | (n27363 & n33657) | (n33656 & n33657);
  assign n33659 = n27158 | n27363;
  assign n33660 = n33656 | n33659;
  assign n27368 = ~n33658 & n33660;
  assign n27369 = n27168 & n27368;
  assign n33580 = (n27100 & n27173) | (n27100 & n36569) | (n27173 & n36569);
  assign n33661 = n27167 & n27369;
  assign n33662 = (n27369 & n33580) | (n27369 & n33661) | (n33580 & n33661);
  assign n27372 = n27167 | n27368;
  assign n33663 = n27168 | n27372;
  assign n33664 = (n27372 & n33580) | (n27372 & n33663) | (n33580 & n33663);
  assign n27374 = ~n33662 & n33664;
  assign n27375 = x137 & x163;
  assign n27376 = n27374 & n27375;
  assign n27377 = n27374 | n27375;
  assign n27378 = ~n27376 & n27377;
  assign n27379 = x136 & x164;
  assign n27380 = n27378 & n27379;
  assign n27381 = n27378 | n27379;
  assign n27382 = ~n27380 & n27381;
  assign n27383 = n36591 | n27382;
  assign n27384 = n36591 & n27382;
  assign n27385 = n27383 & ~n27384;
  assign n27386 = n27190 & n27385;
  assign n27387 = n27303 & n27386;
  assign n27388 = n27189 | n27385;
  assign n27389 = n27192 | n27388;
  assign n27390 = ~n27387 & n27389;
  assign n27391 = x135 & x165;
  assign n27392 = n27390 & n27391;
  assign n27393 = n27390 | n27391;
  assign n27394 = ~n27392 & n27393;
  assign n27395 = x134 & x166;
  assign n27396 = n27394 & n27395;
  assign n27397 = n27394 | n27395;
  assign n27398 = ~n27396 & n27397;
  assign n27399 = n33394 | n33585;
  assign n37587 = n26858 | n26973;
  assign n37588 = n26972 | n37587;
  assign n36620 = n26973 | n33581;
  assign n36621 = (n33244 & n37588) | (n33244 & n36620) | (n37588 & n36620);
  assign n33666 = (n26973 & ~n27092) | (n26973 & n36621) | (~n27092 & n36621);
  assign n27401 = ~n27188 & n27195;
  assign n27402 = n27188 & ~n27195;
  assign n27403 = n27401 | n27402;
  assign n27404 = n27187 & ~n27403;
  assign n27405 = ~n27187 & n27403;
  assign n27406 = n27404 | n27405;
  assign n27407 = n33532 & ~n27406;
  assign n27408 = ~n33532 & n27406;
  assign n27409 = n27407 | n27408;
  assign n27410 = n33666 & n27409;
  assign n33667 = n27196 | n27410;
  assign n33668 = (n27196 & n27399) | (n27196 & n33667) | (n27399 & n33667);
  assign n27413 = n27398 | n33668;
  assign n27414 = n27398 & n33668;
  assign n27415 = n27413 & ~n27414;
  assign n37589 = n33585 & n33666;
  assign n37590 = n27409 & n37589;
  assign n37591 = n27086 & ~n37590;
  assign n37798 = n27086 & ~n33666;
  assign n37799 = (n27086 & ~n27409) | (n27086 & n37798) | (~n27409 & n37798);
  assign n37593 = (~n33394 & n37591) | (~n33394 & n37799) | (n37591 & n37799);
  assign n36625 = n27203 & n37593;
  assign n27418 = n27415 | n36625;
  assign n27419 = n33603 | n27418;
  assign n27420 = n26984 | n36625;
  assign n27421 = n27081 | n27420;
  assign n37594 = ~n27086 & n37590;
  assign n37800 = ~n27086 & n33666;
  assign n37801 = n27409 & n37800;
  assign n37596 = (n33394 & n37594) | (n33394 & n37801) | (n37594 & n37801);
  assign n36627 = (n27086 & n27203) | (n27086 & ~n37596) | (n27203 & ~n37596);
  assign n27423 = n27415 & n36627;
  assign n27424 = n27421 & n27423;
  assign n27425 = n27419 & ~n27424;
  assign n27426 = x133 & x167;
  assign n27427 = n27425 & n27426;
  assign n27428 = n27425 | n27426;
  assign n27429 = ~n27427 & n27428;
  assign n27430 = n33607 & n27429;
  assign n27431 = n33607 | n27429;
  assign n27432 = ~n27430 & n27431;
  assign n27433 = x132 & x168;
  assign n27434 = x131 & x169;
  assign n27435 = n27433 & n27434;
  assign n27436 = n27433 | n27434;
  assign n27437 = ~n27435 & n27436;
  assign n27438 = n27432 & n27437;
  assign n27439 = n27432 | n27437;
  assign n27440 = ~n27438 & n27439;
  assign n33669 = n27223 | n27225;
  assign n33670 = (n27076 & n27223) | (n27076 & n33669) | (n27223 & n33669);
  assign n27442 = n27440 & ~n33670;
  assign n33671 = n27075 | n27223;
  assign n33672 = n33520 | n33671;
  assign n27444 = n27224 & ~n27440;
  assign n27445 = n33672 & n27444;
  assign n27446 = n27442 | n27445;
  assign n27447 = x130 & x170;
  assign n27448 = ~n27446 & n27447;
  assign n27449 = n27446 & ~n27447;
  assign n27450 = n27448 | n27449;
  assign n27451 = ~n33601 & n27450;
  assign n27452 = n33601 & ~n27450;
  assign n27453 = n27451 | n27452;
  assign n27283 = n27069 | n27232;
  assign n27284 = n33518 | n27283;
  assign n33594 = n27071 & ~n27286;
  assign n33595 = (n27071 & ~n27288) | (n27071 & n33594) | (~n27288 & n33594);
  assign n27291 = n27284 & n33595;
  assign n33596 = n27238 | n27291;
  assign n36628 = n27453 & n33596;
  assign n36629 = n27291 & n27453;
  assign n36630 = (n27060 & n36628) | (n27060 & n36629) | (n36628 & n36629);
  assign n36631 = n27453 | n33596;
  assign n36632 = n27291 | n27453;
  assign n36633 = (n27060 & n36631) | (n27060 & n36632) | (n36631 & n36632);
  assign n27456 = ~n36630 & n36633;
  assign n27457 = x129 & x171;
  assign n27458 = n27456 & ~n27457;
  assign n27459 = ~n27456 & n27457;
  assign n27460 = n27458 | n27459;
  assign n27461 = n36587 & n27460;
  assign n27462 = n36587 | n27460;
  assign n27463 = ~n27461 & n27462;
  assign n27464 = n27281 & n27463;
  assign n27465 = n27281 | n27463;
  assign n27466 = ~n27464 & n27465;
  assign n27467 = n33593 & n27466;
  assign n27468 = n33593 | n27466;
  assign n27469 = ~n27467 & n27468;
  assign n27470 = n27279 & n27469;
  assign n27471 = n27279 | n27469;
  assign n27472 = ~n27470 & n27471;
  assign n27473 = n33591 & n27472;
  assign n27474 = n33591 | n27472;
  assign n27475 = ~n27473 & n27474;
  assign n27476 = n27277 & n27475;
  assign n27477 = n27277 | n27475;
  assign n27478 = ~n27476 & n27477;
  assign n27479 = n27276 & n27478;
  assign n27480 = n27276 | n27478;
  assign n27481 = ~n27479 & n27480;
  assign n27482 = n27275 & n27481;
  assign n27483 = n27275 | n27481;
  assign n27484 = ~n27482 & n27483;
  assign n27485 = n33589 & n27484;
  assign n27486 = n33589 | n27484;
  assign n27487 = ~n27485 & n27486;
  assign n27488 = n27482 | n27485;
  assign n27489 = x126 & x175;
  assign n33673 = n27476 | n27478;
  assign n33674 = (n27276 & n27476) | (n27276 & n33673) | (n27476 & n33673);
  assign n27491 = x127 & x174;
  assign n36634 = n27464 | n27466;
  assign n36635 = (n27464 & n33593) | (n27464 & n36634) | (n33593 & n36634);
  assign n27493 = n27059 | n27291;
  assign n27494 = n33506 | n27493;
  assign n27289 = n27286 & n27288;
  assign n27495 = n27284 & ~n27289;
  assign n27496 = n27071 | n27495;
  assign n27497 = n27453 & n27496;
  assign n27498 = n27494 & n27497;
  assign n33675 = n27457 & ~n27498;
  assign n33676 = n36633 & n33675;
  assign n33677 = n27460 | n33676;
  assign n33678 = (n36587 & n33676) | (n36587 & n33677) | (n33676 & n33677);
  assign n36636 = n27288 & n27446;
  assign n36637 = n27296 & n27446;
  assign n36638 = (n33600 & n36636) | (n33600 & n36637) | (n36636 & n36637);
  assign n33679 = n27446 & n27447;
  assign n33680 = (n27447 & n33601) | (n27447 & n33679) | (n33601 & n33679);
  assign n27505 = ~n36638 & n33680;
  assign n27506 = n27498 | n27505;
  assign n27507 = n27429 & ~n27433;
  assign n27508 = ~n27429 & n27433;
  assign n27509 = n27507 | n27508;
  assign n27510 = n33607 | n27509;
  assign n27511 = n33607 & n27509;
  assign n27512 = n27510 & ~n27511;
  assign n36639 = n27512 | n33669;
  assign n36640 = n27223 | n27512;
  assign n36641 = (n27076 & n36639) | (n27076 & n36640) | (n36639 & n36640);
  assign n27514 = n27224 & n27512;
  assign n27515 = n33672 & n27514;
  assign n33681 = n27434 & ~n27515;
  assign n33682 = n36641 & n33681;
  assign n33683 = n27446 | n33682;
  assign n33684 = (n33601 & n33682) | (n33601 & n33683) | (n33682 & n33683);
  assign n27519 = x131 & x170;
  assign n27520 = n27432 & n27433;
  assign n27521 = n27515 | n27520;
  assign n33685 = n27427 | n27429;
  assign n33686 = (n27427 & n33607) | (n27427 & n33685) | (n33607 & n33685);
  assign n27523 = x133 & x168;
  assign n27524 = n27394 & n33668;
  assign n36642 = (n27395 & n27396) | (n27395 & n33668) | (n27396 & n33668);
  assign n27527 = ~n27524 & n36642;
  assign n37597 = n27527 | n36627;
  assign n37598 = (n27415 & n27527) | (n27415 & n37597) | (n27527 & n37597);
  assign n36644 = (n27421 & n27527) | (n27421 & n37598) | (n27527 & n37598);
  assign n36645 = n27392 | n27394;
  assign n36646 = (n27392 & n33668) | (n27392 & n36645) | (n33668 & n36645);
  assign n33791 = n27179 | n27376;
  assign n36647 = (n27376 & n27378) | (n27376 & n33791) | (n27378 & n33791);
  assign n33690 = n27376 | n27378;
  assign n33691 = (n27184 & n36647) | (n27184 & n33690) | (n36647 & n33690);
  assign n27532 = x137 & x164;
  assign n27533 = x138 & x163;
  assign n27539 = n27344 & n27345;
  assign n27540 = n27344 | n27345;
  assign n27541 = ~n27539 & n27540;
  assign n27542 = n33653 & n27541;
  assign n33701 = n27346 & n27541;
  assign n33702 = (n27346 & n33653) | (n27346 & n33701) | (n33653 & n33701);
  assign n27545 = ~n27542 & n33702;
  assign n33692 = n27158 & n27359;
  assign n33703 = n27545 | n33692;
  assign n33704 = n27359 | n27545;
  assign n33705 = (n33656 & n33703) | (n33656 & n33704) | (n33703 & n33704);
  assign n27547 = x139 & x162;
  assign n33706 = n27539 | n33652;
  assign n36650 = n27345 | n27355;
  assign n36651 = (n27344 & n27355) | (n27344 & n36650) | (n27355 & n36650);
  assign n33708 = (n33543 & n33706) | (n33543 & n36651) | (n33706 & n36651);
  assign n27558 = x143 & x158;
  assign n33720 = n27558 & n36599;
  assign n36654 = n27316 & n27323;
  assign n37599 = (n27558 & n33720) | (n27558 & n36654) | (n33720 & n36654);
  assign n37600 = (n27323 & n27558) | (n27323 & n33720) | (n27558 & n33720);
  assign n37601 = (n33610 & n37599) | (n33610 & n37600) | (n37599 & n37600);
  assign n36656 = (n27130 & n27323) | (n27130 & n36654) | (n27323 & n36654);
  assign n36658 = (n27558 & n33720) | (n27558 & n36656) | (n33720 & n36656);
  assign n36659 = (n33483 & n37601) | (n33483 & n36658) | (n37601 & n36658);
  assign n33722 = n27558 | n36599;
  assign n37602 = n33722 | n36654;
  assign n37603 = n27323 | n33722;
  assign n37604 = (n33610 & n37602) | (n33610 & n37603) | (n37602 & n37603);
  assign n36661 = n33722 | n36656;
  assign n36662 = (n33483 & n37604) | (n33483 & n36661) | (n37604 & n36661);
  assign n27561 = ~n36659 & n36662;
  assign n36655 = (n27323 & n33610) | (n27323 & n36654) | (n33610 & n36654);
  assign n33716 = (n33483 & n36655) | (n33483 & n36656) | (n36655 & n36656);
  assign n36664 = n27316 | n27323;
  assign n37605 = n27318 & n36664;
  assign n37606 = (n27318 & n33610) | (n27318 & n37605) | (n33610 & n37605);
  assign n36666 = n27130 | n36664;
  assign n36668 = n27318 & n36666;
  assign n36669 = (n33483 & n37606) | (n33483 & n36668) | (n37606 & n36668);
  assign n27555 = ~n33716 & n36669;
  assign n33724 = n27555 & n27561;
  assign n33712 = n27311 & n27329;
  assign n36663 = (n27138 & n27329) | (n27138 & n33712) | (n27329 & n33712);
  assign n36670 = (n27561 & n33724) | (n27561 & n36663) | (n33724 & n36663);
  assign n36671 = (n27561 & n33712) | (n27561 & n33724) | (n33712 & n33724);
  assign n36672 = (n33546 & n36670) | (n33546 & n36671) | (n36670 & n36671);
  assign n33726 = n27555 | n27561;
  assign n36673 = n33726 | n36663;
  assign n36674 = n33712 | n33726;
  assign n36675 = (n33546 & n36673) | (n33546 & n36674) | (n36673 & n36674);
  assign n27564 = ~n36672 & n36675;
  assign n27565 = x142 & x159;
  assign n27566 = n27564 & n27565;
  assign n27567 = n27564 | n27565;
  assign n27568 = ~n27566 & n27567;
  assign n36652 = n27334 | n36615;
  assign n36653 = (n27334 & n27336) | (n27334 & n36652) | (n27336 & n36652);
  assign n36676 = n27568 & n36653;
  assign n36677 = n27334 & n27568;
  assign n36678 = (n33609 & n36676) | (n33609 & n36677) | (n36676 & n36677);
  assign n36679 = n27568 | n36653;
  assign n36680 = n27334 | n27568;
  assign n36681 = (n33609 & n36679) | (n33609 & n36680) | (n36679 & n36680);
  assign n27571 = ~n36678 & n36681;
  assign n33728 = n27540 & ~n27571;
  assign n33729 = n33708 & n33728;
  assign n33730 = ~n27540 & n27571;
  assign n33731 = (n27571 & ~n33708) | (n27571 & n33730) | (~n33708 & n33730);
  assign n27574 = n33729 | n33731;
  assign n27575 = x141 & x160;
  assign n27576 = x140 & x161;
  assign n27577 = n27575 & ~n27576;
  assign n27578 = ~n27575 & n27576;
  assign n27579 = n27577 | n27578;
  assign n27580 = n27574 & ~n27579;
  assign n27581 = ~n27574 & n27579;
  assign n27582 = n27580 | n27581;
  assign n27583 = n27547 & ~n27582;
  assign n27584 = ~n27547 & n27582;
  assign n27585 = n27583 | n27584;
  assign n27586 = n33705 | n27585;
  assign n27587 = n33705 & n27585;
  assign n27588 = n27586 & ~n27587;
  assign n33693 = (n27359 & n33656) | (n27359 & n33692) | (n33656 & n33692);
  assign n33694 = n27158 | n27359;
  assign n33696 = n27360 & n33694;
  assign n33697 = (n27360 & n33656) | (n27360 & n33696) | (n33656 & n33696);
  assign n27537 = ~n33693 & n33697;
  assign n33699 = n27369 | n27537;
  assign n36682 = n27588 & n33699;
  assign n36648 = n27167 | n27537;
  assign n36649 = (n27369 & n27537) | (n27369 & n36648) | (n27537 & n36648);
  assign n36683 = n27588 & n36649;
  assign n36684 = (n33580 & n36682) | (n33580 & n36683) | (n36682 & n36683);
  assign n36685 = n27588 | n33699;
  assign n36686 = n27588 | n36649;
  assign n36687 = (n33580 & n36685) | (n33580 & n36686) | (n36685 & n36686);
  assign n27591 = ~n36684 & n36687;
  assign n27592 = n27533 & n27591;
  assign n27593 = n27533 | n27591;
  assign n27594 = ~n27592 & n27593;
  assign n27595 = n27532 & n27594;
  assign n27596 = n27532 | n27594;
  assign n27597 = ~n27595 & n27596;
  assign n27598 = ~n33691 & n27597;
  assign n27599 = n33691 & ~n27597;
  assign n27600 = n27598 | n27599;
  assign n27601 = x136 & x165;
  assign n27602 = n27600 | n27601;
  assign n27603 = n27600 & n27601;
  assign n27604 = n27602 & ~n27603;
  assign n33732 = n27179 | n27378;
  assign n33733 = n27184 | n33732;
  assign n37607 = ~n27178 & n27379;
  assign n37608 = (~n27177 & n27379) | (~n27177 & n37607) | (n27379 & n37607);
  assign n36689 = (~n27378 & n27379) | (~n27378 & n37608) | (n27379 & n37608);
  assign n33735 = ~n27378 & n27379;
  assign n33736 = (~n27184 & n36689) | (~n27184 & n33735) | (n36689 & n33735);
  assign n27607 = n33733 & n33736;
  assign n33737 = n27386 | n27607;
  assign n33738 = (n27303 & n27607) | (n27303 & n33737) | (n27607 & n33737);
  assign n27609 = ~n27604 & n33738;
  assign n27610 = n27604 & ~n33738;
  assign n27611 = n27609 | n27610;
  assign n27612 = x135 & x166;
  assign n27613 = n27611 & n27612;
  assign n27614 = n27611 | n27612;
  assign n27615 = ~n27613 & n27614;
  assign n27616 = n36646 | n27615;
  assign n27617 = n36646 & n27615;
  assign n27618 = n27616 & ~n27617;
  assign n27619 = x134 & x167;
  assign n27620 = ~n27618 & n27619;
  assign n27621 = n27618 & ~n27619;
  assign n27622 = n27620 | n27621;
  assign n27623 = n36644 & n27622;
  assign n27624 = n36644 | n27622;
  assign n27625 = ~n27623 & n27624;
  assign n27626 = n27523 & n27625;
  assign n27627 = n27523 | n27625;
  assign n27628 = ~n27626 & n27627;
  assign n27629 = n33686 | n27628;
  assign n27630 = n33686 & n27628;
  assign n27631 = n27629 & ~n27630;
  assign n27632 = x132 & x169;
  assign n27633 = ~n27631 & n27632;
  assign n27634 = n27631 & ~n27632;
  assign n27635 = n27633 | n27634;
  assign n27636 = n27521 | n27635;
  assign n27637 = n27521 & n27635;
  assign n27638 = n27636 & ~n27637;
  assign n27639 = n27519 & n27638;
  assign n27640 = n27519 | n27638;
  assign n27641 = ~n27639 & n27640;
  assign n27642 = ~n33684 & n27641;
  assign n27643 = n33684 & ~n27641;
  assign n27644 = n27642 | n27643;
  assign n27645 = x130 & x171;
  assign n27646 = n27644 & n27645;
  assign n27647 = n27644 | n27645;
  assign n27648 = ~n27646 & n27647;
  assign n27649 = ~n27506 & n27648;
  assign n27650 = n27506 & ~n27648;
  assign n27651 = n27649 | n27650;
  assign n27652 = n33678 | n27651;
  assign n27653 = n33678 & n27651;
  assign n27654 = n27652 & ~n27653;
  assign n27655 = x129 & x172;
  assign n27656 = n27654 & ~n27655;
  assign n27657 = ~n27654 & n27655;
  assign n27658 = n27656 | n27657;
  assign n27659 = n36635 & n27658;
  assign n27660 = n36635 | n27658;
  assign n27661 = ~n27659 & n27660;
  assign n27662 = x128 & x173;
  assign n27663 = n27661 & n27662;
  assign n27664 = n27661 | n27662;
  assign n27665 = ~n27663 & n27664;
  assign n33739 = n27470 | n27472;
  assign n33740 = (n27470 & n33591) | (n27470 & n33739) | (n33591 & n33739);
  assign n27667 = n27665 & n33740;
  assign n27668 = n27665 | n33740;
  assign n27669 = ~n27667 & n27668;
  assign n27670 = n27491 & n27669;
  assign n27671 = n27491 | n27669;
  assign n27672 = ~n27670 & n27671;
  assign n27673 = n33674 & n27672;
  assign n27674 = n33674 | n27672;
  assign n27675 = ~n27673 & n27674;
  assign n27676 = n27489 & n27675;
  assign n27677 = n27489 | n27675;
  assign n27678 = ~n27676 & n27677;
  assign n27679 = n27488 & n27678;
  assign n27680 = n27488 | n27678;
  assign n27681 = ~n27679 & n27680;
  assign n33741 = n27676 | n27678;
  assign n33742 = (n27488 & n27676) | (n27488 & n33741) | (n27676 & n33741);
  assign n33743 = n27243 | n33676;
  assign n33744 = n27246 | n33743;
  assign n33745 = ~n27457 & n27498;
  assign n37802 = n27655 & ~n36633;
  assign n37803 = ~n27457 & n27655;
  assign n37804 = (n33745 & n37802) | (n33745 & n37803) | (n37802 & n37803);
  assign n37610 = (~n27651 & n27655) | (~n27651 & n37804) | (n27655 & n37804);
  assign n36691 = (n27655 & ~n33744) | (n27655 & n37610) | (~n33744 & n37610);
  assign n33748 = n27652 & n36691;
  assign n33749 = n27658 | n33748;
  assign n33750 = (n36635 & n33748) | (n36635 & n33749) | (n33748 & n33749);
  assign n33751 = n27505 | n27644;
  assign n33752 = n27498 | n33751;
  assign n33753 = n27505 & n27644;
  assign n33754 = (n27498 & n27644) | (n27498 & n33753) | (n27644 & n33753);
  assign n27692 = n27645 & ~n33754;
  assign n27693 = n33752 & n27692;
  assign n33746 = (n36633 & n27457) | (n36633 & ~n33745) | (n27457 & ~n33745);
  assign n27685 = n27651 & n33746;
  assign n33755 = n27685 | n27693;
  assign n33756 = (n27693 & n33744) | (n27693 & n33755) | (n33744 & n33755);
  assign n36692 = n27288 | n33682;
  assign n36693 = n27296 | n33682;
  assign n36694 = (n33600 & n36692) | (n33600 & n36693) | (n36692 & n36693);
  assign n33760 = ~n27434 & n27515;
  assign n33761 = (n27434 & n36641) | (n27434 & ~n33760) | (n36641 & ~n33760);
  assign n27698 = n27638 & n33761;
  assign n27699 = n36694 & n27698;
  assign n33757 = n27638 | n33683;
  assign n33758 = n27638 | n33682;
  assign n33759 = (n33601 & n33757) | (n33601 & n33758) | (n33757 & n33758);
  assign n33762 = n27519 & n33759;
  assign n33763 = ~n27699 & n33762;
  assign n27702 = n33754 | n33763;
  assign n33764 = n27520 & n27631;
  assign n33765 = (n27515 & n27631) | (n27515 & n33764) | (n27631 & n33764);
  assign n33766 = n27520 | n27631;
  assign n33768 = n27632 & n33766;
  assign n33769 = (n27515 & n27632) | (n27515 & n33768) | (n27632 & n33768);
  assign n27706 = ~n33765 & n33769;
  assign n36695 = n27706 | n33761;
  assign n36696 = (n27638 & n27706) | (n27638 & n36695) | (n27706 & n36695);
  assign n33771 = (n36694 & n27706) | (n36694 & n36696) | (n27706 & n36696);
  assign n27708 = n33686 | n27625;
  assign n27709 = n27301 | n27427;
  assign n27710 = n27220 | n27709;
  assign n27711 = n27428 & n27625;
  assign n37611 = n27523 & ~n27711;
  assign n37612 = (n27523 & ~n27710) | (n27523 & n37611) | (~n27710 & n37611);
  assign n36698 = n27708 & n37612;
  assign n33772 = n36698 | n33764;
  assign n33773 = n27631 | n36698;
  assign n33774 = (n27515 & n33772) | (n27515 & n33773) | (n33772 & n33773);
  assign n33775 = n27527 & n27618;
  assign n36699 = (n27423 & n27618) | (n27423 & n33775) | (n27618 & n33775);
  assign n36700 = n27618 & n33775;
  assign n36701 = (n27421 & n36699) | (n27421 & n36700) | (n36699 & n36700);
  assign n36702 = n27527 & n27619;
  assign n36703 = (n27618 & n27619) | (n27618 & n36702) | (n27619 & n36702);
  assign n36704 = (n27423 & n27619) | (n27423 & n36703) | (n27619 & n36703);
  assign n36705 = n27619 & n36703;
  assign n36706 = (n27421 & n36704) | (n27421 & n36705) | (n36704 & n36705);
  assign n27719 = ~n36701 & n36706;
  assign n33781 = n27711 | n27719;
  assign n33782 = (n27710 & n27719) | (n27710 & n33781) | (n27719 & n33781);
  assign n27721 = x135 & x167;
  assign n36707 = n27392 | n33667;
  assign n36708 = n27196 | n27392;
  assign n36709 = (n27399 & n36707) | (n27399 & n36708) | (n36707 & n36708);
  assign n27723 = n27393 & n27611;
  assign n27724 = n36709 & n27723;
  assign n33783 = n27392 | n27611;
  assign n36710 = n27394 | n33783;
  assign n36711 = (n33668 & n33783) | (n33668 & n36710) | (n33783 & n36710);
  assign n27726 = ~n27724 & n36711;
  assign n27727 = n27612 & n27726;
  assign n27729 = n27600 & n33738;
  assign n33788 = (n27601 & n27603) | (n27601 & n33738) | (n27603 & n33738);
  assign n27732 = ~n27729 & n33788;
  assign n33789 = n27723 | n27732;
  assign n33790 = (n36709 & n27732) | (n36709 & n33789) | (n27732 & n33789);
  assign n36712 = n27183 | n33791;
  assign n36713 = (n33536 & n33791) | (n33536 & n36712) | (n33791 & n36712);
  assign n33700 = (n33580 & n36649) | (n33580 & n33699) | (n36649 & n33699);
  assign n33795 = n27582 & n33703;
  assign n33796 = n27582 & n33704;
  assign n33797 = (n33656 & n33795) | (n33656 & n33796) | (n33795 & n33796);
  assign n27746 = n27571 & n27575;
  assign n27747 = n27571 | n27575;
  assign n27748 = ~n27746 & n27747;
  assign n36717 = n27540 | n27748;
  assign n36718 = (n27748 & n33708) | (n27748 & n36717) | (n33708 & n36717);
  assign n27549 = n27540 & n33708;
  assign n33803 = n27576 & ~n27748;
  assign n33804 = (~n27549 & n27576) | (~n27549 & n33803) | (n27576 & n33803);
  assign n27752 = n36718 & n33804;
  assign n33816 = n27540 | n27746;
  assign n33805 = n27566 | n27568;
  assign n36719 = (n27566 & n33805) | (n27566 & n36653) | (n33805 & n36653);
  assign n37613 = n27334 | n27566;
  assign n37614 = (n27566 & n27568) | (n27566 & n37613) | (n27568 & n37613);
  assign n36721 = (n33609 & n36719) | (n33609 & n37614) | (n36719 & n37614);
  assign n27756 = x143 & x159;
  assign n37806 = n27558 & n27756;
  assign n37893 = n36599 & n37806;
  assign n37807 = (n36656 & n37893) | (n36656 & n37806) | (n37893 & n37806);
  assign n37616 = n27756 & n37601;
  assign n37617 = (n33483 & n37807) | (n33483 & n37616) | (n37807 & n37616);
  assign n36723 = (n27756 & n33724) | (n27756 & n37617) | (n33724 & n37617);
  assign n36724 = (n27561 & n27756) | (n27561 & n37617) | (n27756 & n37617);
  assign n36725 = (n36663 & n36723) | (n36663 & n36724) | (n36723 & n36724);
  assign n36726 = (n33712 & n36723) | (n33712 & n36724) | (n36723 & n36724);
  assign n36727 = (n33546 & n36725) | (n33546 & n36726) | (n36725 & n36726);
  assign n37809 = n27558 | n27756;
  assign n37894 = (n27756 & n36599) | (n27756 & n37809) | (n36599 & n37809);
  assign n37810 = (n36656 & n37894) | (n36656 & n37809) | (n37894 & n37809);
  assign n37619 = n27756 | n37601;
  assign n37620 = (n33483 & n37810) | (n33483 & n37619) | (n37810 & n37619);
  assign n36729 = n33724 | n37620;
  assign n36730 = n27561 | n37620;
  assign n36731 = (n36663 & n36729) | (n36663 & n36730) | (n36729 & n36730);
  assign n36732 = (n33712 & n36729) | (n33712 & n36730) | (n36729 & n36730);
  assign n36733 = (n33546 & n36731) | (n33546 & n36732) | (n36731 & n36732);
  assign n27759 = ~n36727 & n36733;
  assign n27760 = x142 & x160;
  assign n27761 = n27759 & ~n27760;
  assign n27762 = ~n27759 & n27760;
  assign n27763 = n27761 | n27762;
  assign n27764 = x141 & x161;
  assign n27765 = ~n27763 & n27764;
  assign n27766 = n27763 & ~n27764;
  assign n27767 = n27765 | n27766;
  assign n27768 = n36721 | n27767;
  assign n27769 = n36721 & n27767;
  assign n27770 = n27768 & ~n27769;
  assign n33818 = n27747 & n27770;
  assign n36734 = n33816 & n33818;
  assign n36735 = n27746 & n33818;
  assign n36736 = (n33708 & n36734) | (n33708 & n36735) | (n36734 & n36735);
  assign n33820 = n27747 | n27770;
  assign n36737 = (n27770 & n33816) | (n27770 & n33820) | (n33816 & n33820);
  assign n36738 = (n27746 & n27770) | (n27746 & n33820) | (n27770 & n33820);
  assign n36739 = (n33708 & n36737) | (n33708 & n36738) | (n36737 & n36738);
  assign n27775 = ~n36736 & n36739;
  assign n27776 = x140 & x162;
  assign n27777 = n27775 | n27776;
  assign n27778 = n27775 & n27776;
  assign n27779 = n27777 & ~n27778;
  assign n33822 = n27752 | n27779;
  assign n33823 = n33797 | n33822;
  assign n33824 = n27752 & n27779;
  assign n33825 = (n27779 & n33797) | (n27779 & n33824) | (n33797 & n33824);
  assign n27782 = n33823 & ~n33825;
  assign n27783 = x139 & x163;
  assign n27784 = n27782 | n27783;
  assign n27785 = n27782 & n27783;
  assign n27786 = n27784 & ~n27785;
  assign n33798 = n27582 | n33703;
  assign n33799 = n27582 | n33704;
  assign n33800 = (n33656 & n33798) | (n33656 & n33799) | (n33798 & n33799);
  assign n27743 = n27547 & n33800;
  assign n27744 = ~n33797 & n27743;
  assign n33801 = n27588 | n27744;
  assign n33826 = n27786 | n33801;
  assign n33827 = n27744 | n27786;
  assign n33828 = (n33700 & n33826) | (n33700 & n33827) | (n33826 & n33827);
  assign n33829 = n27786 & n33801;
  assign n33830 = n27744 & n27786;
  assign n33831 = (n33700 & n33829) | (n33700 & n33830) | (n33829 & n33830);
  assign n27789 = n33828 & ~n33831;
  assign n27790 = x138 & x164;
  assign n27791 = ~n27789 & n27790;
  assign n27792 = n27789 & ~n27790;
  assign n27793 = n27791 | n27792;
  assign n36740 = n27377 | n27592;
  assign n36741 = (n27592 & n27594) | (n27592 & n36740) | (n27594 & n36740);
  assign n36742 = n27793 & ~n36741;
  assign n36743 = ~n27592 & n27793;
  assign n36744 = (~n36713 & n36742) | (~n36713 & n36743) | (n36742 & n36743);
  assign n36745 = ~n27793 & n36741;
  assign n36746 = n27592 & ~n27793;
  assign n36747 = (n36713 & n36745) | (n36713 & n36746) | (n36745 & n36746);
  assign n27797 = n36744 | n36747;
  assign n27798 = x137 & x165;
  assign n27799 = n27797 & n27798;
  assign n27800 = n27797 | n27798;
  assign n27801 = ~n27799 & n27800;
  assign n27735 = n27377 & n27594;
  assign n27736 = n36713 & n27735;
  assign n36714 = n27594 | n33690;
  assign n36715 = n27594 | n36647;
  assign n36716 = (n27184 & n36714) | (n27184 & n36715) | (n36714 & n36715);
  assign n27738 = ~n27736 & n36716;
  assign n27739 = n27532 & n27738;
  assign n33793 = n27600 | n27739;
  assign n36748 = n27801 | n33793;
  assign n36749 = n27739 | n27801;
  assign n36750 = (n33738 & n36748) | (n33738 & n36749) | (n36748 & n36749);
  assign n36751 = n27801 & n33793;
  assign n36752 = n27739 & n27801;
  assign n36753 = (n33738 & n36751) | (n33738 & n36752) | (n36751 & n36752);
  assign n27804 = n36750 & ~n36753;
  assign n27805 = x136 & x166;
  assign n27806 = ~n27804 & n27805;
  assign n27807 = n27804 & ~n27805;
  assign n27808 = n27806 | n27807;
  assign n27809 = n33790 | n27808;
  assign n27810 = n33790 & n27808;
  assign n27811 = n27809 & ~n27810;
  assign n37621 = n27727 | n27811;
  assign n37622 = n33775 | n37621;
  assign n33786 = n27618 | n27727;
  assign n36755 = n27811 | n33786;
  assign n36756 = (n27424 & n37622) | (n27424 & n36755) | (n37622 & n36755);
  assign n37623 = n27727 & n27811;
  assign n37624 = (n27811 & n33775) | (n27811 & n37623) | (n33775 & n37623);
  assign n36758 = n27811 & n33786;
  assign n36759 = (n27424 & n37624) | (n27424 & n36758) | (n37624 & n36758);
  assign n27814 = n36756 & ~n36759;
  assign n27815 = n27721 & n27814;
  assign n27816 = n27721 | n27814;
  assign n27817 = ~n27815 & n27816;
  assign n27818 = n33782 & n27817;
  assign n27819 = n33782 | n27817;
  assign n27820 = ~n27818 & n27819;
  assign n27821 = x134 & x168;
  assign n27822 = n27820 & n27821;
  assign n27823 = n27820 | n27821;
  assign n27824 = ~n27822 & n27823;
  assign n27825 = x133 & x169;
  assign n27826 = n27824 & n27825;
  assign n27827 = n27824 | n27825;
  assign n27828 = ~n27826 & n27827;
  assign n27829 = n33774 | n27828;
  assign n27830 = n33774 & n27828;
  assign n27831 = n27829 & ~n27830;
  assign n27832 = n33771 & n27831;
  assign n27833 = n33771 | n27831;
  assign n27834 = ~n27832 & n27833;
  assign n27835 = x132 & x170;
  assign n27836 = n27834 & n27835;
  assign n27837 = n27834 | n27835;
  assign n27838 = ~n27836 & n27837;
  assign n27839 = n27702 | n27838;
  assign n27840 = n27702 & n27838;
  assign n27841 = n27839 & ~n27840;
  assign n27842 = x131 & x171;
  assign n27843 = n27841 & ~n27842;
  assign n27844 = ~n27841 & n27842;
  assign n27845 = n27843 | n27844;
  assign n27846 = n33756 & n27845;
  assign n27847 = n33756 | n27845;
  assign n27848 = ~n27846 & n27847;
  assign n27849 = x130 & x172;
  assign n27850 = n27848 & n27849;
  assign n27851 = n27848 | n27849;
  assign n27852 = ~n27850 & n27851;
  assign n27853 = n33750 | n27852;
  assign n27854 = n33750 & n27852;
  assign n27855 = n27853 & ~n27854;
  assign n27856 = x129 & x173;
  assign n27857 = n27855 & ~n27856;
  assign n27858 = ~n27855 & n27856;
  assign n27859 = n27857 | n27858;
  assign n27860 = x128 & x174;
  assign n27861 = n27859 & n27860;
  assign n27862 = n27859 | n27860;
  assign n27863 = ~n27861 & n27862;
  assign n36760 = n27663 | n27665;
  assign n36761 = (n27663 & n33740) | (n27663 & n36760) | (n33740 & n36760);
  assign n27865 = n27863 | n36761;
  assign n27866 = n27863 & n36761;
  assign n27867 = n27865 & ~n27866;
  assign n33834 = n27670 | n27672;
  assign n33835 = (n27670 & n33674) | (n27670 & n33834) | (n33674 & n33834);
  assign n27869 = n27867 & n33835;
  assign n27870 = n27867 | n33835;
  assign n27871 = ~n27869 & n27870;
  assign n27872 = x127 & x175;
  assign n27873 = n27871 & n27872;
  assign n27874 = n27871 | n27872;
  assign n27875 = ~n27873 & n27874;
  assign n27876 = n33742 & n27875;
  assign n27877 = n33742 | n27875;
  assign n27878 = ~n27876 & n27877;
  assign n33836 = n27873 | n27875;
  assign n33837 = (n27873 & n33742) | (n27873 & n33836) | (n33742 & n33836);
  assign n27880 = n27859 | n36761;
  assign n33838 = ~n27859 & n27860;
  assign n33839 = (n27860 & ~n36761) | (n27860 & n33838) | (~n36761 & n33838);
  assign n27883 = n27880 & n33839;
  assign n33840 = n27867 | n27883;
  assign n33841 = (n27883 & n33835) | (n27883 & n33840) | (n33835 & n33840);
  assign n27885 = x129 & x174;
  assign n37811 = ~n27655 & n36633;
  assign n37812 = n27457 & ~n27655;
  assign n37813 = (~n33745 & n37811) | (~n33745 & n37812) | (n37811 & n37812);
  assign n37626 = n27651 & n37813;
  assign n36765 = n33744 & n37626;
  assign n33845 = (n27652 & n27655) | (n27652 & ~n36765) | (n27655 & ~n36765);
  assign n27888 = n27845 & ~n27849;
  assign n27889 = ~n27845 & n27849;
  assign n27890 = n27888 | n27889;
  assign n27891 = n33756 | n27890;
  assign n27892 = n33756 & n27890;
  assign n27893 = n27891 & ~n27892;
  assign n27894 = n33845 & n27893;
  assign n33842 = n27464 | n33748;
  assign n36762 = n27466 | n33842;
  assign n36763 = (n33593 & n33842) | (n33593 & n36762) | (n33842 & n36762);
  assign n36766 = n27856 & ~n36763;
  assign n36767 = (n27856 & ~n27894) | (n27856 & n36766) | (~n27894 & n36766);
  assign n33847 = n27853 & n36767;
  assign n33848 = n27859 | n33847;
  assign n33849 = (n36761 & n33847) | (n36761 & n33848) | (n33847 & n33848);
  assign n27895 = n36763 & n27894;
  assign n33850 = n27505 | n33763;
  assign n33851 = n27498 | n33850;
  assign n33852 = n27519 | n33759;
  assign n33853 = (n27519 & ~n27699) | (n27519 & n33852) | (~n27699 & n33852);
  assign n27902 = ~n27831 & n27835;
  assign n27903 = n27831 & ~n27835;
  assign n27904 = n27902 | n27903;
  assign n27905 = ~n33771 & n27904;
  assign n27906 = n33771 & ~n27904;
  assign n27907 = n27905 | n27906;
  assign n27908 = n33853 & n27907;
  assign n27909 = n33851 & n27908;
  assign n36768 = n27842 & ~n27909;
  assign n36769 = n27839 & n36768;
  assign n27912 = n27846 | n36769;
  assign n33854 = n27836 | n33851;
  assign n27914 = n36698 | n27824;
  assign n27915 = n33765 | n27914;
  assign n33856 = n27520 | n36698;
  assign n33857 = n27515 | n33856;
  assign n37627 = ~n27523 & n27711;
  assign n37628 = n27710 & n37627;
  assign n36771 = (n27523 & n27708) | (n27523 & ~n37628) | (n27708 & ~n37628);
  assign n27918 = n27824 & n36771;
  assign n27919 = n33857 & n27918;
  assign n27920 = n27915 & ~n27919;
  assign n27921 = n27825 & n27920;
  assign n33858 = n27831 | n27921;
  assign n33859 = (n27921 & n33771) | (n27921 & n33858) | (n33771 & n33858);
  assign n36772 = n27822 | n33856;
  assign n36773 = n27515 | n36772;
  assign n33861 = (n27822 & n27918) | (n27822 & n36773) | (n27918 & n36773);
  assign n27925 = n27612 | n27726;
  assign n27926 = n27811 & n27925;
  assign n33862 = n27527 | n27727;
  assign n33864 = n27926 & n33862;
  assign n36774 = n27721 & ~n33864;
  assign n36775 = n27721 & ~n27926;
  assign n36776 = (~n27424 & n36774) | (~n27424 & n36775) | (n36774 & n36775);
  assign n27929 = n36756 & n36776;
  assign n33866 = n27817 | n27929;
  assign n33867 = (n27929 & n33782) | (n27929 & n33866) | (n33782 & n33866);
  assign n33833 = (n27592 & n36713) | (n27592 & n36741) | (n36713 & n36741);
  assign n33710 = (n27334 & n33609) | (n27334 & n36653) | (n33609 & n36653);
  assign n33883 = n27763 | n33805;
  assign n33884 = n27566 | n27763;
  assign n33885 = (n33710 & n33883) | (n33710 & n33884) | (n33883 & n33884);
  assign n33886 = n27763 & n33805;
  assign n33887 = n27566 & n27763;
  assign n33888 = (n33710 & n33886) | (n33710 & n33887) | (n33886 & n33887);
  assign n27945 = n33885 & ~n33888;
  assign n33889 = n27747 & n27945;
  assign n36777 = n33816 & n33889;
  assign n36778 = n27746 & n33889;
  assign n36779 = (n33708 & n36777) | (n33708 & n36778) | (n36777 & n36778);
  assign n27947 = n27746 | n27945;
  assign n33891 = n27748 | n27947;
  assign n36780 = n27764 & n33891;
  assign n36781 = n27764 & n27947;
  assign n36782 = (n27549 & n36780) | (n27549 & n36781) | (n36780 & n36781);
  assign n27950 = ~n36779 & n36782;
  assign n33881 = n27752 & n27775;
  assign n33893 = n27950 | n33881;
  assign n33894 = n27775 | n27950;
  assign n33895 = (n33797 & n33893) | (n33797 & n33894) | (n33893 & n33894);
  assign n27952 = x141 & x162;
  assign n27953 = x142 & x161;
  assign n33817 = (n27746 & n33708) | (n27746 & n33816) | (n33708 & n33816);
  assign n27959 = x143 & x160;
  assign n33900 = n27566 & n27759;
  assign n36787 = (n27568 & n27759) | (n27568 & n33900) | (n27759 & n33900);
  assign n36788 = (n33900 & n36653) | (n33900 & n36787) | (n36653 & n36787);
  assign n36789 = (n27334 & n33900) | (n27334 & n36787) | (n33900 & n36787);
  assign n36790 = (n33609 & n36788) | (n33609 & n36789) | (n36788 & n36789);
  assign n33904 = n27959 & n36727;
  assign n33905 = (n27959 & n36790) | (n27959 & n33904) | (n36790 & n33904);
  assign n33906 = n27959 | n36727;
  assign n33907 = n36790 | n33906;
  assign n27963 = ~n33905 & n33907;
  assign n33897 = n27566 | n27759;
  assign n36783 = n27568 | n33897;
  assign n36784 = (n33897 & n36653) | (n33897 & n36783) | (n36653 & n36783);
  assign n36785 = (n27334 & n33897) | (n27334 & n36783) | (n33897 & n36783);
  assign n36786 = (n33609 & n36784) | (n33609 & n36785) | (n36784 & n36785);
  assign n27956 = n27760 & ~n36790;
  assign n27957 = n36786 & n27956;
  assign n36792 = n27957 & n27963;
  assign n37629 = (n27963 & n33889) | (n27963 & n36792) | (n33889 & n36792);
  assign n36793 = (n33817 & n37629) | (n33817 & n36792) | (n37629 & n36792);
  assign n36795 = n27957 | n27963;
  assign n37630 = n33889 | n36795;
  assign n36796 = (n33817 & n37630) | (n33817 & n36795) | (n37630 & n36795);
  assign n27966 = ~n36793 & n36796;
  assign n27967 = n27953 & n27966;
  assign n27968 = n27953 | n27966;
  assign n27969 = ~n27967 & n27968;
  assign n27970 = n27952 & ~n27969;
  assign n27971 = ~n27952 & n27969;
  assign n27972 = n27970 | n27971;
  assign n27973 = n33895 | n27972;
  assign n27974 = n33895 & n27972;
  assign n27975 = n27973 & ~n27974;
  assign n33882 = (n27775 & n33797) | (n27775 & n33881) | (n33797 & n33881);
  assign n33908 = n27752 | n27775;
  assign n33909 = n33797 | n33908;
  assign n27977 = ~n33882 & n33909;
  assign n27980 = n27776 | n27977;
  assign n27978 = n27776 & n27977;
  assign n33911 = n27744 | n27978;
  assign n33913 = n27980 & n33911;
  assign n33910 = n27978 | n33801;
  assign n33914 = n27980 & n33910;
  assign n33915 = (n33700 & n33913) | (n33700 & n33914) | (n33913 & n33914);
  assign n27982 = n27975 & n33915;
  assign n33870 = n27782 & n33801;
  assign n33916 = n27978 | n33870;
  assign n33871 = n27744 & n27782;
  assign n33917 = n27978 | n33871;
  assign n33918 = (n33700 & n33916) | (n33700 & n33917) | (n33916 & n33917);
  assign n27984 = n27975 | n33918;
  assign n27985 = ~n27982 & n27984;
  assign n27986 = x140 & x163;
  assign n27987 = n27985 & n27986;
  assign n27988 = n27985 | n27986;
  assign n27989 = ~n27987 & n27988;
  assign n33872 = (n33700 & n33870) | (n33700 & n33871) | (n33870 & n33871);
  assign n36797 = (n27783 & n27785) | (n27783 & n33801) | (n27785 & n33801);
  assign n33874 = n27744 | n27782;
  assign n33877 = n27783 & n33874;
  assign n33878 = (n33700 & n36797) | (n33700 & n33877) | (n36797 & n33877);
  assign n27940 = ~n33872 & n33878;
  assign n33879 = n27789 | n27940;
  assign n33919 = n27989 | n33879;
  assign n33920 = n27940 | n27989;
  assign n33921 = (n33833 & n33919) | (n33833 & n33920) | (n33919 & n33920);
  assign n33922 = n27989 & n33879;
  assign n33923 = n27940 & n27989;
  assign n33924 = (n33833 & n33922) | (n33833 & n33923) | (n33922 & n33923);
  assign n27992 = n33921 & ~n33924;
  assign n27993 = x139 & x164;
  assign n27994 = x138 & x165;
  assign n27995 = n27993 & n27994;
  assign n27996 = n27993 | n27994;
  assign n27997 = ~n27995 & n27996;
  assign n27998 = n27992 & n27997;
  assign n27999 = n27992 | n27997;
  assign n28000 = ~n27998 & n27999;
  assign n28002 = n27532 | n27738;
  assign n28003 = n27797 & n28002;
  assign n33925 = n27739 & n28003;
  assign n33926 = (n28003 & n33738) | (n28003 & n33925) | (n33738 & n33925);
  assign n36798 = n27789 | n36741;
  assign n36799 = n27592 | n27789;
  assign n36800 = (n36713 & n36798) | (n36713 & n36799) | (n36798 & n36799);
  assign n36801 = (n27790 & n27791) | (n27790 & ~n36741) | (n27791 & ~n36741);
  assign n36802 = (~n27592 & n27790) | (~n27592 & n27791) | (n27790 & n27791);
  assign n36803 = (~n36713 & n36801) | (~n36713 & n36802) | (n36801 & n36802);
  assign n28007 = n36800 & n36803;
  assign n33928 = ~n28000 & n28007;
  assign n33929 = (~n28000 & n33926) | (~n28000 & n33928) | (n33926 & n33928);
  assign n33930 = n28000 & ~n28007;
  assign n33931 = ~n33926 & n33930;
  assign n28011 = n33929 | n33931;
  assign n33932 = n27797 | n33793;
  assign n33933 = n27739 | n27797;
  assign n33934 = (n33738 & n33932) | (n33738 & n33933) | (n33932 & n33933);
  assign n28013 = ~n33926 & n33934;
  assign n28014 = n27798 & n28013;
  assign n28015 = n28011 | n28014;
  assign n33935 = n27804 | n28015;
  assign n33936 = (n28015 & n33790) | (n28015 & n33935) | (n33790 & n33935);
  assign n28018 = n27798 | n28013;
  assign n28019 = n28011 & n28018;
  assign n33937 = n28014 & n28019;
  assign n33938 = (n28019 & n33790) | (n28019 & n33937) | (n33790 & n33937);
  assign n28021 = n33936 & ~n33938;
  assign n28022 = x137 & x166;
  assign n28023 = n28021 & n28022;
  assign n28024 = n28021 | n28022;
  assign n28025 = ~n28023 & n28024;
  assign n33865 = (n27424 & n27926) | (n27424 & n33864) | (n27926 & n33864);
  assign n27931 = n33790 & n27804;
  assign n33868 = n27804 & n27805;
  assign n33869 = (n27805 & n33790) | (n27805 & n33868) | (n33790 & n33868);
  assign n27934 = ~n27931 & n33869;
  assign n33939 = n27934 & n28025;
  assign n33940 = (n28025 & n33865) | (n28025 & n33939) | (n33865 & n33939);
  assign n33941 = n27934 | n28025;
  assign n33942 = n33865 | n33941;
  assign n28028 = ~n33940 & n33942;
  assign n28029 = x136 & x167;
  assign n28030 = n28028 & n28029;
  assign n28031 = n28028 | n28029;
  assign n28032 = ~n28030 & n28031;
  assign n28033 = x135 & x168;
  assign n28034 = n28032 & n28033;
  assign n28035 = n28032 | n28033;
  assign n28036 = ~n28034 & n28035;
  assign n28037 = n33867 | n28036;
  assign n28038 = n33867 & n28036;
  assign n28039 = n28037 & ~n28038;
  assign n28040 = x134 & x169;
  assign n28041 = n28039 | n28040;
  assign n28042 = n28039 & n28040;
  assign n28043 = n28041 & ~n28042;
  assign n28044 = ~n33861 & n28043;
  assign n28045 = n33861 & ~n28043;
  assign n28046 = n28044 | n28045;
  assign n28047 = x133 & x170;
  assign n28048 = n28046 & n28047;
  assign n28049 = n28046 | n28047;
  assign n28050 = ~n28048 & n28049;
  assign n28051 = n33859 | n28050;
  assign n28052 = n33859 & n28050;
  assign n28053 = n28051 & ~n28052;
  assign n36804 = n27908 & n28053;
  assign n36805 = n27836 & n28053;
  assign n36806 = (n33854 & n36804) | (n33854 & n36805) | (n36804 & n36805);
  assign n36807 = n27908 | n28053;
  assign n36808 = n27836 | n28053;
  assign n36809 = (n33854 & n36807) | (n33854 & n36808) | (n36807 & n36808);
  assign n28056 = ~n36806 & n36809;
  assign n28057 = x132 & x171;
  assign n28058 = n28056 & n28057;
  assign n28059 = n28056 | n28057;
  assign n28060 = ~n28058 & n28059;
  assign n28061 = x131 & x172;
  assign n28062 = n28060 & n28061;
  assign n28063 = n28060 | n28061;
  assign n28064 = ~n28062 & n28063;
  assign n28065 = n27912 | n28064;
  assign n28066 = n27912 & n28064;
  assign n28067 = n28065 & ~n28066;
  assign n33943 = n27850 & n28067;
  assign n33944 = (n27895 & n28067) | (n27895 & n33943) | (n28067 & n33943);
  assign n33945 = n27850 | n28067;
  assign n33946 = n27895 | n33945;
  assign n28070 = ~n33944 & n33946;
  assign n28071 = x130 & x173;
  assign n28072 = n28070 & n28071;
  assign n28073 = n28070 | n28071;
  assign n28074 = ~n28072 & n28073;
  assign n28075 = n33849 | n28074;
  assign n28076 = n33849 & n28074;
  assign n28077 = n28075 & ~n28076;
  assign n28078 = n27885 & n28077;
  assign n28079 = n27885 | n28077;
  assign n28080 = ~n28078 & n28079;
  assign n28081 = ~n33841 & n28080;
  assign n28082 = n33841 & ~n28080;
  assign n28083 = n28081 | n28082;
  assign n28084 = x128 & x175;
  assign n28085 = n28083 & n28084;
  assign n28086 = n28083 | n28084;
  assign n28087 = ~n28085 & n28086;
  assign n28088 = n33837 & n28087;
  assign n28089 = n33837 | n28087;
  assign n28090 = ~n28088 & n28089;
  assign n28091 = n33841 & n28080;
  assign n28092 = n27663 | n33847;
  assign n36810 = n27665 | n28092;
  assign n36811 = (n28092 & n33740) | (n28092 & n36810) | (n33740 & n36810);
  assign n36812 = ~n27856 & n36763;
  assign n36813 = n27894 & n36812;
  assign n33948 = (n27853 & n27856) | (n27853 & ~n36813) | (n27856 & ~n36813);
  assign n36814 = n27850 | n36763;
  assign n36815 = (n27850 & n27894) | (n27850 & n36814) | (n27894 & n36814);
  assign n28095 = ~n28067 & n28071;
  assign n28096 = n28067 & ~n28071;
  assign n28097 = n28095 | n28096;
  assign n28098 = ~n36815 & n28097;
  assign n28099 = n36815 & ~n28097;
  assign n28100 = n28098 | n28099;
  assign n28101 = n33948 & n28100;
  assign n33951 = n28072 | n28101;
  assign n33952 = (n28072 & n36811) | (n28072 & n33951) | (n36811 & n33951);
  assign n28107 = n33756 | n36769;
  assign n36816 = ~n27842 & n27909;
  assign n36817 = (n27839 & n27842) | (n27839 & ~n36816) | (n27842 & ~n36816);
  assign n28109 = n28060 & n36817;
  assign n28110 = n28107 & n28109;
  assign n28111 = n36769 | n28060;
  assign n28112 = n27846 | n28111;
  assign n28113 = ~n28110 & n28112;
  assign n28114 = n28061 & n28113;
  assign n36818 = n28058 | n36769;
  assign n36819 = n33756 | n36818;
  assign n33954 = (n28058 & n28109) | (n28058 & n36819) | (n28109 & n36819);
  assign n33955 = n27706 | n27825;
  assign n33956 = (n27706 & n27920) | (n27706 & n33955) | (n27920 & n33955);
  assign n28117 = n27699 | n33956;
  assign n28121 = n33861 & n28039;
  assign n33957 = (n28040 & n28042) | (n28040 & n33861) | (n28042 & n33861);
  assign n28124 = ~n28121 & n33957;
  assign n28118 = n27825 | n27920;
  assign n28119 = n28046 & n28118;
  assign n33958 = n28119 | n28124;
  assign n33959 = (n28117 & n28124) | (n28117 & n33958) | (n28124 & n33958);
  assign n28126 = n27719 | n27929;
  assign n33960 = n27711 | n28126;
  assign n33961 = (n27710 & n28126) | (n27710 & n33960) | (n28126 & n33960);
  assign n36820 = ~n27721 & n33864;
  assign n36821 = ~n27721 & n27926;
  assign n36822 = (n27424 & n36820) | (n27424 & n36821) | (n36820 & n36821);
  assign n33963 = (n27721 & n36756) | (n27721 & ~n36822) | (n36756 & ~n36822);
  assign n28130 = n28022 & n28029;
  assign n28131 = n28022 | n28029;
  assign n28132 = ~n28130 & n28131;
  assign n28133 = n28021 & ~n28132;
  assign n28134 = ~n28021 & n28132;
  assign n28135 = n28133 | n28134;
  assign n33964 = ~n27934 & n28135;
  assign n33965 = ~n33865 & n33964;
  assign n33966 = n27934 & ~n28135;
  assign n33967 = (~n28135 & n33865) | (~n28135 & n33966) | (n33865 & n33966);
  assign n28138 = n33965 | n33967;
  assign n28139 = n33963 & n28138;
  assign n33968 = n28030 | n28139;
  assign n33969 = (n28030 & n33961) | (n28030 & n33968) | (n33961 & n33968);
  assign n33970 = n27934 | n28023;
  assign n36823 = n33864 | n33970;
  assign n36824 = n27926 | n33970;
  assign n36825 = (n27424 & n36823) | (n27424 & n36824) | (n36823 & n36824);
  assign n36826 = (n27940 & n33879) | (n27940 & n36741) | (n33879 & n36741);
  assign n36827 = (n27592 & n27940) | (n27592 & n33879) | (n27940 & n33879);
  assign n36828 = (n36713 & n36826) | (n36713 & n36827) | (n36826 & n36827);
  assign n28143 = n27989 & n27993;
  assign n28144 = n27989 | n27993;
  assign n28145 = ~n28143 & n28144;
  assign n28146 = n36828 | n28145;
  assign n28147 = n36828 & n28145;
  assign n28148 = n28146 & ~n28147;
  assign n33972 = n28007 & n28148;
  assign n33973 = (n28148 & n33926) | (n28148 & n33972) | (n33926 & n33972);
  assign n36829 = n27994 & n28007;
  assign n36830 = (n27994 & n28148) | (n27994 & n36829) | (n28148 & n36829);
  assign n33977 = (n27994 & n33926) | (n27994 & n36830) | (n33926 & n36830);
  assign n28152 = ~n33973 & n33977;
  assign n28153 = n33938 | n28152;
  assign n28154 = n27992 & n27993;
  assign n33978 = n28154 | n33972;
  assign n33979 = n28148 | n28154;
  assign n33980 = (n33926 & n33978) | (n33926 & n33979) | (n33978 & n33979);
  assign n28159 = x142 & x162;
  assign n33902 = n27957 | n33889;
  assign n28161 = x143 & x161;
  assign n36833 = n27959 & n28161;
  assign n37631 = n36727 & n36833;
  assign n36834 = (n36790 & n37631) | (n36790 & n36833) | (n37631 & n36833);
  assign n36831 = (n27963 & n28161) | (n27963 & n36834) | (n28161 & n36834);
  assign n36835 = (n33902 & n36831) | (n33902 & n36834) | (n36831 & n36834);
  assign n36836 = (n27957 & n36831) | (n27957 & n36834) | (n36831 & n36834);
  assign n36837 = (n33817 & n36835) | (n33817 & n36836) | (n36835 & n36836);
  assign n36840 = n27959 | n28161;
  assign n37632 = (n28161 & n36727) | (n28161 & n36840) | (n36727 & n36840);
  assign n36841 = (n36790 & n37632) | (n36790 & n36840) | (n37632 & n36840);
  assign n36838 = n27963 | n36841;
  assign n36842 = (n33902 & n36838) | (n33902 & n36841) | (n36838 & n36841);
  assign n36843 = (n27957 & n36838) | (n27957 & n36841) | (n36838 & n36841);
  assign n36844 = (n33817 & n36842) | (n33817 & n36843) | (n36842 & n36843);
  assign n28164 = ~n36837 & n36844;
  assign n28165 = n28159 & n28164;
  assign n28166 = n28159 | n28164;
  assign n28167 = ~n28165 & n28166;
  assign n33984 = n27967 | n27969;
  assign n36845 = n28167 | n33984;
  assign n36846 = n27967 | n28167;
  assign n36847 = (n33895 & n36845) | (n33895 & n36846) | (n36845 & n36846);
  assign n36848 = n28167 & n33984;
  assign n36849 = n27967 & n28167;
  assign n36850 = (n33895 & n36848) | (n33895 & n36849) | (n36848 & n36849);
  assign n28170 = n36847 & ~n36850;
  assign n28171 = x141 & x163;
  assign n28172 = ~n28170 & n28171;
  assign n28173 = n28170 & ~n28171;
  assign n28174 = n28172 | n28173;
  assign n36851 = n27969 | n33893;
  assign n36852 = n27969 | n33894;
  assign n36853 = (n33797 & n36851) | (n33797 & n36852) | (n36851 & n36852);
  assign n33994 = (n27952 & n27970) | (n27952 & ~n33895) | (n27970 & ~n33895);
  assign n28177 = n36853 & n33994;
  assign n33995 = n27975 | n28177;
  assign n36854 = n28174 & n33995;
  assign n36855 = n28174 & n28177;
  assign n36856 = (n33915 & n36854) | (n33915 & n36855) | (n36854 & n36855);
  assign n36857 = n28174 | n33995;
  assign n36858 = n28174 | n28177;
  assign n36859 = (n33915 & n36857) | (n33915 & n36858) | (n36857 & n36858);
  assign n28181 = ~n36856 & n36859;
  assign n28184 = n27987 | n28181;
  assign n34000 = n28184 | n33923;
  assign n34001 = n28184 | n33922;
  assign n34002 = (n33833 & n34000) | (n33833 & n34001) | (n34000 & n34001);
  assign n28187 = x140 & x164;
  assign n28188 = x139 & x165;
  assign n28189 = n28187 & n28188;
  assign n28190 = n28187 | n28188;
  assign n28191 = ~n28189 & n28190;
  assign n28182 = n27988 & n28181;
  assign n36860 = n27940 | n27986;
  assign n36861 = (n27940 & n27985) | (n27940 & n36860) | (n27985 & n36860);
  assign n33997 = n28182 & n36861;
  assign n33981 = n27987 | n33879;
  assign n33998 = n28182 & n33981;
  assign n33999 = (n33833 & n33997) | (n33833 & n33998) | (n33997 & n33998);
  assign n36862 = n28191 & ~n33999;
  assign n36863 = n34002 & n36862;
  assign n36864 = ~n28191 & n33999;
  assign n36865 = (n28191 & n34002) | (n28191 & ~n36864) | (n34002 & ~n36864);
  assign n28194 = ~n36863 & n36865;
  assign n28195 = n33980 | n28194;
  assign n28196 = n33980 & n28194;
  assign n28197 = n28195 & ~n28196;
  assign n28198 = x138 & x166;
  assign n28199 = ~n28197 & n28198;
  assign n28200 = n28197 & ~n28198;
  assign n28201 = n28199 | n28200;
  assign n28202 = n28153 | n28201;
  assign n28203 = n28153 & n28201;
  assign n28204 = n28202 & ~n28203;
  assign n28205 = n28024 & n28204;
  assign n28206 = n36825 & n28205;
  assign n28207 = n28023 | n28204;
  assign n36866 = n28207 | n33939;
  assign n36867 = n28025 | n28207;
  assign n36868 = (n33865 & n36866) | (n33865 & n36867) | (n36866 & n36867);
  assign n28209 = ~n28206 & n36868;
  assign n28210 = x137 & x167;
  assign n28211 = n28209 & n28210;
  assign n28212 = n28209 | n28210;
  assign n28213 = ~n28211 & n28212;
  assign n28214 = n33969 & n28213;
  assign n28215 = n33969 | n28213;
  assign n28216 = ~n28214 & n28215;
  assign n28217 = x136 & x168;
  assign n28218 = n28216 & n28217;
  assign n28219 = n28216 | n28217;
  assign n28220 = ~n28218 & n28219;
  assign n28221 = n33867 | n28032;
  assign n37633 = n28033 & ~n33963;
  assign n37634 = (n28033 & ~n28138) | (n28033 & n37633) | (~n28138 & n37633);
  assign n36870 = (n28033 & ~n33961) | (n28033 & n37634) | (~n33961 & n37634);
  assign n34004 = n28221 & n36870;
  assign n28224 = n28220 | n34004;
  assign n28225 = n28121 | n28224;
  assign n28232 = x135 & x169;
  assign n28226 = n27822 | n34004;
  assign n34005 = n28226 | n33857;
  assign n34006 = (n27918 & n28226) | (n27918 & n34005) | (n28226 & n34005);
  assign n37635 = ~n28033 & n33963;
  assign n37636 = n28138 & n37635;
  assign n37895 = n28232 & n37636;
  assign n37896 = n33961 & n37895;
  assign n37815 = ~n28033 & n28232;
  assign n37816 = (~n28221 & n37896) | (~n28221 & n37815) | (n37896 & n37815);
  assign n37638 = (~n28220 & n28232) | (~n28220 & n37816) | (n28232 & n37816);
  assign n36874 = (n28232 & ~n34006) | (n28232 & n37638) | (~n34006 & n37638);
  assign n34010 = n28225 & n36874;
  assign n37897 = n28232 | n37636;
  assign n37898 = (n28232 & n33961) | (n28232 & n37897) | (n33961 & n37897);
  assign n37818 = n28033 & ~n28232;
  assign n37819 = (n28221 & ~n37898) | (n28221 & n37818) | (~n37898 & n37818);
  assign n37640 = n28220 & n37819;
  assign n36876 = n34006 & n37640;
  assign n34012 = (n28225 & n28232) | (n28225 & ~n36876) | (n28232 & ~n36876);
  assign n28235 = ~n34010 & n34012;
  assign n28236 = n33959 & n28235;
  assign n28237 = n33959 | n28235;
  assign n28238 = ~n28236 & n28237;
  assign n28239 = x134 & x170;
  assign n28240 = n28238 & n28239;
  assign n28241 = n28238 | n28239;
  assign n28242 = ~n28240 & n28241;
  assign n28243 = x133 & x171;
  assign n28244 = n28242 & n28243;
  assign n28245 = n28242 | n28243;
  assign n28246 = ~n28244 & n28245;
  assign n28247 = n27921 | n28046;
  assign n28248 = n27832 | n28247;
  assign n34013 = n28047 & ~n28119;
  assign n34014 = (n28047 & ~n28117) | (n28047 & n34013) | (~n28117 & n34013);
  assign n28250 = n28248 & n34014;
  assign n34015 = n28053 | n28250;
  assign n36877 = (n27908 & n28250) | (n27908 & n34015) | (n28250 & n34015);
  assign n36878 = (n27836 & n28250) | (n27836 & n34015) | (n28250 & n34015);
  assign n36879 = (n33854 & n36877) | (n33854 & n36878) | (n36877 & n36878);
  assign n28252 = n28246 | n36879;
  assign n28253 = n28246 & n36879;
  assign n28254 = n28252 & ~n28253;
  assign n28255 = x132 & x172;
  assign n28256 = ~n28254 & n28255;
  assign n28257 = n28254 & ~n28255;
  assign n28258 = n28256 | n28257;
  assign n28259 = n33954 | n28258;
  assign n28260 = n33954 & n28258;
  assign n28261 = n28259 & ~n28260;
  assign n28262 = n28114 | n28261;
  assign n28263 = n33944 | n28262;
  assign n28270 = x131 & x173;
  assign n36880 = n27849 | n28061;
  assign n36881 = (n27848 & n28061) | (n27848 & n36880) | (n28061 & n36880);
  assign n34018 = (n27850 & n28113) | (n27850 & n36881) | (n28113 & n36881);
  assign n36882 = n34018 | n36763;
  assign n36883 = (n27894 & n34018) | (n27894 & n36882) | (n34018 & n36882);
  assign n28266 = n28061 | n28113;
  assign n28267 = n28261 & n28266;
  assign n28268 = n36883 & n28267;
  assign n36884 = n28268 & ~n28270;
  assign n36885 = (n28263 & n28270) | (n28263 & ~n36884) | (n28270 & ~n36884);
  assign n36886 = ~n28268 & n28270;
  assign n36887 = n28263 & n36886;
  assign n28273 = n36885 & ~n36887;
  assign n28274 = n33952 & n28273;
  assign n28275 = n33952 | n28273;
  assign n28276 = ~n28274 & n28275;
  assign n28277 = x130 & x174;
  assign n28278 = n28276 & n28277;
  assign n28279 = n28276 | n28277;
  assign n28280 = ~n28278 & n28279;
  assign n36888 = n27885 & ~n33948;
  assign n36889 = (n27885 & ~n28100) | (n27885 & n36888) | (~n28100 & n36888);
  assign n33950 = (n27885 & ~n36811) | (n27885 & n36889) | (~n36811 & n36889);
  assign n28104 = n28075 & n33950;
  assign n34019 = n28104 & n28280;
  assign n34020 = (n28091 & n28280) | (n28091 & n34019) | (n28280 & n34019);
  assign n34021 = n28104 | n28280;
  assign n34022 = n28091 | n34021;
  assign n28283 = ~n34020 & n34022;
  assign n28284 = x129 & x175;
  assign n28285 = n28283 | n28284;
  assign n28286 = n28283 & n28284;
  assign n28287 = n28285 & ~n28286;
  assign n34023 = n28085 | n28087;
  assign n34024 = (n28085 & n33837) | (n28085 & n34023) | (n33837 & n34023);
  assign n28289 = n28287 & ~n34024;
  assign n28290 = ~n28287 & n34024;
  assign n28291 = n28289 | n28290;
  assign n28294 = n33954 & n28254;
  assign n34027 = n28254 & n28255;
  assign n34028 = (n28255 & n33954) | (n28255 & n34027) | (n33954 & n34027);
  assign n28297 = ~n28294 & n34028;
  assign n28298 = n28268 | n28297;
  assign n28299 = n28242 | n36879;
  assign n28300 = n27836 | n28250;
  assign n28301 = n27909 | n28300;
  assign n28120 = n28117 & n28119;
  assign n28302 = ~n28120 & n28248;
  assign n28303 = n28047 | n28302;
  assign n28304 = n28232 & n28239;
  assign n28305 = n28232 | n28239;
  assign n28306 = ~n28304 & n28305;
  assign n37899 = ~n28306 & n37636;
  assign n37900 = n33961 & n37899;
  assign n37821 = n28033 | n28306;
  assign n37822 = (n28221 & ~n37900) | (n28221 & n37821) | (~n37900 & n37821);
  assign n37642 = (n28220 & n28306) | (n28220 & n37822) | (n28306 & n37822);
  assign n36891 = (n28306 & n34006) | (n28306 & n37642) | (n34006 & n37642);
  assign n34030 = n28225 & ~n36891;
  assign n37901 = n28306 & ~n37636;
  assign n37902 = (n28306 & ~n33961) | (n28306 & n37901) | (~n33961 & n37901);
  assign n37824 = n28033 & n28306;
  assign n37825 = (n28221 & n37902) | (n28221 & n37824) | (n37902 & n37824);
  assign n37644 = n28220 & n37825;
  assign n36893 = n34006 & n37644;
  assign n34032 = (~n28225 & n28306) | (~n28225 & n36893) | (n28306 & n36893);
  assign n28309 = n34030 | n34032;
  assign n28310 = ~n33959 & n28309;
  assign n28311 = n33959 & ~n28309;
  assign n28312 = n28310 | n28311;
  assign n28313 = n28303 & n28312;
  assign n28314 = n28301 & n28313;
  assign n28315 = n28299 & ~n28314;
  assign n28316 = n28243 & n28315;
  assign n34033 = n28254 | n28316;
  assign n34034 = (n28316 & n33954) | (n28316 & n34033) | (n33954 & n34033);
  assign n34035 = n28240 | n28313;
  assign n34036 = (n28240 & n28301) | (n28240 & n34035) | (n28301 & n34035);
  assign n34037 = n28235 | n34010;
  assign n34038 = (n33959 & n34010) | (n33959 & n34037) | (n34010 & n34037);
  assign n28320 = x137 & x168;
  assign n34039 = n28152 & n28197;
  assign n34040 = (n28197 & n33938) | (n28197 & n34039) | (n33938 & n34039);
  assign n36894 = n28152 & n28198;
  assign n36895 = (n28197 & n28198) | (n28197 & n36894) | (n28198 & n36894);
  assign n34044 = (n28198 & n33938) | (n28198 & n36895) | (n33938 & n36895);
  assign n28324 = ~n34040 & n34044;
  assign n36896 = n28024 | n28324;
  assign n36897 = (n28204 & n28324) | (n28204 & n36896) | (n28324 & n36896);
  assign n34046 = (n28324 & n36825) | (n28324 & n36897) | (n36825 & n36897);
  assign n36898 = n28187 & ~n33999;
  assign n36899 = n34002 & n36898;
  assign n36900 = ~n28187 & n33999;
  assign n36901 = (n28187 & n34002) | (n28187 & ~n36900) | (n34002 & ~n36900);
  assign n28328 = ~n36899 & n36901;
  assign n28329 = n33980 & n28328;
  assign n34047 = n28188 & n28328;
  assign n34048 = (n28188 & n33980) | (n28188 & n34047) | (n33980 & n34047);
  assign n28332 = ~n28329 & n34048;
  assign n34049 = n28332 | n34039;
  assign n34050 = n28197 | n28332;
  assign n34051 = (n33938 & n34049) | (n33938 & n34050) | (n34049 & n34050);
  assign n28335 = x141 & x164;
  assign n28336 = x140 & x165;
  assign n28337 = n28335 & n28336;
  assign n28338 = n28335 | n28336;
  assign n28339 = ~n28337 & n28338;
  assign n34054 = n28170 & n33995;
  assign n34055 = n28170 & n28177;
  assign n34056 = (n33915 & n34054) | (n33915 & n34055) | (n34054 & n34055);
  assign n37645 = n28170 & n28171;
  assign n37646 = (n28171 & n33995) | (n28171 & n37645) | (n33995 & n37645);
  assign n34058 = n28170 | n28177;
  assign n36903 = n28171 & n34058;
  assign n36904 = (n33915 & n37646) | (n33915 & n36903) | (n37646 & n36903);
  assign n28343 = ~n34056 & n36904;
  assign n34060 = n28343 | n33998;
  assign n28345 = x142 & x163;
  assign n28352 = x143 & x162;
  assign n34067 = n28352 & n36837;
  assign n36907 = n28352 & n36837;
  assign n36908 = (n28164 & n28352) | (n28164 & n36907) | (n28352 & n36907);
  assign n36910 = (n27967 & n34067) | (n27967 & n36908) | (n34067 & n36908);
  assign n37647 = n34067 | n36908;
  assign n37648 = (n27969 & n36910) | (n27969 & n37647) | (n36910 & n37647);
  assign n36911 = (n33895 & n37648) | (n33895 & n36910) | (n37648 & n36910);
  assign n34070 = n28352 | n36837;
  assign n36912 = n28352 | n36837;
  assign n36913 = n28164 | n36912;
  assign n36915 = (n27967 & n34070) | (n27967 & n36913) | (n34070 & n36913);
  assign n37649 = n34070 | n36913;
  assign n37650 = (n27969 & n36915) | (n27969 & n37649) | (n36915 & n37649);
  assign n36916 = (n33895 & n37650) | (n33895 & n36915) | (n37650 & n36915);
  assign n28355 = ~n36911 & n36916;
  assign n36918 = n27967 & n28164;
  assign n37651 = (n27969 & n28164) | (n27969 & n36918) | (n28164 & n36918);
  assign n36919 = (n33895 & n37651) | (n33895 & n36918) | (n37651 & n36918);
  assign n36921 = (n27967 & n28159) | (n27967 & n28165) | (n28159 & n28165);
  assign n37653 = (n27969 & n36921) | (n27969 & n28159) | (n36921 & n28159);
  assign n36922 = (n33895 & n37653) | (n33895 & n36921) | (n37653 & n36921);
  assign n28349 = ~n36919 & n36922;
  assign n34072 = n28349 & n28355;
  assign n36923 = (n28355 & n34054) | (n28355 & n34072) | (n34054 & n34072);
  assign n36924 = (n28355 & n34055) | (n28355 & n34072) | (n34055 & n34072);
  assign n36925 = (n33915 & n36923) | (n33915 & n36924) | (n36923 & n36924);
  assign n34074 = n28349 | n28355;
  assign n36926 = n34054 | n34074;
  assign n36927 = n34055 | n34074;
  assign n36928 = (n33915 & n36926) | (n33915 & n36927) | (n36926 & n36927);
  assign n28358 = ~n36925 & n36928;
  assign n28359 = n28345 & n28358;
  assign n28360 = n28345 | n28358;
  assign n28361 = ~n28359 & n28360;
  assign n36905 = n28343 | n36861;
  assign n36906 = (n28182 & n28343) | (n28182 & n36905) | (n28343 & n36905);
  assign n36929 = n28361 & n36906;
  assign n36930 = n28361 & n33833;
  assign n36931 = (n34060 & n36929) | (n34060 & n36930) | (n36929 & n36930);
  assign n36932 = n28361 | n36906;
  assign n36933 = n28361 | n33833;
  assign n36934 = (n34060 & n36932) | (n34060 & n36933) | (n36932 & n36933);
  assign n28364 = ~n36931 & n36934;
  assign n28365 = n28339 & n28364;
  assign n28366 = n28339 | n28364;
  assign n28367 = ~n28365 & n28366;
  assign n34052 = n36899 | n28328;
  assign n34076 = n28367 | n34052;
  assign n34077 = n36899 | n28367;
  assign n34078 = (n33980 & n34076) | (n33980 & n34077) | (n34076 & n34077);
  assign n34079 = n28367 & n34052;
  assign n34080 = n36899 & n28367;
  assign n34081 = (n33980 & n34079) | (n33980 & n34080) | (n34079 & n34080);
  assign n28370 = n34078 & ~n34081;
  assign n28371 = x139 & x166;
  assign n28372 = n28370 | n28371;
  assign n28373 = n28370 & n28371;
  assign n28374 = n28372 & ~n28373;
  assign n28375 = n34051 | n28374;
  assign n28376 = n34051 & n28374;
  assign n28377 = n28375 & ~n28376;
  assign n28378 = x138 & x167;
  assign n28379 = ~n28377 & n28378;
  assign n28380 = n28377 & ~n28378;
  assign n28381 = n28379 | n28380;
  assign n28382 = n34046 & n28381;
  assign n28383 = n34046 | n28381;
  assign n28384 = ~n28382 & n28383;
  assign n28385 = n28211 | n28384;
  assign n34082 = n28213 | n28385;
  assign n34083 = (n28385 & n33969) | (n28385 & n34082) | (n33969 & n34082);
  assign n34084 = n28211 | n33968;
  assign n28388 = n28212 & n28384;
  assign n34085 = n28030 | n28211;
  assign n36935 = n28388 & n34085;
  assign n36936 = n28388 & n33961;
  assign n36937 = (n34084 & n36935) | (n34084 & n36936) | (n36935 & n36936);
  assign n28390 = n34083 & ~n36937;
  assign n28391 = ~n28320 & n28390;
  assign n28392 = n28320 & ~n28390;
  assign n28393 = n28391 | n28392;
  assign n28394 = x136 & x169;
  assign n28395 = n28393 & n28394;
  assign n28396 = n28393 | n28394;
  assign n28397 = ~n28395 & n28396;
  assign n36872 = n33961 & n37636;
  assign n34008 = (n28033 & n28221) | (n28033 & ~n36872) | (n28221 & ~n36872);
  assign n37654 = n28218 | n34008;
  assign n37655 = (n28218 & n28220) | (n28218 & n37654) | (n28220 & n37654);
  assign n36939 = (n28218 & n34006) | (n28218 & n37655) | (n34006 & n37655);
  assign n28399 = ~n28397 & n36939;
  assign n28400 = n28397 & ~n36939;
  assign n28401 = n28399 | n28400;
  assign n28402 = x135 & x170;
  assign n28403 = n28401 & n28402;
  assign n28404 = n28401 | n28402;
  assign n28405 = ~n28403 & n28404;
  assign n28406 = n34038 | n28405;
  assign n28407 = n34038 & n28405;
  assign n28408 = n28406 & ~n28407;
  assign n28409 = n34036 & n28408;
  assign n28410 = n34036 | n28408;
  assign n28411 = ~n28409 & n28410;
  assign n28412 = x134 & x171;
  assign n28413 = n28411 & n28412;
  assign n28414 = n28411 | n28412;
  assign n28415 = ~n28413 & n28414;
  assign n28416 = x133 & x172;
  assign n28417 = n28415 & n28416;
  assign n28418 = n28415 | n28416;
  assign n28419 = ~n28417 & n28418;
  assign n28420 = n34034 | n28419;
  assign n28421 = n34034 & n28419;
  assign n28422 = n28420 & ~n28421;
  assign n28423 = x132 & x173;
  assign n28424 = ~n28422 & n28423;
  assign n28425 = n28422 & ~n28423;
  assign n28426 = n28424 | n28425;
  assign n28427 = ~n28298 & n28426;
  assign n28428 = n28298 & ~n28426;
  assign n28429 = n28427 | n28428;
  assign n28430 = n36887 | n28429;
  assign n28431 = n28274 | n28430;
  assign n28102 = n36811 & n28101;
  assign n28432 = n28072 | n36887;
  assign n28433 = n28102 | n28432;
  assign n28434 = n36885 & n28429;
  assign n28435 = n28433 & n28434;
  assign n28436 = n28431 & ~n28435;
  assign n28437 = x131 & x174;
  assign n28438 = n28436 & n28437;
  assign n28439 = n28436 | n28437;
  assign n28440 = ~n28438 & n28439;
  assign n28441 = n28278 | n28440;
  assign n28442 = n34020 | n28441;
  assign n28447 = x130 & x175;
  assign n34087 = n28104 | n28278;
  assign n36940 = n28080 | n34087;
  assign n36941 = (n33841 & n34087) | (n33841 & n36940) | (n34087 & n36940);
  assign n28444 = n28279 & n28440;
  assign n28445 = n36941 & n28444;
  assign n36942 = n28445 & ~n28447;
  assign n36943 = (n28442 & n28447) | (n28442 & ~n36942) | (n28447 & ~n36942);
  assign n36944 = ~n28445 & n28447;
  assign n36945 = n28442 & n36944;
  assign n28450 = n36943 & ~n36945;
  assign n34025 = n28285 & n28286;
  assign n36946 = n28450 & n34025;
  assign n36947 = n28285 & n28450;
  assign n36948 = (n34024 & n36946) | (n34024 & n36947) | (n36946 & n36947);
  assign n36949 = n28450 | n34025;
  assign n36950 = n28285 | n28450;
  assign n36951 = (n34024 & n36949) | (n34024 & n36950) | (n36949 & n36950);
  assign n28453 = ~n36948 & n36951;
  assign n34026 = (n28285 & n34024) | (n28285 & n34025) | (n34024 & n34025);
  assign n34091 = n28297 | n28422;
  assign n34092 = n28268 | n34091;
  assign n34093 = n28297 & n28422;
  assign n34094 = (n28268 & n28422) | (n28268 & n34093) | (n28422 & n34093);
  assign n28457 = n28423 & ~n34094;
  assign n28458 = n34092 & n28457;
  assign n34095 = n28434 | n28458;
  assign n34096 = (n28433 & n28458) | (n28433 & n34095) | (n28458 & n34095);
  assign n28462 = n28058 | n28316;
  assign n28463 = n28110 | n28462;
  assign n28464 = n28243 | n28315;
  assign n28465 = n28415 & n28464;
  assign n28466 = n28463 & n28465;
  assign n28467 = n28416 & ~n28466;
  assign n28460 = n28316 | n28415;
  assign n28461 = n28294 | n28460;
  assign n34097 = n28297 | n28461;
  assign n34098 = (n28297 & n28467) | (n28297 & n34097) | (n28467 & n34097);
  assign n28470 = n28268 | n34098;
  assign n28471 = n28461 & ~n28466;
  assign n28472 = n28416 | n28471;
  assign n28474 = n34038 | n28401;
  assign n28475 = n33959 | n34010;
  assign n28476 = n34012 & n28401;
  assign n28477 = n28475 & n28476;
  assign n28478 = n28474 & ~n28477;
  assign n28479 = n28402 & n28478;
  assign n34099 = n28408 | n28479;
  assign n34100 = (n28479 & n34036) | (n28479 & n34099) | (n34036 & n34099);
  assign n28229 = n28220 & n34008;
  assign n34101 = n28218 & n28393;
  assign n36952 = (n28229 & n28393) | (n28229 & n34101) | (n28393 & n34101);
  assign n36953 = n28393 & n34101;
  assign n36954 = (n34006 & n36952) | (n34006 & n36953) | (n36952 & n36953);
  assign n37656 = n28217 & n28394;
  assign n37657 = n28216 & n37656;
  assign n36956 = (n28393 & n28394) | (n28393 & n37657) | (n28394 & n37657);
  assign n36957 = (n28229 & n28394) | (n28229 & n36956) | (n28394 & n36956);
  assign n37826 = n28394 & n37656;
  assign n37827 = n28216 & n37826;
  assign n37659 = (n28393 & n28394) | (n28393 & n37827) | (n28394 & n37827);
  assign n36959 = (n34006 & n36957) | (n34006 & n37659) | (n36957 & n37659);
  assign n28484 = ~n36954 & n36959;
  assign n36960 = n28484 | n34012;
  assign n36961 = (n28401 & n28484) | (n28401 & n36960) | (n28484 & n36960);
  assign n34108 = (n28475 & n28484) | (n28475 & n36961) | (n28484 & n36961);
  assign n28486 = n28320 & n28390;
  assign n34110 = n28393 | n28486;
  assign n34165 = n28218 | n28486;
  assign n36962 = (n28393 & n28486) | (n28393 & n34165) | (n28486 & n34165);
  assign n36963 = (n28229 & n34110) | (n28229 & n36962) | (n34110 & n36962);
  assign n36964 = n34110 & n36962;
  assign n36965 = (n34006 & n36963) | (n34006 & n36964) | (n36963 & n36964);
  assign n34086 = (n33961 & n34084) | (n33961 & n34085) | (n34084 & n34085);
  assign n28489 = n34051 & n28370;
  assign n34112 = (n28371 & n28373) | (n28371 & n34051) | (n28373 & n34051);
  assign n28492 = ~n28489 & n34112;
  assign n34113 = n28377 | n28492;
  assign n36966 = (n28492 & n34113) | (n28492 & n36897) | (n34113 & n36897);
  assign n36967 = (n28324 & n28492) | (n28324 & n34113) | (n28492 & n34113);
  assign n36968 = (n36825 & n36966) | (n36825 & n36967) | (n36966 & n36967);
  assign n28494 = n28335 & n28364;
  assign n28495 = n28335 | n28364;
  assign n28496 = ~n28494 & n28495;
  assign n34115 = n28496 | n34052;
  assign n34116 = n36899 | n28496;
  assign n34117 = (n33980 & n34115) | (n33980 & n34116) | (n34115 & n34116);
  assign n34118 = n28496 & n34052;
  assign n34119 = n36899 & n28496;
  assign n34120 = (n33980 & n34118) | (n33980 & n34119) | (n34118 & n34119);
  assign n28499 = n28336 & ~n34120;
  assign n28500 = n34117 & n28499;
  assign n34121 = n28370 | n28500;
  assign n34122 = (n28500 & n34051) | (n28500 & n34121) | (n34051 & n34121);
  assign n28503 = x142 & x164;
  assign n28504 = x141 & x165;
  assign n28505 = n28503 & n28504;
  assign n28506 = n28503 | n28504;
  assign n28507 = ~n28505 & n28506;
  assign n28510 = x143 & x163;
  assign n37660 = n28510 & n37648;
  assign n37661 = n28510 & n36910;
  assign n37662 = (n33895 & n37660) | (n33895 & n37661) | (n37660 & n37661);
  assign n36970 = (n28510 & n34072) | (n28510 & n37662) | (n34072 & n37662);
  assign n36971 = (n28355 & n28510) | (n28355 & n37662) | (n28510 & n37662);
  assign n36972 = (n34054 & n36970) | (n34054 & n36971) | (n36970 & n36971);
  assign n36973 = (n34055 & n36970) | (n34055 & n36971) | (n36970 & n36971);
  assign n36974 = (n33915 & n36972) | (n33915 & n36973) | (n36972 & n36973);
  assign n37663 = n28510 | n37648;
  assign n37664 = n28510 | n36910;
  assign n37665 = (n33895 & n37663) | (n33895 & n37664) | (n37663 & n37664);
  assign n36976 = n34072 | n37665;
  assign n36977 = n28355 | n37665;
  assign n36978 = (n34054 & n36976) | (n34054 & n36977) | (n36976 & n36977);
  assign n36979 = (n34055 & n36976) | (n34055 & n36977) | (n36976 & n36977);
  assign n36980 = (n33915 & n36978) | (n33915 & n36979) | (n36978 & n36979);
  assign n28513 = ~n36974 & n36980;
  assign n34135 = n28359 & n28513;
  assign n36981 = (n28361 & n28513) | (n28361 & n34135) | (n28513 & n34135);
  assign n36982 = (n34135 & n36906) | (n34135 & n36981) | (n36906 & n36981);
  assign n36983 = (n33833 & n34135) | (n33833 & n36981) | (n34135 & n36981);
  assign n36984 = (n34060 & n36982) | (n34060 & n36983) | (n36982 & n36983);
  assign n34138 = n28359 | n28513;
  assign n36985 = n28361 | n34138;
  assign n36986 = (n34138 & n36906) | (n34138 & n36985) | (n36906 & n36985);
  assign n36987 = (n33833 & n34138) | (n33833 & n36985) | (n34138 & n36985);
  assign n36988 = (n34060 & n36986) | (n34060 & n36987) | (n36986 & n36987);
  assign n28516 = ~n36984 & n36988;
  assign n28517 = n28507 & n28516;
  assign n28518 = n28507 | n28516;
  assign n28519 = ~n28517 & n28518;
  assign n34140 = n28494 | n28519;
  assign n34141 = n34120 | n34140;
  assign n34142 = n28494 & n28519;
  assign n34143 = (n28519 & n34120) | (n28519 & n34142) | (n34120 & n34142);
  assign n28522 = n34141 & ~n34143;
  assign n28523 = x140 & x166;
  assign n28524 = n28522 | n28523;
  assign n28525 = n28522 & n28523;
  assign n28526 = n28524 & ~n28525;
  assign n28527 = n34122 | n28526;
  assign n28528 = n34122 & n28526;
  assign n28529 = n28527 & ~n28528;
  assign n28530 = x139 & x167;
  assign n28531 = n28529 | n28530;
  assign n28532 = n28529 & n28530;
  assign n28533 = n28531 & ~n28532;
  assign n28534 = n36968 | n28533;
  assign n28535 = n36968 & n28533;
  assign n28536 = n28534 & ~n28535;
  assign n36989 = n28377 | n36897;
  assign n36990 = n28324 | n28377;
  assign n36991 = (n36825 & n36989) | (n36825 & n36990) | (n36989 & n36990);
  assign n36992 = (n28378 & n28379) | (n28378 & ~n36897) | (n28379 & ~n36897);
  assign n37666 = ~n28324 & n28378;
  assign n37667 = (~n28377 & n28378) | (~n28377 & n37666) | (n28378 & n37666);
  assign n36994 = (~n36825 & n36992) | (~n36825 & n37667) | (n36992 & n37667);
  assign n28539 = n36991 & n36994;
  assign n36996 = n28536 & ~n28539;
  assign n37668 = ~n28388 & n36996;
  assign n36997 = (~n34086 & n37668) | (~n34086 & n36996) | (n37668 & n36996);
  assign n36999 = ~n28536 & n28539;
  assign n37669 = (n28388 & ~n28536) | (n28388 & n36999) | (~n28536 & n36999);
  assign n37000 = (n34086 & n37669) | (n34086 & n36999) | (n37669 & n36999);
  assign n28543 = n36997 | n37000;
  assign n28544 = x138 & x168;
  assign n28545 = n28543 & n28544;
  assign n28546 = n28543 | n28544;
  assign n28547 = ~n28545 & n28546;
  assign n28548 = x137 & x169;
  assign n28549 = n28547 & n28548;
  assign n28550 = n28547 | n28548;
  assign n28551 = ~n28549 & n28550;
  assign n28552 = n36965 | n28551;
  assign n28553 = n36965 & n28551;
  assign n28554 = n28552 & ~n28553;
  assign n28555 = x136 & x170;
  assign n28556 = n28554 | n28555;
  assign n28557 = n28554 & n28555;
  assign n28558 = n28556 & ~n28557;
  assign n28559 = ~n34108 & n28558;
  assign n28560 = n34108 & ~n28558;
  assign n28561 = n28559 | n28560;
  assign n28562 = x135 & x171;
  assign n28563 = n28561 & n28562;
  assign n28564 = n28561 | n28562;
  assign n28565 = ~n28563 & n28564;
  assign n28566 = n34100 | n28565;
  assign n28567 = n34100 & n28565;
  assign n28568 = n28566 & ~n28567;
  assign n28569 = x134 & x172;
  assign n28570 = ~n28568 & n28569;
  assign n28571 = n28568 & ~n28569;
  assign n28572 = n28570 | n28571;
  assign n34147 = ~n28413 & n28572;
  assign n34148 = ~n28466 & n34147;
  assign n34149 = n28413 & ~n28572;
  assign n34150 = (n28466 & ~n28572) | (n28466 & n34149) | (~n28572 & n34149);
  assign n28575 = n34148 | n34150;
  assign n28576 = n28472 & n28575;
  assign n28577 = n28470 & n28576;
  assign n28468 = n28461 & n28467;
  assign n28578 = n28468 | n28575;
  assign n28579 = n34094 | n28578;
  assign n28580 = ~n28577 & n28579;
  assign n28581 = x133 & x173;
  assign n28582 = n28580 | n28581;
  assign n28583 = n28580 & n28581;
  assign n28584 = n28582 & ~n28583;
  assign n28585 = n34096 & n28584;
  assign n28586 = n34096 | n28584;
  assign n28587 = ~n28585 & n28586;
  assign n28588 = x132 & x174;
  assign n28589 = n28587 | n28588;
  assign n28590 = n28587 & n28588;
  assign n28591 = n28589 & ~n28590;
  assign n28592 = n28438 | n28591;
  assign n28593 = n28445 | n28592;
  assign n28594 = n28278 | n28438;
  assign n37001 = n28594 | n34019;
  assign n37002 = n28280 | n28594;
  assign n37003 = (n28091 & n37001) | (n28091 & n37002) | (n37001 & n37002);
  assign n28596 = n28439 & n28591;
  assign n28597 = n37003 & n28596;
  assign n28598 = n28593 & ~n28597;
  assign n28599 = x131 & x175;
  assign n28600 = n28598 & n28599;
  assign n28601 = n28598 | n28599;
  assign n28602 = ~n28600 & n28601;
  assign n34089 = n36945 | n28450;
  assign n37004 = n28602 | n34089;
  assign n37005 = n28602 | n36945;
  assign n37006 = (n34026 & n37004) | (n34026 & n37005) | (n37004 & n37005);
  assign n37007 = n28602 & n34089;
  assign n37008 = n28602 & n36945;
  assign n37009 = (n34026 & n37007) | (n34026 & n37008) | (n37007 & n37008);
  assign n28605 = n37006 & ~n37009;
  assign n28606 = n28590 | n28597;
  assign n34151 = n28413 & n28568;
  assign n34152 = (n28466 & n28568) | (n28466 & n34151) | (n28568 & n34151);
  assign n34153 = n28413 | n28568;
  assign n34155 = n28569 & n34153;
  assign n34156 = (n28466 & n28569) | (n28466 & n34155) | (n28569 & n34155);
  assign n28610 = ~n34152 & n34156;
  assign n34157 = n28576 | n28610;
  assign n34158 = (n28470 & n28610) | (n28470 & n34157) | (n28610 & n34157);
  assign n28612 = n34100 | n28561;
  assign n28613 = n34036 | n28479;
  assign n28614 = n28402 | n28478;
  assign n28615 = n28561 & n28614;
  assign n28616 = n28613 & n28615;
  assign n28617 = n28612 & ~n28616;
  assign n28618 = n28562 & n28617;
  assign n34159 = n28618 | n34151;
  assign n34160 = n28568 | n28618;
  assign n34161 = (n28466 & n34159) | (n28466 & n34160) | (n34159 & n34160);
  assign n37010 = n28554 & n36961;
  assign n37011 = n28484 & n28554;
  assign n37012 = (n28475 & n37010) | (n28475 & n37011) | (n37010 & n37011);
  assign n37013 = (n28555 & n28557) | (n28555 & n36961) | (n28557 & n36961);
  assign n37670 = n28484 & n28555;
  assign n37671 = (n28554 & n28555) | (n28554 & n37670) | (n28555 & n37670);
  assign n37015 = (n28475 & n37013) | (n28475 & n37671) | (n37013 & n37671);
  assign n28623 = ~n37012 & n37015;
  assign n34163 = n28615 | n28623;
  assign n34164 = (n28613 & n28623) | (n28613 & n34163) | (n28623 & n34163);
  assign n28625 = n36965 | n28547;
  assign n37016 = n28229 | n34165;
  assign n37017 = (n34006 & n34165) | (n34006 & n37016) | (n34165 & n37016);
  assign n37672 = ~n28320 & n28548;
  assign n37673 = ~n28390 & n37672;
  assign n37019 = (~n28547 & n28548) | (~n28547 & n37673) | (n28548 & n37673);
  assign n34168 = (n28548 & ~n37017) | (n28548 & n37019) | (~n37017 & n37019);
  assign n28631 = n28625 & n34168;
  assign n34171 = n28529 & n34113;
  assign n34172 = n28492 & n28529;
  assign n34173 = (n34046 & n34171) | (n34046 & n34172) | (n34171 & n34172);
  assign n37022 = n28492 & n28530;
  assign n37023 = (n28529 & n28530) | (n28529 & n37022) | (n28530 & n37022);
  assign n34174 = n28529 | n34113;
  assign n34178 = n28530 & n34174;
  assign n34179 = (n34046 & n37023) | (n34046 & n34178) | (n37023 & n34178);
  assign n28637 = ~n34173 & n34179;
  assign n34145 = n28388 | n28539;
  assign n34180 = n28536 | n28637;
  assign n37024 = (n28637 & n34145) | (n28637 & n34180) | (n34145 & n34180);
  assign n37025 = (n28539 & n28637) | (n28539 & n34180) | (n28637 & n34180);
  assign n37026 = (n34086 & n37024) | (n34086 & n37025) | (n37024 & n37025);
  assign n34182 = n28522 & n34121;
  assign n34183 = n28500 & n28522;
  assign n34184 = (n34051 & n34182) | (n34051 & n34183) | (n34182 & n34183);
  assign n28644 = n28503 & n28516;
  assign n28645 = n28503 | n28516;
  assign n28646 = ~n28644 & n28645;
  assign n34191 = n28494 & n28646;
  assign n34192 = (n28646 & n34120) | (n28646 & n34191) | (n34120 & n34191);
  assign n37674 = n28335 & n28504;
  assign n37675 = n28364 & n37674;
  assign n37028 = (n28504 & n28646) | (n28504 & n37675) | (n28646 & n37675);
  assign n34196 = (n28504 & n34120) | (n28504 & n37028) | (n34120 & n37028);
  assign n28650 = ~n34192 & n34196;
  assign n28653 = x142 & x165;
  assign n28655 = x143 & x164;
  assign n34200 = n28655 & n36974;
  assign n34201 = (n28655 & n36984) | (n28655 & n34200) | (n36984 & n34200);
  assign n34202 = n28655 | n36974;
  assign n34203 = n36984 | n34202;
  assign n28658 = ~n34201 & n34203;
  assign n28659 = n28653 & n28658;
  assign n28660 = n28653 | n28658;
  assign n28661 = ~n28659 & n28660;
  assign n34198 = n28644 | n28646;
  assign n37031 = n28661 | n34198;
  assign n37029 = n28494 | n28644;
  assign n37030 = (n28644 & n28646) | (n28644 & n37029) | (n28646 & n37029);
  assign n37032 = n28661 | n37030;
  assign n37033 = (n34120 & n37031) | (n34120 & n37032) | (n37031 & n37032);
  assign n37034 = n28661 & n34198;
  assign n37035 = n28661 & n37030;
  assign n37036 = (n34120 & n37034) | (n34120 & n37035) | (n37034 & n37035);
  assign n28664 = n37033 & ~n37036;
  assign n28665 = x141 & x166;
  assign n28666 = ~n28664 & n28665;
  assign n28667 = n28664 & ~n28665;
  assign n28668 = n28666 | n28667;
  assign n37037 = n28650 | n28668;
  assign n37038 = n34184 | n37037;
  assign n37039 = n28650 & n28668;
  assign n37040 = (n28668 & n34184) | (n28668 & n37039) | (n34184 & n37039);
  assign n28671 = n37038 & ~n37040;
  assign n34185 = n28522 | n34121;
  assign n34186 = n28500 | n28522;
  assign n34187 = (n34051 & n34185) | (n34051 & n34186) | (n34185 & n34186);
  assign n28641 = ~n34184 & n34187;
  assign n28672 = n28523 | n28641;
  assign n28673 = n28671 & n28672;
  assign n28642 = n28523 & n28641;
  assign n34189 = n28492 | n28642;
  assign n37041 = n28673 & n34189;
  assign n34188 = n28642 | n34113;
  assign n37042 = n28673 & n34188;
  assign n37043 = (n34046 & n37041) | (n34046 & n37042) | (n37041 & n37042);
  assign n28675 = n28642 | n28671;
  assign n37044 = n28675 | n34172;
  assign n37045 = n28675 | n34171;
  assign n37046 = (n34046 & n37044) | (n34046 & n37045) | (n37044 & n37045);
  assign n28677 = ~n37043 & n37046;
  assign n28678 = x140 & x167;
  assign n28679 = n28677 & n28678;
  assign n28680 = n28677 | n28678;
  assign n28681 = ~n28679 & n28680;
  assign n28682 = ~n37026 & n28681;
  assign n28683 = n37026 & ~n28681;
  assign n28684 = n28682 | n28683;
  assign n28685 = x139 & x168;
  assign n28686 = x138 & x169;
  assign n28687 = n28685 & n28686;
  assign n28688 = n28685 | n28686;
  assign n28689 = ~n28687 & n28688;
  assign n28690 = n28684 & n28689;
  assign n28691 = n28684 | n28689;
  assign n28692 = ~n28690 & n28691;
  assign n28627 = n28320 | n28390;
  assign n37020 = n28545 | n28627;
  assign n37021 = (n28545 & n28547) | (n28545 & n37020) | (n28547 & n37020);
  assign n37047 = n28692 & ~n37021;
  assign n37048 = ~n28545 & n28692;
  assign n37049 = (~n37017 & n37047) | (~n37017 & n37048) | (n37047 & n37048);
  assign n37050 = ~n28692 & n37021;
  assign n37051 = n28545 & ~n28692;
  assign n37052 = (n37017 & n37050) | (n37017 & n37051) | (n37050 & n37051);
  assign n28695 = n37049 | n37052;
  assign n28696 = n28631 | n28695;
  assign n34204 = n28554 | n28696;
  assign n34205 = (n28696 & n34108) | (n28696 & n34204) | (n34108 & n34204);
  assign n28698 = n28484 | n28631;
  assign n34206 = n28476 | n28698;
  assign n34207 = (n28475 & n28698) | (n28475 & n34206) | (n28698 & n34206);
  assign n28628 = n28547 & n28627;
  assign n28629 = n37017 & n28628;
  assign n28700 = n28625 & ~n28629;
  assign n28701 = n28548 | n28700;
  assign n28702 = n28695 & n28701;
  assign n28703 = n34207 & n28702;
  assign n28704 = n34205 & ~n28703;
  assign n28705 = x137 & x170;
  assign n28706 = n28704 | n28705;
  assign n28707 = n28704 & n28705;
  assign n28708 = n28706 & ~n28707;
  assign n28709 = n34164 & n28708;
  assign n28710 = n34164 | n28708;
  assign n28711 = ~n28709 & n28710;
  assign n28712 = x136 & x171;
  assign n28713 = n28711 & n28712;
  assign n28714 = n28711 | n28712;
  assign n28715 = ~n28713 & n28714;
  assign n28716 = x135 & x172;
  assign n28717 = n28715 & n28716;
  assign n28718 = n28715 | n28716;
  assign n28719 = ~n28717 & n28718;
  assign n28720 = ~n34161 & n28719;
  assign n28721 = n34161 & ~n28719;
  assign n28722 = n28720 | n28721;
  assign n28723 = x134 & x173;
  assign n28724 = n28722 | n28723;
  assign n28725 = n28722 & n28723;
  assign n28726 = n28724 & ~n28725;
  assign n28727 = ~n34158 & n28726;
  assign n28728 = n34158 & ~n28726;
  assign n28729 = n28727 | n28728;
  assign n28730 = n28583 | n28729;
  assign n28731 = n28585 | n28730;
  assign n28732 = n28458 | n28583;
  assign n28733 = n28435 | n28732;
  assign n28734 = n28582 & n28729;
  assign n28735 = n28733 & n28734;
  assign n28736 = n28731 & ~n28735;
  assign n28737 = x133 & x174;
  assign n28738 = n28736 & n28737;
  assign n28739 = n28736 | n28737;
  assign n28740 = ~n28738 & n28739;
  assign n28741 = x132 & x175;
  assign n28742 = n28740 & ~n28741;
  assign n28743 = ~n28740 & n28741;
  assign n28744 = n28742 | n28743;
  assign n28745 = n28606 & n28744;
  assign n28746 = n28606 | n28744;
  assign n28747 = ~n28745 & n28746;
  assign n28748 = n28600 | n28747;
  assign n28749 = n37009 | n28748;
  assign n28750 = n36945 | n28600;
  assign n28751 = n36948 | n28750;
  assign n28752 = n28601 & n28747;
  assign n28753 = n28751 & n28752;
  assign n28754 = n28749 & ~n28753;
  assign n34208 = n28590 & n28740;
  assign n34209 = (n28597 & n28740) | (n28597 & n34208) | (n28740 & n34208);
  assign n34210 = n28590 | n28740;
  assign n34211 = n28597 | n34210;
  assign n28757 = n28741 & n34211;
  assign n28758 = ~n34209 & n28757;
  assign n34212 = n28752 | n28758;
  assign n34213 = (n28751 & n28758) | (n28751 & n34212) | (n28758 & n34212);
  assign n28760 = n34158 & n28722;
  assign n34214 = (n28723 & n28725) | (n28723 & n34158) | (n28725 & n34158);
  assign n28763 = ~n28760 & n34214;
  assign n37053 = n28582 | n28763;
  assign n37054 = (n28729 & n28763) | (n28729 & n37053) | (n28763 & n37053);
  assign n34216 = (n28733 & n28763) | (n28733 & n37054) | (n28763 & n37054);
  assign n34217 = n28413 | n28618;
  assign n34218 = n28466 | n34217;
  assign n28766 = n28562 | n28617;
  assign n28767 = n28715 & n28766;
  assign n28768 = n34218 & n28767;
  assign n28769 = n34161 | n28715;
  assign n28770 = ~n28768 & n28769;
  assign n28771 = n28716 & n28770;
  assign n28772 = n34158 | n28771;
  assign n28773 = n28713 | n28768;
  assign n28774 = n28684 & n28685;
  assign n28775 = n28684 | n28685;
  assign n28776 = ~n28774 & n28775;
  assign n37055 = n28776 & n37021;
  assign n37056 = n28545 & n28776;
  assign n37057 = (n37017 & n37055) | (n37017 & n37056) | (n37055 & n37056);
  assign n34170 = (n28545 & n37017) | (n28545 & n37021) | (n37017 & n37021);
  assign n34219 = n28686 & n28776;
  assign n34220 = (n28686 & n34170) | (n28686 & n34219) | (n34170 & n34219);
  assign n28780 = ~n37057 & n34220;
  assign n34221 = n28702 | n28780;
  assign n34222 = (n28780 & n34207) | (n28780 & n34221) | (n34207 & n34221);
  assign n28782 = x139 & x169;
  assign n28783 = x138 & x170;
  assign n28784 = n28782 & n28783;
  assign n28785 = n28782 | n28783;
  assign n28786 = ~n28784 & n28785;
  assign n28788 = x140 & x168;
  assign n34225 = n28679 | n34180;
  assign n34226 = n28637 | n28679;
  assign n37058 = (n34145 & n34225) | (n34145 & n34226) | (n34225 & n34226);
  assign n37059 = (n28539 & n34225) | (n28539 & n34226) | (n34225 & n34226);
  assign n37060 = (n34086 & n37058) | (n34086 & n37059) | (n37058 & n37059);
  assign n34190 = (n34046 & n34188) | (n34046 & n34189) | (n34188 & n34189);
  assign n34228 = n28650 & n28664;
  assign n34229 = (n28664 & n34184) | (n28664 & n34228) | (n34184 & n34228);
  assign n34230 = n28650 | n28664;
  assign n34232 = n28665 & n34230;
  assign n34233 = (n28665 & n34184) | (n28665 & n34232) | (n34184 & n34232);
  assign n28794 = ~n34229 & n34233;
  assign n28801 = x142 & x166;
  assign n28803 = x143 & x165;
  assign n37069 = n28655 & n28803;
  assign n37676 = n36974 & n37069;
  assign n37070 = (n36984 & n37676) | (n36984 & n37069) | (n37676 & n37069);
  assign n37067 = (n28658 & n28803) | (n28658 & n37070) | (n28803 & n37070);
  assign n37071 = (n34198 & n37067) | (n34198 & n37070) | (n37067 & n37070);
  assign n37072 = (n37030 & n37067) | (n37030 & n37070) | (n37067 & n37070);
  assign n37073 = (n34120 & n37071) | (n34120 & n37072) | (n37071 & n37072);
  assign n37076 = n28655 | n28803;
  assign n37677 = (n28803 & n36974) | (n28803 & n37076) | (n36974 & n37076);
  assign n37077 = (n36984 & n37677) | (n36984 & n37076) | (n37677 & n37076);
  assign n37074 = n28658 | n37077;
  assign n37078 = (n34198 & n37074) | (n34198 & n37077) | (n37074 & n37077);
  assign n37079 = (n37030 & n37074) | (n37030 & n37077) | (n37074 & n37077);
  assign n37080 = (n34120 & n37078) | (n34120 & n37079) | (n37078 & n37079);
  assign n28806 = ~n37073 & n37080;
  assign n28807 = n28801 & n28806;
  assign n28808 = n28801 | n28806;
  assign n28809 = ~n28807 & n28808;
  assign n37678 = n28644 & n28658;
  assign n37679 = (n28646 & n28658) | (n28646 & n37678) | (n28658 & n37678);
  assign n37062 = n28658 & n37030;
  assign n37063 = (n34120 & n37679) | (n34120 & n37062) | (n37679 & n37062);
  assign n37064 = (n28653 & n28659) | (n28653 & n34198) | (n28659 & n34198);
  assign n37065 = (n28653 & n28659) | (n28653 & n37030) | (n28659 & n37030);
  assign n37066 = (n34120 & n37064) | (n34120 & n37065) | (n37064 & n37065);
  assign n28799 = ~n37063 & n37066;
  assign n34237 = n28799 | n34228;
  assign n37081 = n28809 | n34237;
  assign n34238 = n28664 | n28799;
  assign n37082 = n28809 | n34238;
  assign n37083 = (n34184 & n37081) | (n34184 & n37082) | (n37081 & n37082);
  assign n37084 = n28809 & n34237;
  assign n37085 = n28809 & n34238;
  assign n37086 = (n34184 & n37084) | (n34184 & n37085) | (n37084 & n37085);
  assign n28812 = n37083 & ~n37086;
  assign n37088 = ~n28794 & n28812;
  assign n37680 = ~n28673 & n37088;
  assign n37089 = (~n34190 & n37680) | (~n34190 & n37088) | (n37680 & n37088);
  assign n37091 = n28794 & ~n28812;
  assign n37681 = (n28673 & ~n28812) | (n28673 & n37091) | (~n28812 & n37091);
  assign n37092 = (n34190 & n37681) | (n34190 & n37091) | (n37681 & n37091);
  assign n28815 = n37089 | n37092;
  assign n28816 = x141 & x167;
  assign n28817 = n28815 & n28816;
  assign n28818 = n28815 | n28816;
  assign n28819 = ~n28817 & n28818;
  assign n37093 = n28680 & n28819;
  assign n37094 = n37060 & n37093;
  assign n37095 = n28680 | n28819;
  assign n37096 = (n28819 & n37060) | (n28819 & n37095) | (n37060 & n37095);
  assign n28822 = ~n37094 & n37096;
  assign n28823 = n28788 & n28822;
  assign n28824 = n28788 | n28822;
  assign n28825 = ~n28823 & n28824;
  assign n34223 = n28774 | n28776;
  assign n34248 = n28825 & n34223;
  assign n34249 = n28774 & n28825;
  assign n34250 = (n34170 & n34248) | (n34170 & n34249) | (n34248 & n34249);
  assign n34251 = n28825 | n34223;
  assign n34252 = n28774 | n28825;
  assign n34253 = (n34170 & n34251) | (n34170 & n34252) | (n34251 & n34252);
  assign n28828 = ~n34250 & n34253;
  assign n28829 = ~n28786 & n28828;
  assign n28830 = n28786 & ~n28828;
  assign n28831 = n28829 | n28830;
  assign n28832 = n34222 | n28831;
  assign n28833 = n34222 & n28831;
  assign n28834 = n28832 & ~n28833;
  assign n28835 = n28707 | n28834;
  assign n34254 = n28708 | n28835;
  assign n34255 = (n28835 & n34164) | (n28835 & n34254) | (n34164 & n34254);
  assign n28838 = n28706 & n28834;
  assign n34256 = n28707 & n28838;
  assign n34257 = (n28838 & n34164) | (n28838 & n34256) | (n34164 & n34256);
  assign n28840 = n34255 & ~n34257;
  assign n28841 = x137 & x171;
  assign n28842 = n28840 & n28841;
  assign n28843 = n28840 | n28841;
  assign n28844 = ~n28842 & n28843;
  assign n28845 = x136 & x172;
  assign n28846 = n28844 & ~n28845;
  assign n28847 = ~n28844 & n28845;
  assign n28848 = n28846 | n28847;
  assign n28849 = ~n28773 & n28848;
  assign n28850 = n28773 & ~n28848;
  assign n28851 = n28849 | n28850;
  assign n28852 = n28716 | n28770;
  assign n28853 = n28851 & n28852;
  assign n28854 = n28772 & n28853;
  assign n28855 = n28771 | n28851;
  assign n28856 = n28760 | n28855;
  assign n28857 = ~n28854 & n28856;
  assign n28858 = x135 & x173;
  assign n28859 = n28857 | n28858;
  assign n28860 = n28857 & n28858;
  assign n28861 = n28859 & ~n28860;
  assign n28862 = n34216 & n28861;
  assign n28863 = n34216 | n28861;
  assign n28864 = ~n28862 & n28863;
  assign n28865 = x134 & x174;
  assign n28866 = n28864 & n28865;
  assign n28867 = n28864 | n28865;
  assign n28868 = ~n28866 & n28867;
  assign n28869 = n28738 | n28868;
  assign n28870 = n34209 | n28869;
  assign n28871 = n28590 | n28738;
  assign n28872 = n28597 | n28871;
  assign n28873 = n28739 & n28868;
  assign n28874 = n28872 & n28873;
  assign n28875 = n28870 & ~n28874;
  assign n28876 = x133 & x175;
  assign n28877 = n28875 & n28876;
  assign n28878 = n28875 | n28876;
  assign n28879 = ~n28877 & n28878;
  assign n28880 = n34213 | n28879;
  assign n28881 = n34213 & n28879;
  assign n28882 = n28880 & ~n28881;
  assign n34258 = n28860 | n28861;
  assign n34259 = (n28860 & n34216) | (n28860 & n34258) | (n34216 & n34258);
  assign n29001 = n28713 | n28842;
  assign n37097 = (n28842 & n28844) | (n28842 & n29001) | (n28844 & n29001);
  assign n34267 = n28842 | n28844;
  assign n34268 = (n28768 & n37097) | (n28768 & n34267) | (n37097 & n34267);
  assign n28902 = x139 & x170;
  assign n28906 = x140 & x169;
  assign n28790 = n28680 & n37060;
  assign n34234 = n28673 | n28794;
  assign n34235 = (n28794 & n34190) | (n28794 & n34234) | (n34190 & n34234);
  assign n28910 = x143 & x166;
  assign n34278 = n28910 & n37073;
  assign n37098 = n28910 & n37073;
  assign n37099 = (n28806 & n28910) | (n28806 & n37098) | (n28910 & n37098);
  assign n37100 = (n34237 & n34278) | (n34237 & n37099) | (n34278 & n37099);
  assign n37101 = (n34238 & n34278) | (n34238 & n37099) | (n34278 & n37099);
  assign n37102 = (n34184 & n37100) | (n34184 & n37101) | (n37100 & n37101);
  assign n34281 = n28910 | n37073;
  assign n37103 = n28910 | n37073;
  assign n37104 = n28806 | n37103;
  assign n37105 = (n34237 & n34281) | (n34237 & n37104) | (n34281 & n37104);
  assign n37106 = (n34238 & n34281) | (n34238 & n37104) | (n34281 & n37104);
  assign n37107 = (n34184 & n37105) | (n34184 & n37106) | (n37105 & n37106);
  assign n28913 = ~n37102 & n37107;
  assign n28914 = x142 & x167;
  assign n28915 = n28913 & ~n28914;
  assign n28916 = ~n28913 & n28914;
  assign n28917 = n28915 | n28916;
  assign n37682 = n28799 | n28806;
  assign n37683 = n34228 | n37682;
  assign n37109 = n28806 | n34238;
  assign n37110 = (n34184 & n37683) | (n34184 & n37109) | (n37683 & n37109);
  assign n34283 = n28801 & ~n28806;
  assign n37111 = (n28801 & ~n34237) | (n28801 & n34283) | (~n34237 & n34283);
  assign n37112 = (n28801 & ~n34238) | (n28801 & n34283) | (~n34238 & n34283);
  assign n37113 = (~n34184 & n37111) | (~n34184 & n37112) | (n37111 & n37112);
  assign n28921 = n37110 & n37113;
  assign n34285 = n28812 | n28921;
  assign n34287 = n28917 & n34285;
  assign n34288 = n28917 & n28921;
  assign n34289 = (n34235 & n34287) | (n34235 & n34288) | (n34287 & n34288);
  assign n34290 = n28917 | n34285;
  assign n34291 = n28917 | n28921;
  assign n34292 = (n34235 & n34290) | (n34235 & n34291) | (n34290 & n34291);
  assign n28925 = ~n34289 & n34292;
  assign n28926 = x141 & x168;
  assign n28927 = n28925 & n28926;
  assign n28928 = n28925 | n28926;
  assign n28929 = ~n28927 & n28928;
  assign n34273 = n28817 | n28819;
  assign n37114 = n28929 & n34273;
  assign n37115 = n28817 & n28929;
  assign n37116 = (n28790 & n37114) | (n28790 & n37115) | (n37114 & n37115);
  assign n37117 = n28929 | n34273;
  assign n37118 = n28817 | n28929;
  assign n37119 = (n28790 & n37117) | (n28790 & n37118) | (n37117 & n37118);
  assign n28932 = ~n37116 & n37119;
  assign n28933 = n28906 & n28932;
  assign n28934 = n28906 | n28932;
  assign n28935 = ~n28933 & n28934;
  assign n34293 = n28823 | n28935;
  assign n34294 = n34250 | n34293;
  assign n34295 = n28823 & n28935;
  assign n34296 = (n28935 & n34250) | (n28935 & n34295) | (n34250 & n34295);
  assign n28938 = n34294 & ~n34296;
  assign n34224 = (n28774 & n34170) | (n28774 & n34223) | (n34170 & n34223);
  assign n28891 = n28782 | n28825;
  assign n28892 = n28782 & n28825;
  assign n28893 = n28891 & ~n28892;
  assign n28894 = n34224 | n28893;
  assign n28895 = n34224 & n28893;
  assign n28896 = n28894 & ~n28895;
  assign n28903 = n28782 & n28828;
  assign n34271 = n28896 | n28903;
  assign n34297 = n28938 | n34271;
  assign n34298 = n28903 | n28938;
  assign n34299 = (n34222 & n34297) | (n34222 & n34298) | (n34297 & n34298);
  assign n34300 = n28938 & n34271;
  assign n34301 = n28903 & n28938;
  assign n34302 = (n34222 & n34300) | (n34222 & n34301) | (n34300 & n34301);
  assign n28941 = n34299 & ~n34302;
  assign n28942 = n28902 & n28941;
  assign n28943 = n28902 | n28941;
  assign n28944 = ~n28942 & n28943;
  assign n28897 = n34222 & n28896;
  assign n34269 = n28783 & n28896;
  assign n34270 = (n28783 & n34222) | (n28783 & n34269) | (n34222 & n34269);
  assign n28900 = ~n28897 & n34270;
  assign n34303 = n28900 & n28944;
  assign n34304 = (n28944 & n34257) | (n28944 & n34303) | (n34257 & n34303);
  assign n34305 = n28900 | n28944;
  assign n34306 = n34257 | n34305;
  assign n28947 = ~n34304 & n34306;
  assign n28948 = x138 & x171;
  assign n28949 = n28947 & n28948;
  assign n28950 = n28947 | n28948;
  assign n28951 = ~n28949 & n28950;
  assign n28952 = x137 & x172;
  assign n28953 = n28951 & n28952;
  assign n28954 = n28951 | n28952;
  assign n28955 = ~n28953 & n28954;
  assign n28956 = n34268 | n28955;
  assign n28957 = n34268 & n28955;
  assign n28958 = n28956 & ~n28957;
  assign n34260 = n28713 & n28844;
  assign n34261 = (n28768 & n28844) | (n28768 & n34260) | (n28844 & n34260);
  assign n37684 = n28712 & n28845;
  assign n37685 = n28711 & n37684;
  assign n37121 = (n28844 & n28845) | (n28844 & n37685) | (n28845 & n37685);
  assign n34265 = (n28768 & n28845) | (n28768 & n37121) | (n28845 & n37121);
  assign n28888 = ~n34261 & n34265;
  assign n34307 = n28888 & n28958;
  assign n34308 = (n28854 & n28958) | (n28854 & n34307) | (n28958 & n34307);
  assign n34309 = n28888 | n28958;
  assign n34310 = n28854 | n34309;
  assign n28961 = ~n34308 & n34310;
  assign n28962 = x136 & x173;
  assign n28963 = n28961 & n28962;
  assign n28964 = n28961 | n28962;
  assign n28965 = ~n28963 & n28964;
  assign n28966 = n34259 | n28965;
  assign n28967 = n34259 & n28965;
  assign n28968 = n28966 & ~n28967;
  assign n28969 = x135 & x174;
  assign n28970 = n28968 & ~n28969;
  assign n28971 = ~n28968 & n28969;
  assign n28972 = n28970 | n28971;
  assign n34311 = n28866 & n28972;
  assign n34312 = (n28874 & n28972) | (n28874 & n34311) | (n28972 & n34311);
  assign n34313 = n28866 | n28972;
  assign n34314 = n28874 | n34313;
  assign n28975 = ~n34312 & n34314;
  assign n28976 = x134 & x175;
  assign n28977 = n28975 & n28976;
  assign n28978 = n28975 | n28976;
  assign n28979 = ~n28977 & n28978;
  assign n28980 = n28877 | n28979;
  assign n28981 = n28881 | n28980;
  assign n28982 = n28758 | n28877;
  assign n28983 = n28753 | n28982;
  assign n28883 = n28866 | n28874;
  assign n28984 = n28972 & ~n28976;
  assign n28985 = ~n28972 & n28976;
  assign n28986 = n28984 | n28985;
  assign n28987 = n28883 & n28986;
  assign n28988 = n28883 | n28986;
  assign n28989 = ~n28987 & n28988;
  assign n28990 = n28878 & n28989;
  assign n28991 = n28983 & n28990;
  assign n28992 = n28981 & ~n28991;
  assign n34315 = n28977 | n28990;
  assign n34316 = (n28977 & n28983) | (n28977 & n34315) | (n28983 & n34315);
  assign n34317 = n28763 | n28858;
  assign n34318 = (n28763 & n28857) | (n28763 & n34317) | (n28857 & n34317);
  assign n34319 = n28734 | n34318;
  assign n34320 = (n28733 & n34318) | (n28733 & n34319) | (n34318 & n34319);
  assign n28996 = n28859 & n34320;
  assign n34321 = n28963 | n28965;
  assign n34322 = (n28963 & n28996) | (n28963 & n34321) | (n28996 & n34321);
  assign n28999 = n28842 | n28951;
  assign n29000 = n34261 | n28999;
  assign n29003 = n28902 & ~n28948;
  assign n29004 = ~n28902 & n28948;
  assign n29005 = n29003 | n29004;
  assign n29006 = n28941 & n29005;
  assign n29007 = n28941 | n29005;
  assign n29008 = ~n29006 & n29007;
  assign n34323 = n28900 & n29008;
  assign n34324 = (n29008 & n34257) | (n29008 & n34323) | (n34257 & n34323);
  assign n34325 = n28900 | n29008;
  assign n34326 = n34257 | n34325;
  assign n34327 = ~n34324 & n34326;
  assign n34328 = n28843 & n34327;
  assign n34329 = n29001 & n34328;
  assign n37122 = ~n28952 & n34329;
  assign n37123 = ~n28952 & n34328;
  assign n37124 = (n28768 & n37122) | (n28768 & n37123) | (n37122 & n37123);
  assign n34335 = (n28952 & n29000) | (n28952 & ~n37124) | (n29000 & ~n37124);
  assign n34336 = n28949 | n34329;
  assign n34337 = n28949 | n34328;
  assign n34338 = (n28768 & n34336) | (n28768 & n34337) | (n34336 & n34337);
  assign n34339 = n28823 | n28932;
  assign n34340 = n34250 | n34339;
  assign n29023 = n28824 & n28932;
  assign n34344 = n28906 & ~n29023;
  assign n34342 = n28774 | n28823;
  assign n37125 = n28776 | n34342;
  assign n37126 = (n28906 & n34344) | (n28906 & ~n37125) | (n34344 & ~n37125);
  assign n37127 = (n28906 & ~n34342) | (n28906 & n34344) | (~n34342 & n34344);
  assign n37128 = (~n34170 & n37126) | (~n34170 & n37127) | (n37126 & n37127);
  assign n29026 = n34340 & n37128;
  assign n34343 = (n34170 & n37125) | (n34170 & n34342) | (n37125 & n34342);
  assign n34274 = (n28790 & n28817) | (n28790 & n34273) | (n28817 & n34273);
  assign n29038 = x142 & x168;
  assign n34354 = n28913 & n28921;
  assign n34362 = n37102 | n34354;
  assign n37129 = n28913 | n37102;
  assign n37130 = (n34285 & n37102) | (n34285 & n37129) | (n37102 & n37129);
  assign n37131 = (n34234 & n34362) | (n34234 & n37130) | (n34362 & n37130);
  assign n37132 = (n28794 & n34362) | (n28794 & n37130) | (n34362 & n37130);
  assign n37133 = (n34190 & n37131) | (n34190 & n37132) | (n37131 & n37132);
  assign n29040 = x143 & x167;
  assign n29041 = n37133 & n29040;
  assign n29042 = n37133 | n29040;
  assign n29043 = ~n29041 & n29042;
  assign n29044 = ~n29038 & n29043;
  assign n29045 = n29038 & ~n29043;
  assign n29046 = n29044 | n29045;
  assign n34350 = n28913 | n34285;
  assign n34351 = n28913 | n28921;
  assign n37134 = (n34234 & n34350) | (n34234 & n34351) | (n34350 & n34351);
  assign n37135 = (n28794 & n34350) | (n28794 & n34351) | (n34350 & n34351);
  assign n37136 = (n34190 & n37134) | (n34190 & n37135) | (n37134 & n37135);
  assign n34357 = n28914 & ~n34354;
  assign n37137 = (n28914 & n28916) | (n28914 & ~n34285) | (n28916 & ~n34285);
  assign n37138 = (~n34234 & n34357) | (~n34234 & n37137) | (n34357 & n37137);
  assign n37139 = (~n28794 & n34357) | (~n28794 & n37137) | (n34357 & n37137);
  assign n37140 = (~n34190 & n37138) | (~n34190 & n37139) | (n37138 & n37139);
  assign n29036 = n37136 & n37140;
  assign n34359 = n28925 | n29036;
  assign n34364 = n29046 | n34359;
  assign n34365 = n29036 | n29046;
  assign n34366 = (n34274 & n34364) | (n34274 & n34365) | (n34364 & n34365);
  assign n34367 = n29046 & n34359;
  assign n34368 = n29036 & n29046;
  assign n34369 = (n34274 & n34367) | (n34274 & n34368) | (n34367 & n34368);
  assign n29049 = n34366 & ~n34369;
  assign n29050 = x141 & x169;
  assign n29051 = n29049 | n29050;
  assign n29052 = n29049 & n29050;
  assign n29053 = n29051 & ~n29052;
  assign n37142 = n28817 | n28925;
  assign n37686 = n28819 | n37142;
  assign n37143 = (n28790 & n37686) | (n28790 & n37142) | (n37686 & n37142);
  assign n34346 = ~n28925 & n28926;
  assign n37144 = (n28926 & ~n34273) | (n28926 & n34346) | (~n34273 & n34346);
  assign n37145 = (~n28817 & n28926) | (~n28817 & n34346) | (n28926 & n34346);
  assign n37146 = (~n28790 & n37144) | (~n28790 & n37145) | (n37144 & n37145);
  assign n29031 = n37143 & n37146;
  assign n34348 = n29023 | n29031;
  assign n34370 = n29053 | n34348;
  assign n34371 = n29031 | n29053;
  assign n34372 = (n34343 & n34370) | (n34343 & n34371) | (n34370 & n34371);
  assign n34373 = n29053 & n34348;
  assign n34374 = n29031 & n29053;
  assign n34375 = (n34343 & n34373) | (n34343 & n34374) | (n34373 & n34374);
  assign n29056 = n34372 & ~n34375;
  assign n29057 = x140 & x170;
  assign n29058 = n29056 | n29057;
  assign n29059 = n29056 & n29057;
  assign n29060 = n29058 & ~n29059;
  assign n34376 = n29026 | n29060;
  assign n34377 = n34302 | n34376;
  assign n34378 = n29026 & n29060;
  assign n34379 = (n29060 & n34302) | (n29060 & n34378) | (n34302 & n34378);
  assign n29063 = n34377 & ~n34379;
  assign n29064 = x139 & x171;
  assign n29065 = n29063 | n29064;
  assign n29066 = n29063 & n29064;
  assign n29067 = n29065 & ~n29066;
  assign n34380 = n28942 | n29067;
  assign n34381 = n34304 | n34380;
  assign n34382 = n28942 & n29067;
  assign n34383 = (n29067 & n34304) | (n29067 & n34382) | (n34304 & n34382);
  assign n29071 = n34381 & ~n34383;
  assign n29072 = x138 & x172;
  assign n29073 = ~n29071 & n29072;
  assign n29074 = n29071 & ~n29072;
  assign n29075 = n29073 | n29074;
  assign n29076 = ~n34338 & n29075;
  assign n29077 = n34338 & ~n29075;
  assign n29078 = n29076 | n29077;
  assign n29079 = n34335 & n29078;
  assign n34331 = n28952 & ~n34329;
  assign n34332 = n28952 & ~n34328;
  assign n34333 = (~n28768 & n34331) | (~n28768 & n34332) | (n34331 & n34332);
  assign n29015 = n29000 & n34333;
  assign n29016 = n28888 | n29015;
  assign n34384 = n29016 & n29079;
  assign n34385 = (n28854 & n29079) | (n28854 & n34384) | (n29079 & n34384);
  assign n29081 = n29015 | n29078;
  assign n34386 = n29081 | n34307;
  assign n34387 = n28958 | n29081;
  assign n34388 = (n28854 & n34386) | (n28854 & n34387) | (n34386 & n34387);
  assign n29083 = ~n34385 & n34388;
  assign n29084 = x137 & x173;
  assign n29085 = n29083 | n29084;
  assign n29086 = n29083 & n29084;
  assign n29087 = n29085 & ~n29086;
  assign n29088 = n34322 & n29087;
  assign n29089 = n34322 | n29087;
  assign n29090 = ~n29088 & n29089;
  assign n29091 = x136 & x174;
  assign n29092 = n29090 & n29091;
  assign n29093 = n29090 | n29091;
  assign n29094 = ~n29092 & n29093;
  assign n28997 = n28965 & n28996;
  assign n29095 = n28966 & ~n28997;
  assign n29096 = n28969 & n29095;
  assign n29097 = n29094 | n29096;
  assign n29098 = n34312 | n29097;
  assign n29099 = n28866 | n29096;
  assign n29100 = n28874 | n29099;
  assign n29101 = n28969 | n29095;
  assign n29102 = n29094 & n29101;
  assign n29103 = n29100 & n29102;
  assign n29104 = n29098 & ~n29103;
  assign n29105 = x135 & x175;
  assign n29106 = n29104 & n29105;
  assign n29107 = n29104 | n29105;
  assign n29108 = ~n29106 & n29107;
  assign n29109 = n34316 | n29108;
  assign n29110 = n34316 & n29108;
  assign n29111 = n29109 & ~n29110;
  assign n34409 = n29049 & n34348;
  assign n34410 = n29031 & n29049;
  assign n34411 = (n34343 & n34409) | (n34343 & n34410) | (n34409 & n34410);
  assign n37687 = (n29050 & n29052) | (n29050 & n34348) | (n29052 & n34348);
  assign n37688 = n29031 & n29050;
  assign n37689 = (n29049 & n29050) | (n29049 & n37688) | (n29050 & n37688);
  assign n37149 = (n34343 & n37687) | (n34343 & n37689) | (n37687 & n37689);
  assign n29133 = ~n34411 & n37149;
  assign n34407 = n29026 & n29056;
  assign n34415 = n29133 | n34407;
  assign n34416 = n29056 | n29133;
  assign n34417 = (n34302 & n34415) | (n34302 & n34416) | (n34415 & n34416);
  assign n34418 = n29043 & n34359;
  assign n34419 = n29036 & n29043;
  assign n37150 = (n34273 & n34418) | (n34273 & n34419) | (n34418 & n34419);
  assign n37151 = (n28817 & n34418) | (n28817 & n34419) | (n34418 & n34419);
  assign n37152 = (n28790 & n37150) | (n28790 & n37151) | (n37150 & n37151);
  assign n37153 = n29036 & n29038;
  assign n37154 = (n29038 & n29043) | (n29038 & n37153) | (n29043 & n37153);
  assign n37155 = n29038 & n29043;
  assign n37156 = (n29038 & n34359) | (n29038 & n37155) | (n34359 & n37155);
  assign n37157 = (n34273 & n37154) | (n34273 & n37156) | (n37154 & n37156);
  assign n37158 = (n28817 & n37154) | (n28817 & n37156) | (n37154 & n37156);
  assign n37159 = (n28790 & n37157) | (n28790 & n37158) | (n37157 & n37158);
  assign n29138 = ~n37152 & n37159;
  assign n29140 = x142 & x169;
  assign n29142 = x143 & x168;
  assign n37160 = n29041 | n29043;
  assign n37161 = (n29041 & n34359) | (n29041 & n37160) | (n34359 & n37160);
  assign n34430 = n29142 & n37161;
  assign n37162 = n29036 | n29041;
  assign n37163 = (n29041 & n29043) | (n29041 & n37162) | (n29043 & n37162);
  assign n34431 = n29142 & n37163;
  assign n34432 = (n34274 & n34430) | (n34274 & n34431) | (n34430 & n34431);
  assign n34433 = n29142 | n37161;
  assign n34434 = n29142 | n37163;
  assign n34435 = (n34274 & n34433) | (n34274 & n34434) | (n34433 & n34434);
  assign n29145 = ~n34432 & n34435;
  assign n29146 = n29140 & n29145;
  assign n29147 = n29140 | n29145;
  assign n29148 = ~n29146 & n29147;
  assign n34436 = n29138 | n29148;
  assign n34437 = n34411 | n34436;
  assign n34438 = n29138 & n29148;
  assign n34439 = (n29148 & n34411) | (n29148 & n34438) | (n34411 & n34438);
  assign n29151 = n34437 & ~n34439;
  assign n29152 = x141 & x170;
  assign n29153 = ~n29151 & n29152;
  assign n29154 = n29151 & ~n29152;
  assign n29155 = n29153 | n29154;
  assign n29156 = n34417 | n29155;
  assign n29157 = n34417 & n29155;
  assign n29158 = n29156 & ~n29157;
  assign n34401 = ~n29026 & n29056;
  assign n34402 = ~n34302 & n34401;
  assign n34403 = n29026 & ~n29056;
  assign n34404 = (~n29056 & n34302) | (~n29056 & n34403) | (n34302 & n34403);
  assign n29126 = n34402 | n34404;
  assign n29159 = n29057 | n29126;
  assign n29160 = n29158 & n29159;
  assign n29127 = n29057 & n29126;
  assign n34405 = n28942 | n29127;
  assign n34440 = n29160 & n34405;
  assign n34441 = (n29160 & n34304) | (n29160 & n34440) | (n34304 & n34440);
  assign n29162 = n29127 | n29158;
  assign n34393 = n28942 & n29063;
  assign n34442 = n29162 | n34393;
  assign n34443 = n29063 | n29162;
  assign n34444 = (n34304 & n34442) | (n34304 & n34443) | (n34442 & n34443);
  assign n29164 = ~n34441 & n34444;
  assign n29165 = x140 & x171;
  assign n29166 = x139 & x172;
  assign n29167 = n29165 & n29166;
  assign n29168 = n29165 | n29166;
  assign n29169 = ~n29167 & n29168;
  assign n29170 = n29164 & n29169;
  assign n29171 = n29164 | n29169;
  assign n29172 = ~n29170 & n29171;
  assign n34394 = (n29063 & n34304) | (n29063 & n34393) | (n34304 & n34393);
  assign n34395 = n28942 | n29063;
  assign n34397 = n29064 & n34395;
  assign n34398 = (n29064 & n34304) | (n29064 & n34397) | (n34304 & n34397);
  assign n29122 = ~n34394 & n34398;
  assign n34399 = n29071 | n29122;
  assign n34445 = n29172 | n34399;
  assign n34446 = n29122 | n29172;
  assign n34447 = (n34338 & n34445) | (n34338 & n34446) | (n34445 & n34446);
  assign n34448 = n29172 & n34399;
  assign n34449 = n29122 & n29172;
  assign n34450 = (n34338 & n34448) | (n34338 & n34449) | (n34448 & n34449);
  assign n29175 = n34447 & ~n34450;
  assign n29176 = x138 & x173;
  assign n29177 = n29175 | n29176;
  assign n29178 = n29175 & n29176;
  assign n29179 = n29177 & ~n29178;
  assign n29114 = n34338 & n29071;
  assign n34391 = n29071 & n29072;
  assign n34392 = (n29072 & n34338) | (n29072 & n34391) | (n34338 & n34391);
  assign n29117 = ~n29114 & n34392;
  assign n34451 = n29117 & ~n29179;
  assign n34452 = (~n29179 & n34385) | (~n29179 & n34451) | (n34385 & n34451);
  assign n34453 = ~n29117 & n29179;
  assign n34454 = ~n34385 & n34453;
  assign n29182 = n34452 | n34454;
  assign n34456 = n29086 | n29182;
  assign n37164 = n29087 | n34456;
  assign n34457 = (n34322 & n37164) | (n34322 & n34456) | (n37164 & n34456);
  assign n34459 = n29086 & n29182;
  assign n37165 = (n29087 & n29182) | (n29087 & n34459) | (n29182 & n34459);
  assign n34460 = (n34322 & n37165) | (n34322 & n34459) | (n37165 & n34459);
  assign n29185 = n34457 & ~n34460;
  assign n29186 = x137 & x174;
  assign n29187 = n29185 & ~n29186;
  assign n29188 = ~n29185 & n29186;
  assign n29189 = n29187 | n29188;
  assign n34461 = n29092 & n29189;
  assign n34462 = (n29103 & n29189) | (n29103 & n34461) | (n29189 & n34461);
  assign n34463 = n29092 | n29189;
  assign n34464 = n29103 | n34463;
  assign n29192 = ~n34462 & n34464;
  assign n29193 = x136 & x175;
  assign n29194 = n29192 & n29193;
  assign n29195 = n29192 | n29193;
  assign n29196 = ~n29194 & n29195;
  assign n29197 = n29106 | n29196;
  assign n29198 = n29110 | n29197;
  assign n29199 = n28977 | n29106;
  assign n29200 = n28991 | n29199;
  assign n29112 = n29092 | n29103;
  assign n29201 = n29189 & ~n29193;
  assign n29202 = ~n29189 & n29193;
  assign n29203 = n29201 | n29202;
  assign n29204 = n29112 & n29203;
  assign n29205 = n29112 | n29203;
  assign n29206 = n29107 & n29205;
  assign n29207 = ~n29204 & n29206;
  assign n29208 = n29200 & n29207;
  assign n29209 = n29198 & ~n29208;
  assign n34465 = n29194 | n29207;
  assign n34466 = (n29194 & n29200) | (n29194 & n34465) | (n29200 & n34465);
  assign n29211 = x138 & x174;
  assign n29216 = n28963 | n29086;
  assign n34473 = n28965 | n29216;
  assign n34474 = (n28996 & n29216) | (n28996 & n34473) | (n29216 & n34473);
  assign n34486 = n29151 & n34416;
  assign n34487 = n29151 & n34415;
  assign n34488 = (n34302 & n34486) | (n34302 & n34487) | (n34486 & n34487);
  assign n34492 = n29138 & n29145;
  assign n37166 = (n29145 & n34409) | (n29145 & n34492) | (n34409 & n34492);
  assign n37167 = (n29145 & n34410) | (n29145 & n34492) | (n34410 & n34492);
  assign n37168 = (n34343 & n37166) | (n34343 & n37167) | (n37166 & n37167);
  assign n37169 = n29138 & n29140;
  assign n37170 = (n29140 & n29145) | (n29140 & n37169) | (n29145 & n37169);
  assign n37171 = (n29140 & n34409) | (n29140 & n37170) | (n34409 & n37170);
  assign n37172 = (n29140 & n34410) | (n29140 & n37170) | (n34410 & n37170);
  assign n37173 = (n34343 & n37171) | (n34343 & n37172) | (n37171 & n37172);
  assign n29237 = ~n37168 & n37173;
  assign n29239 = x142 & x170;
  assign n29241 = x143 & x169;
  assign n37174 = n29138 | n34432;
  assign n37175 = (n29145 & n34432) | (n29145 & n37174) | (n34432 & n37174);
  assign n34501 = n29241 & n37175;
  assign n37828 = n29142 & n29241;
  assign n37829 = n37161 & n37828;
  assign n37830 = n37163 & n37828;
  assign n37692 = (n34274 & n37829) | (n34274 & n37830) | (n37829 & n37830);
  assign n37177 = (n29145 & n29241) | (n29145 & n37692) | (n29241 & n37692);
  assign n37178 = (n34409 & n34501) | (n34409 & n37177) | (n34501 & n37177);
  assign n37179 = (n34410 & n34501) | (n34410 & n37177) | (n34501 & n37177);
  assign n37180 = (n34343 & n37178) | (n34343 & n37179) | (n37178 & n37179);
  assign n34504 = n29241 | n37175;
  assign n37831 = n29142 | n29241;
  assign n37832 = (n29241 & n37161) | (n29241 & n37831) | (n37161 & n37831);
  assign n37833 = (n29241 & n37163) | (n29241 & n37831) | (n37163 & n37831);
  assign n37695 = (n34274 & n37832) | (n34274 & n37833) | (n37832 & n37833);
  assign n37182 = n29145 | n37695;
  assign n37183 = (n34409 & n34504) | (n34409 & n37182) | (n34504 & n37182);
  assign n37184 = (n34410 & n34504) | (n34410 & n37182) | (n34504 & n37182);
  assign n37185 = (n34343 & n37183) | (n34343 & n37184) | (n37183 & n37184);
  assign n29244 = ~n37180 & n37185;
  assign n29245 = n29239 & n29244;
  assign n29246 = n29239 | n29244;
  assign n29247 = ~n29245 & n29246;
  assign n34507 = n29237 | n29247;
  assign n34508 = n34488 | n34507;
  assign n34509 = n29237 & n29247;
  assign n34510 = (n29247 & n34488) | (n29247 & n34509) | (n34488 & n34509);
  assign n29250 = n34508 & ~n34510;
  assign n34489 = n29151 | n34416;
  assign n34490 = n29151 | n34415;
  assign n34491 = (n34302 & n34489) | (n34302 & n34490) | (n34489 & n34490);
  assign n29231 = n29152 & n34491;
  assign n29232 = ~n34488 & n29231;
  assign n34511 = n29232 & n29250;
  assign n34512 = (n29250 & n34441) | (n29250 & n34511) | (n34441 & n34511);
  assign n34513 = n29232 | n29250;
  assign n34514 = n34441 | n34513;
  assign n29253 = ~n34512 & n34514;
  assign n29254 = x141 & x171;
  assign n29255 = n29253 & n29254;
  assign n29256 = n29253 | n29254;
  assign n29257 = ~n29255 & n29256;
  assign n29258 = x140 & x172;
  assign n29259 = n29257 & ~n29258;
  assign n29260 = ~n29257 & n29258;
  assign n29261 = n29259 | n29260;
  assign n29221 = n29164 & n29165;
  assign n29222 = n29164 | n29165;
  assign n29223 = ~n29221 & n29222;
  assign n34477 = n29223 & n34399;
  assign n34478 = n29122 & n29223;
  assign n34479 = (n34338 & n34477) | (n34338 & n34478) | (n34477 & n34478);
  assign n29262 = n29221 | n34479;
  assign n29263 = n29261 & n29262;
  assign n29264 = n29261 | n29262;
  assign n29265 = ~n29263 & n29264;
  assign n34480 = n29223 | n34399;
  assign n34481 = n29122 | n29223;
  assign n34482 = (n34338 & n34480) | (n34338 & n34481) | (n34480 & n34481);
  assign n29226 = n29166 & n34482;
  assign n29227 = ~n34479 & n29226;
  assign n34484 = n29175 | n29227;
  assign n34515 = n29265 & ~n34484;
  assign n34467 = n29117 & n29175;
  assign n34483 = n29227 | n34467;
  assign n34516 = n29265 & ~n34483;
  assign n34517 = (~n34385 & n34515) | (~n34385 & n34516) | (n34515 & n34516);
  assign n34518 = ~n29265 & n34484;
  assign n34519 = ~n29265 & n34483;
  assign n34520 = (n34385 & n34518) | (n34385 & n34519) | (n34518 & n34519);
  assign n29268 = n34517 | n34520;
  assign n29269 = x139 & x173;
  assign n29270 = n29268 & n29269;
  assign n29271 = n29268 | n29269;
  assign n29272 = ~n29270 & n29271;
  assign n34468 = (n29175 & n34385) | (n29175 & n34467) | (n34385 & n34467);
  assign n34469 = n29117 | n29175;
  assign n34471 = n29176 & n34469;
  assign n34472 = (n29176 & n34385) | (n29176 & n34471) | (n34385 & n34471);
  assign n29215 = ~n34468 & n34472;
  assign n29218 = n29085 & n29182;
  assign n34475 = n29215 | n29218;
  assign n34521 = n29272 & n34475;
  assign n34522 = n29215 & n29272;
  assign n34523 = (n34474 & n34521) | (n34474 & n34522) | (n34521 & n34522);
  assign n34524 = n29272 | n34475;
  assign n34525 = n29215 | n29272;
  assign n34526 = (n34474 & n34524) | (n34474 & n34525) | (n34524 & n34525);
  assign n29275 = ~n34523 & n34526;
  assign n29276 = n29211 & n29275;
  assign n29277 = n29211 | n29275;
  assign n29278 = ~n29276 & n29277;
  assign n29219 = n34474 & n29218;
  assign n29279 = n34457 & ~n29219;
  assign n29280 = n29186 & n29279;
  assign n29281 = n29278 | n29280;
  assign n34527 = n29281 | n34461;
  assign n34528 = n29189 | n29281;
  assign n34529 = (n29103 & n34527) | (n29103 & n34528) | (n34527 & n34528);
  assign n29285 = n29186 | n29279;
  assign n29286 = n29278 & n29285;
  assign n29283 = n29092 | n29280;
  assign n34530 = n29283 & n29286;
  assign n34531 = (n29103 & n29286) | (n29103 & n34530) | (n29286 & n34530);
  assign n29288 = n34529 & ~n34531;
  assign n29289 = x137 & x175;
  assign n29290 = n29288 & n29289;
  assign n29291 = n29288 | n29289;
  assign n29292 = ~n29290 & n29291;
  assign n29293 = n34466 & n29292;
  assign n29294 = n34466 | n29292;
  assign n29295 = ~n29293 & n29294;
  assign n29296 = n29276 | n34531;
  assign n29297 = x138 & x175;
  assign n34532 = n29265 & n34484;
  assign n34533 = n29265 & n34483;
  assign n34534 = (n34385 & n34532) | (n34385 & n34533) | (n34532 & n34533);
  assign n34535 = n29221 | n29257;
  assign n34536 = n34479 | n34535;
  assign n34537 = n29221 & n29257;
  assign n34538 = (n29257 & n34479) | (n29257 & n34537) | (n34479 & n34537);
  assign n29302 = n29258 & ~n34538;
  assign n29303 = n34536 & n29302;
  assign n29305 = x142 & x171;
  assign n29312 = x143 & x170;
  assign n34539 = n29237 & n29244;
  assign n37186 = n29312 & n37180;
  assign n37187 = (n29312 & n34539) | (n29312 & n37186) | (n34539 & n37186);
  assign n37188 = (n29244 & n29312) | (n29244 & n37186) | (n29312 & n37186);
  assign n34553 = (n34488 & n37187) | (n34488 & n37188) | (n37187 & n37188);
  assign n37189 = n29312 | n37180;
  assign n37190 = n34539 | n37189;
  assign n37191 = n29244 | n37189;
  assign n34556 = (n34488 & n37190) | (n34488 & n37191) | (n37190 & n37191);
  assign n29315 = ~n34553 & n34556;
  assign n34540 = (n29244 & n34488) | (n29244 & n34539) | (n34488 & n34539);
  assign n34541 = n29237 | n29244;
  assign n34543 = n29239 & n34541;
  assign n34544 = (n29239 & n34488) | (n29239 & n34543) | (n34488 & n34543);
  assign n29309 = ~n34540 & n34544;
  assign n37192 = n29309 & n29315;
  assign n37193 = (n29315 & n34511) | (n29315 & n37192) | (n34511 & n37192);
  assign n34546 = n29250 | n29309;
  assign n34558 = n29315 & n34546;
  assign n34559 = (n34441 & n37193) | (n34441 & n34558) | (n37193 & n34558);
  assign n37194 = n29309 | n29315;
  assign n37195 = n34511 | n37194;
  assign n34561 = n29315 | n34546;
  assign n34562 = (n34441 & n37195) | (n34441 & n34561) | (n37195 & n34561);
  assign n29318 = ~n34559 & n34562;
  assign n29319 = n29305 & n29318;
  assign n29320 = n29305 | n29318;
  assign n29321 = ~n29319 & n29320;
  assign n34564 = n29122 | n29221;
  assign n29323 = n29250 | n29254;
  assign n29324 = n29250 & n29254;
  assign n29325 = n29323 & ~n29324;
  assign n34566 = n29232 | n29325;
  assign n34567 = n34441 | n34566;
  assign n34568 = n29232 & n29325;
  assign n34569 = (n29325 & n34441) | (n29325 & n34568) | (n34441 & n34568);
  assign n34570 = n34567 & ~n34569;
  assign n34571 = n29222 & n34570;
  assign n34572 = n34564 & n34571;
  assign n34563 = n29221 | n34399;
  assign n34573 = n34563 & n34571;
  assign n34574 = (n34338 & n34572) | (n34338 & n34573) | (n34572 & n34573);
  assign n34575 = n29255 & n29321;
  assign n34576 = (n29321 & n34574) | (n29321 & n34575) | (n34574 & n34575);
  assign n34577 = n29255 | n29321;
  assign n34578 = n34574 | n34577;
  assign n29334 = ~n34576 & n34578;
  assign n29335 = x141 & x172;
  assign n29336 = n29334 & n29335;
  assign n29337 = n29334 | n29335;
  assign n29338 = ~n29336 & n29337;
  assign n34579 = ~n29303 & n29338;
  assign n34580 = ~n34534 & n34579;
  assign n34581 = n29303 & ~n29338;
  assign n34582 = (~n29338 & n34534) | (~n29338 & n34581) | (n34534 & n34581);
  assign n29341 = n34580 | n34582;
  assign n29342 = x140 & x173;
  assign n29343 = n29341 & n29342;
  assign n29344 = n29341 | n29342;
  assign n29345 = ~n29343 & n29344;
  assign n34583 = n29270 & n29345;
  assign n34584 = (n29345 & n34523) | (n29345 & n34583) | (n34523 & n34583);
  assign n34585 = n29270 | n29345;
  assign n34586 = n34523 | n34585;
  assign n29348 = ~n34584 & n34586;
  assign n29349 = x139 & x174;
  assign n29350 = n29348 & n29349;
  assign n29351 = n29348 | n29349;
  assign n29352 = ~n29350 & n29351;
  assign n29353 = ~n29297 & n29352;
  assign n29354 = n29297 & ~n29352;
  assign n29355 = n29353 | n29354;
  assign n29356 = n29296 | n29355;
  assign n29357 = n29296 & n29355;
  assign n29358 = n29356 & ~n29357;
  assign n29359 = n29290 | n29358;
  assign n34587 = n29292 | n29359;
  assign n34588 = (n29359 & n34466) | (n29359 & n34587) | (n34466 & n34587);
  assign n29361 = n29194 | n29290;
  assign n34589 = n29207 | n29361;
  assign n34590 = (n29200 & n29361) | (n29200 & n34589) | (n29361 & n34589);
  assign n29363 = n29291 & n29358;
  assign n29364 = n34590 & n29363;
  assign n29365 = n34588 & ~n29364;
  assign n34602 = n29303 & n29338;
  assign n34603 = (n29338 & n34534) | (n29338 & n34602) | (n34534 & n34602);
  assign n29375 = x142 & x172;
  assign n29377 = x143 & x171;
  assign n37697 = n29312 & n29377;
  assign n37834 = n37180 & n37697;
  assign n37698 = (n34539 & n37834) | (n34539 & n37697) | (n37834 & n37697);
  assign n37203 = n29377 & n37188;
  assign n37204 = (n34488 & n37698) | (n34488 & n37203) | (n37698 & n37203);
  assign n37699 = (n29315 & n29377) | (n29315 & n37204) | (n29377 & n37204);
  assign n37904 = n29377 & n37697;
  assign n37922 = n37180 & n37904;
  assign n37905 = (n34539 & n37922) | (n34539 & n37904) | (n37922 & n37904);
  assign n37837 = (n34488 & n37203) | (n34488 & n37905) | (n37203 & n37905);
  assign n37701 = (n34546 & n37699) | (n34546 & n37837) | (n37699 & n37837);
  assign n37206 = (n29377 & n37193) | (n29377 & n37204) | (n37193 & n37204);
  assign n37207 = (n34441 & n37701) | (n34441 & n37206) | (n37701 & n37206);
  assign n37703 = n29312 | n29377;
  assign n37838 = (n29377 & n37180) | (n29377 & n37703) | (n37180 & n37703);
  assign n37704 = (n34539 & n37838) | (n34539 & n37703) | (n37838 & n37703);
  assign n37209 = n29377 | n37188;
  assign n37210 = (n34488 & n37704) | (n34488 & n37209) | (n37704 & n37209);
  assign n37705 = n29315 | n37210;
  assign n37706 = (n34546 & n37210) | (n34546 & n37705) | (n37210 & n37705);
  assign n37212 = n37193 | n37210;
  assign n37213 = (n34441 & n37706) | (n34441 & n37212) | (n37706 & n37212);
  assign n29380 = ~n37207 & n37213;
  assign n29381 = n29375 & n29380;
  assign n29382 = n29375 | n29380;
  assign n29383 = ~n29381 & n29382;
  assign n34608 = n29319 | n29383;
  assign n34609 = n34576 | n34608;
  assign n34610 = n29319 & n29383;
  assign n34611 = (n29383 & n34576) | (n29383 & n34610) | (n34576 & n34610);
  assign n29386 = n34609 & ~n34611;
  assign n29387 = x141 & x173;
  assign n29388 = ~n29386 & n29387;
  assign n29389 = n29386 & ~n29387;
  assign n29390 = n29388 | n29389;
  assign n34612 = n29336 | n29390;
  assign n34613 = n34603 | n34612;
  assign n34614 = n29336 & n29390;
  assign n34615 = (n29390 & n34603) | (n29390 & n34614) | (n34603 & n34614);
  assign n29393 = n34613 & ~n34615;
  assign n29394 = n29343 | n29393;
  assign n29395 = n34584 | n29394;
  assign n29400 = x140 & x174;
  assign n29397 = n29344 & n29393;
  assign n34616 = n29270 | n29343;
  assign n34618 = n29397 & n34616;
  assign n34619 = (n29397 & n34523) | (n29397 & n34618) | (n34523 & n34618);
  assign n34620 = n29400 & ~n34619;
  assign n34621 = n29395 & n34620;
  assign n34622 = ~n29400 & n34619;
  assign n34623 = (n29395 & n29400) | (n29395 & ~n34622) | (n29400 & ~n34622);
  assign n29403 = ~n34621 & n34623;
  assign n34600 = n29350 | n29352;
  assign n37214 = n29403 & n34600;
  assign n37200 = n29276 | n29350;
  assign n37201 = (n29350 & n29352) | (n29350 & n37200) | (n29352 & n37200);
  assign n37215 = n29403 & n37201;
  assign n37216 = (n34531 & n37214) | (n34531 & n37215) | (n37214 & n37215);
  assign n37217 = n29403 | n34600;
  assign n37218 = n29403 | n37201;
  assign n37219 = (n34531 & n37217) | (n34531 & n37218) | (n37217 & n37218);
  assign n29406 = ~n37216 & n37219;
  assign n29407 = x139 & x175;
  assign n29408 = n29406 & n29407;
  assign n29409 = n29406 | n29407;
  assign n29410 = ~n29408 & n29409;
  assign n34591 = n29276 & n29352;
  assign n34592 = (n29352 & n34531) | (n29352 & n34591) | (n34531 & n34591);
  assign n37707 = n29211 & n29297;
  assign n37708 = n29275 & n37707;
  assign n37197 = (n29297 & n29352) | (n29297 & n37708) | (n29352 & n37708);
  assign n34596 = (n29297 & n34531) | (n29297 & n37197) | (n34531 & n37197);
  assign n29369 = ~n34592 & n34596;
  assign n37198 = n29291 | n29369;
  assign n37199 = (n29358 & n29369) | (n29358 & n37198) | (n29369 & n37198);
  assign n37220 = n29410 & n37199;
  assign n37221 = n29369 & n29410;
  assign n37222 = (n34590 & n37220) | (n34590 & n37221) | (n37220 & n37221);
  assign n37223 = n29410 | n37199;
  assign n37224 = n29369 | n29410;
  assign n37225 = (n34590 & n37223) | (n34590 & n37224) | (n37223 & n37224);
  assign n29413 = ~n37222 & n37225;
  assign n34598 = (n29369 & n34590) | (n29369 & n37199) | (n34590 & n37199);
  assign n29422 = x143 & x172;
  assign n37226 = n29380 | n37207;
  assign n37227 = (n29319 & n37207) | (n29319 & n37226) | (n37207 & n37226);
  assign n34635 = n29422 & n37227;
  assign n37228 = n29422 & n37207;
  assign n37229 = (n29380 & n29422) | (n29380 & n37228) | (n29422 & n37228);
  assign n34637 = (n34576 & n34635) | (n34576 & n37229) | (n34635 & n37229);
  assign n34638 = n29422 | n37227;
  assign n37230 = n29422 | n37207;
  assign n37231 = n29380 | n37230;
  assign n34640 = (n34576 & n34638) | (n34576 & n37231) | (n34638 & n37231);
  assign n29425 = ~n34637 & n34640;
  assign n34626 = n29319 & n29380;
  assign n34627 = (n29380 & n34576) | (n29380 & n34626) | (n34576 & n34626);
  assign n34628 = n29319 | n29380;
  assign n34629 = n34576 | n34628;
  assign n29418 = ~n34627 & n34629;
  assign n29426 = n29375 | n29418;
  assign n29427 = n29425 & n29426;
  assign n29419 = n29375 & n29418;
  assign n34630 = n29336 | n29419;
  assign n34641 = n29427 & n34630;
  assign n34642 = (n29427 & n34603) | (n29427 & n34641) | (n34603 & n34641);
  assign n29430 = n29419 | n29425;
  assign n34643 = n29336 & n29386;
  assign n34645 = n29430 | n34643;
  assign n37232 = n29386 | n29425;
  assign n37233 = n29419 | n37232;
  assign n34647 = (n34603 & n34645) | (n34603 & n37233) | (n34645 & n37233);
  assign n29432 = ~n34642 & n34647;
  assign n29433 = x142 & x173;
  assign n29434 = n29432 & n29433;
  assign n29435 = n29432 | n29433;
  assign n29436 = ~n29434 & n29435;
  assign n34648 = n29336 | n29386;
  assign n34649 = n34603 | n34648;
  assign n34650 = n29387 & ~n34643;
  assign n34651 = (n29388 & ~n34603) | (n29388 & n34650) | (~n34603 & n34650);
  assign n29439 = n34649 & n34651;
  assign n34652 = n29436 & n29439;
  assign n34653 = (n29436 & n34619) | (n29436 & n34652) | (n34619 & n34652);
  assign n34654 = n29436 | n29439;
  assign n34655 = n34619 | n34654;
  assign n29443 = ~n34653 & n34655;
  assign n29444 = x141 & x174;
  assign n29445 = n29443 & n29444;
  assign n29446 = n29443 | n29444;
  assign n29447 = ~n29445 & n29446;
  assign n29448 = n34623 & n29447;
  assign n34601 = (n34531 & n37201) | (n34531 & n34600) | (n37201 & n34600);
  assign n37234 = n34621 & n34623;
  assign n37235 = n29447 & n37234;
  assign n34657 = (n29448 & n34601) | (n29448 & n37235) | (n34601 & n37235);
  assign n29450 = n34621 | n29447;
  assign n37236 = n29403 | n34621;
  assign n37237 = n29447 | n37236;
  assign n34659 = (n29450 & n34601) | (n29450 & n37237) | (n34601 & n37237);
  assign n29452 = ~n34657 & n34659;
  assign n29453 = x140 & x175;
  assign n29454 = n29452 & n29453;
  assign n29455 = n29452 | n29453;
  assign n29456 = ~n29454 & n29455;
  assign n34624 = n29408 | n29410;
  assign n37238 = n29456 | n34624;
  assign n37239 = n29408 | n29456;
  assign n37240 = (n34598 & n37238) | (n34598 & n37239) | (n37238 & n37239);
  assign n37241 = n29456 & n34624;
  assign n37242 = n29408 & n29456;
  assign n37243 = (n34598 & n37241) | (n34598 & n37242) | (n37241 & n37242);
  assign n29459 = n37240 & ~n37243;
  assign n29463 = x143 & x173;
  assign n37709 = n29422 & n29463;
  assign n37710 = n37227 & n37709;
  assign n37245 = n29463 & n37229;
  assign n37246 = (n34576 & n37710) | (n34576 & n37245) | (n37710 & n37245);
  assign n34663 = (n29463 & n34642) | (n29463 & n37246) | (n34642 & n37246);
  assign n37711 = n29422 | n29463;
  assign n37712 = (n29463 & n37227) | (n29463 & n37711) | (n37227 & n37711);
  assign n37248 = n29463 | n37229;
  assign n37249 = (n34576 & n37712) | (n34576 & n37248) | (n37712 & n37248);
  assign n34665 = n34642 | n37249;
  assign n29466 = ~n34663 & n34665;
  assign n29469 = n29434 | n29466;
  assign n29470 = n34653 | n29469;
  assign n29472 = x142 & x174;
  assign n29467 = n29435 & n29466;
  assign n34660 = n29434 | n29439;
  assign n34666 = n29467 & n34660;
  assign n34667 = (n29467 & n34619) | (n29467 & n34666) | (n34619 & n34666);
  assign n34668 = n29472 & ~n34667;
  assign n34669 = n29470 & n34668;
  assign n34670 = ~n29472 & n34667;
  assign n34671 = (n29470 & n29472) | (n29470 & ~n34670) | (n29472 & ~n34670);
  assign n29475 = ~n34669 & n34671;
  assign n29476 = x141 & x175;
  assign n29477 = n29475 & ~n29476;
  assign n29478 = ~n29475 & n29476;
  assign n29479 = n29477 | n29478;
  assign n34672 = n29445 & n29479;
  assign n34673 = (n29479 & n34657) | (n29479 & n34672) | (n34657 & n34672);
  assign n34674 = n29445 | n29479;
  assign n34675 = n34657 | n34674;
  assign n29482 = ~n34673 & n34675;
  assign n29483 = n29454 | n29482;
  assign n34625 = (n29408 & n34598) | (n29408 & n34624) | (n34598 & n34624);
  assign n34676 = n29456 | n29483;
  assign n34677 = (n29483 & n34625) | (n29483 & n34676) | (n34625 & n34676);
  assign n29485 = n29408 | n29454;
  assign n34678 = n29410 | n29485;
  assign n34679 = (n29485 & n34598) | (n29485 & n34678) | (n34598 & n34678);
  assign n29487 = n29455 & n29482;
  assign n29488 = n34679 & n29487;
  assign n29489 = n34677 & ~n29488;
  assign n29497 = x143 & x174;
  assign n37839 = n29497 & n37709;
  assign n37840 = n37227 & n37839;
  assign n37251 = n29463 & n29497;
  assign n37841 = n37229 & n37251;
  assign n37715 = (n34576 & n37840) | (n34576 & n37841) | (n37840 & n37841);
  assign n37252 = (n34642 & n37715) | (n34642 & n37251) | (n37715 & n37251);
  assign n34691 = (n29497 & n34667) | (n29497 & n37252) | (n34667 & n37252);
  assign n37842 = n29497 | n37709;
  assign n37843 = (n29497 & n37227) | (n29497 & n37842) | (n37227 & n37842);
  assign n37254 = n29463 | n29497;
  assign n37844 = (n29497 & n37229) | (n29497 & n37254) | (n37229 & n37254);
  assign n37718 = (n34576 & n37843) | (n34576 & n37844) | (n37843 & n37844);
  assign n37255 = (n34642 & n37718) | (n34642 & n37254) | (n37718 & n37254);
  assign n34693 = n34667 | n37255;
  assign n29500 = ~n34691 & n34693;
  assign n29503 = n34669 | n29500;
  assign n34680 = n29445 & n29475;
  assign n34696 = n29503 | n34680;
  assign n34697 = n29475 | n29503;
  assign n34698 = (n34657 & n34696) | (n34657 & n34697) | (n34696 & n34697);
  assign n29506 = x142 & x175;
  assign n29501 = n34671 & n29500;
  assign n34688 = n29445 | n34669;
  assign n34694 = n29501 & n34688;
  assign n37256 = (n29501 & n34694) | (n29501 & n37235) | (n34694 & n37235);
  assign n37257 = (n29448 & n29501) | (n29448 & n34694) | (n29501 & n34694);
  assign n37258 = (n34601 & n37256) | (n34601 & n37257) | (n37256 & n37257);
  assign n37259 = n29506 & ~n37258;
  assign n37260 = n34698 & n37259;
  assign n37261 = ~n29506 & n37258;
  assign n37262 = (n29506 & n34698) | (n29506 & ~n37261) | (n34698 & ~n37261);
  assign n29509 = ~n37260 & n37262;
  assign n37263 = (n29475 & n34680) | (n29475 & n37235) | (n34680 & n37235);
  assign n37264 = (n29448 & n29475) | (n29448 & n34680) | (n29475 & n34680);
  assign n37265 = (n34601 & n37263) | (n34601 & n37264) | (n37263 & n37264);
  assign n37719 = n29444 & n29476;
  assign n37720 = n29443 & n37719;
  assign n37267 = (n29475 & n29476) | (n29475 & n37720) | (n29476 & n37720);
  assign n37268 = (n29476 & n37235) | (n29476 & n37267) | (n37235 & n37267);
  assign n37269 = (n29448 & n29476) | (n29448 & n37267) | (n29476 & n37267);
  assign n37270 = (n34601 & n37268) | (n34601 & n37269) | (n37268 & n37269);
  assign n29493 = ~n37265 & n37270;
  assign n34686 = n29487 | n29493;
  assign n34699 = n29509 & n34686;
  assign n34700 = n29493 & n29509;
  assign n34701 = (n34679 & n34699) | (n34679 & n34700) | (n34699 & n34700);
  assign n34702 = n29509 | n34686;
  assign n34703 = n29493 | n29509;
  assign n34704 = (n34679 & n34702) | (n34679 & n34703) | (n34702 & n34703);
  assign n29512 = ~n34701 & n34704;
  assign n29515 = x143 & x175;
  assign n37722 = n29497 & n29515;
  assign n37933 = n37709 & n37722;
  assign n37924 = n37227 & n37933;
  assign n37846 = n29515 & n37251;
  assign n37925 = n37229 & n37846;
  assign n37908 = (n34576 & n37924) | (n34576 & n37925) | (n37924 & n37925);
  assign n37847 = (n34642 & n37908) | (n34642 & n37846) | (n37908 & n37846);
  assign n37723 = (n34667 & n37847) | (n34667 & n37722) | (n37847 & n37722);
  assign n37274 = (n29515 & n34694) | (n29515 & n37723) | (n34694 & n37723);
  assign n37275 = (n29501 & n29515) | (n29501 & n37723) | (n29515 & n37723);
  assign n34713 = (n34657 & n37274) | (n34657 & n37275) | (n37274 & n37275);
  assign n37725 = n29497 | n29515;
  assign n37934 = (n29515 & n37709) | (n29515 & n37725) | (n37709 & n37725);
  assign n37927 = (n29515 & n37227) | (n29515 & n37934) | (n37227 & n37934);
  assign n37849 = n29515 | n37251;
  assign n37928 = (n29515 & n37229) | (n29515 & n37849) | (n37229 & n37849);
  assign n37911 = (n34576 & n37927) | (n34576 & n37928) | (n37927 & n37928);
  assign n37850 = (n34642 & n37911) | (n34642 & n37849) | (n37911 & n37849);
  assign n37726 = (n34667 & n37850) | (n34667 & n37725) | (n37850 & n37725);
  assign n37277 = n34694 | n37726;
  assign n37278 = n29501 | n37726;
  assign n34716 = (n34657 & n37277) | (n34657 & n37278) | (n37277 & n37278);
  assign n29518 = ~n34713 & n34716;
  assign n29519 = n37262 & n29518;
  assign n37271 = n29493 | n37260;
  assign n37272 = n29487 | n37271;
  assign n37279 = n29519 & n37272;
  assign n34706 = n29493 | n37260;
  assign n37280 = n29519 & n34706;
  assign n37281 = (n34679 & n37279) | (n34679 & n37280) | (n37279 & n37280);
  assign n29521 = n37260 | n29518;
  assign n29522 = n34701 | n29521;
  assign n29523 = ~n37281 & n29522;
  assign n34717 = n29519 | n34713;
  assign n37282 = (n34713 & n34717) | (n34713 & n37272) | (n34717 & n37272);
  assign n37283 = (n34706 & n34713) | (n34706 & n34717) | (n34713 & n34717);
  assign n37284 = (n34679 & n37282) | (n34679 & n37283) | (n37282 & n37283);
  assign y0 = n17;
  assign y1 = n22;
  assign y2 = n34;
  assign y3 = n54;
  assign y4 = n82;
  assign y5 = n118;
  assign y6 = n162;
  assign y7 = n214;
  assign y8 = n266;
  assign y9 = n314;
  assign y10 = n355;
  assign y11 = n388;
  assign y12 = n413;
  assign y13 = n430;
  assign y14 = n439;
  assign y15 = n723;
  assign y16 = n827;
  assign y17 = n832;
  assign y18 = n844;
  assign y19 = n864;
  assign y20 = n892;
  assign y21 = n928;
  assign y22 = n972;
  assign y23 = n1024;
  assign y24 = n1084;
  assign y25 = n1152;
  assign y26 = n1228;
  assign y27 = n1312;
  assign y28 = n1404;
  assign y29 = n1504;
  assign y30 = n1612;
  assign y31 = n1728;
  assign y32 = n1844;
  assign y33 = n1956;
  assign y34 = n2061;
  assign y35 = n2158;
  assign y36 = n2247;
  assign y37 = n2328;
  assign y38 = n2401;
  assign y39 = n2466;
  assign y40 = n2523;
  assign y41 = n2572;
  assign y42 = n2613;
  assign y43 = n2646;
  assign y44 = n2671;
  assign y45 = n2688;
  assign y46 = n2697;
  assign y47 = n3896;
  assign y48 = n4203;
  assign y49 = n4208;
  assign y50 = n4220;
  assign y51 = n4240;
  assign y52 = n4268;
  assign y53 = n4304;
  assign y54 = n4348;
  assign y55 = n4400;
  assign y56 = n4460;
  assign y57 = n4528;
  assign y58 = n4604;
  assign y59 = n4688;
  assign y60 = n4780;
  assign y61 = n4880;
  assign y62 = n4988;
  assign y63 = n5104;
  assign y64 = n5228;
  assign y65 = n5360;
  assign y66 = n5500;
  assign y67 = n5648;
  assign y68 = n5804;
  assign y69 = n5968;
  assign y70 = n6140;
  assign y71 = n6320;
  assign y72 = n6508;
  assign y73 = n6704;
  assign y74 = n6908;
  assign y75 = n7120;
  assign y76 = n7340;
  assign y77 = n7568;
  assign y78 = n7804;
  assign y79 = n8048;
  assign y80 = n8292;
  assign y81 = n8532;
  assign y82 = n8765;
  assign y83 = n8990;
  assign y84 = n9207;
  assign y85 = n9416;
  assign y86 = n9617;
  assign y87 = n9810;
  assign y88 = n9995;
  assign y89 = n10172;
  assign y90 = n10341;
  assign y91 = n10502;
  assign y92 = n10655;
  assign y93 = n10800;
  assign y94 = n10937;
  assign y95 = n11066;
  assign y96 = n11187;
  assign y97 = n11300;
  assign y98 = n11405;
  assign y99 = n11502;
  assign y100 = n11591;
  assign y101 = n11672;
  assign y102 = n11745;
  assign y103 = n11810;
  assign y104 = n11867;
  assign y105 = n11916;
  assign y106 = n11957;
  assign y107 = n11990;
  assign y108 = n12015;
  assign y109 = n12032;
  assign y110 = n12041;
  assign y111 = n17673;
  assign y112 = n18337;
  assign y113 = n18342;
  assign y114 = n18354;
  assign y115 = n18375;
  assign y116 = n18406;
  assign y117 = n18443;
  assign y118 = n18501;
  assign y119 = n18555;
  assign y120 = n18636;
  assign y121 = n18724;
  assign y122 = n18822;
  assign y123 = n18943;
  assign y124 = n19056;
  assign y125 = n19182;
  assign y126 = n19324;
  assign y127 = n19476;
  assign y128 = n19640;
  assign y129 = n19815;
  assign y130 = n20011;
  assign y131 = n20209;
  assign y132 = n20411;
  assign y133 = n20640;
  assign y134 = n20885;
  assign y135 = n21142;
  assign y136 = n21404;
  assign y137 = n21705;
  assign y138 = n22005;
  assign y139 = n22327;
  assign y140 = n22642;
  assign y141 = n22983;
  assign y142 = n23325;
  assign y143 = n23674;
  assign y144 = n24028;
  assign y145 = n24382;
  assign y146 = n24708;
  assign y147 = n25030;
  assign y148 = n25331;
  assign y149 = n25641;
  assign y150 = n25945;
  assign y151 = n26275;
  assign y152 = n26506;
  assign y153 = n26792;
  assign y154 = n27047;
  assign y155 = n27273;
  assign y156 = n27487;
  assign y157 = n27681;
  assign y158 = n27878;
  assign y159 = n28090;
  assign y160 = n28291;
  assign y161 = n28453;
  assign y162 = n28605;
  assign y163 = n28754;
  assign y164 = n28882;
  assign y165 = n28992;
  assign y166 = n29111;
  assign y167 = n29209;
  assign y168 = n29295;
  assign y169 = n29365;
  assign y170 = n29413;
  assign y171 = n29459;
  assign y172 = n29489;
  assign y173 = n29512;
  assign y174 = n29523;
  assign y175 = n37284;
endmodule

