module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159, y160, y161, y162, y163, y164, y165, y166, y167, y168, y169, y170, y171, y172, y173, y174, y175, y176, y177, y178, y179, y180, y181, y182, y183, y184, y185, y186, y187, y188, y189, y190, y191, y192, y193, y194, y195, y196, y197, y198, y199, y200, y201, y202, y203, y204, y205, y206, y207, y208, y209, y210, y211, y212, y213, y214, y215, y216, y217, y218, y219, y220, y221, y222, y223, y224, y225, y226, y227, y228, y229, y230, y231, y232, y233, y234, y235, y236, y237, y238, y239);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159, y160, y161, y162, y163, y164, y165, y166, y167, y168, y169, y170, y171, y172, y173, y174, y175, y176, y177, y178, y179, y180, y181, y182, y183, y184, y185, y186, y187, y188, y189, y190, y191, y192, y193, y194, y195, y196, y197, y198, y199, y200, y201, y202, y203, y204, y205, y206, y207, y208, y209, y210, y211, y212, y213, y214, y215, y216, y217, y218, y219, y220, y221, y222, y223, y224, y225, y226, y227, y228, y229, y230, y231, y232, y233, y234, y235, y236, y237, y238, y239;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246, n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254, n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318, n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326, n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386, n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534, n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587, n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598, n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606, n42607, n42608, n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626, n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794, n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817, n42818, n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841, n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866, n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890, n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913, n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938, n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982, n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019, n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043, n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091, n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099, n43100, n43101, n43102, n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114, n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129, n43130, n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178, n43179, n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187, n43188, n43189, n43190, n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201, n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270, n43271, n43272, n43273, n43274, n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282, n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307, n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345, n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379, n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417, n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451, n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489, n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523, n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534, n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550, n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561, n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595, n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606, n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667, n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678, n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705, n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739, n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763, n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777, n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811, n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849, n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883, n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921, n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955, n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971, n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979, n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993, n43994, n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002, n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027, n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042, n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051, n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062, n44063, n44064, n44065, n44066, n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099, n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44136, n44137, n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146, n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44209, n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258, n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267, n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282, n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330, n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339, n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347, n44348, n44349, n44350, n44351, n44352, n44353, n44354, n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387, n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411, n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419, n44420, n44421, n44422, n44423, n44424, n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459, n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496, n44497, n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546, n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555, n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569, n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627, n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641, n44642, n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650, n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675, n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690, n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699, n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710, n44711, n44712, n44713, n44714, n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747, n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762, n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771, n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779, n44780, n44781, n44782, n44783, n44784, n44785, n44786, n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819, n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854, n44855, n44856, n44857, n44858, n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891, n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926, n44927, n44928, n44929, n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963, n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001, n45002, n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010, n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035, n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050, n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067, n45068, n45069, n45070, n45071, n45072, n45073, n45074, n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107, n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122, n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131, n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139, n45140, n45141, n45142, n45143, n45144, n45145, n45146, n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154, n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179, n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194, n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218, n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250, n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258, n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266, n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274, n45275, n45276, n45277, n45278, n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286, n45287, n45288, n45289, n45290, n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306, n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338, n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352, n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360, n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378, n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386, n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395, n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418, n45419, n45420, n45421, n45422, n45423, n45424, n45425, n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433, n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442, n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466, n45467, n45468, n45469, n45470, n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482, n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45496, n45497, n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505, n45506, n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514, n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522, n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530, n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538, n45539, n45540, n45541, n45542, n45543, n45544, n45545, n45546, n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562, n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570, n45571, n45572, n45573, n45574, n45575, n45576, n45577, n45578, n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586, n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594, n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602, n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610, n45611, n45612, n45613, n45614, n45615, n45616, n45617, n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626, n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638, n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648, n45649, n45650, n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674, n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682, n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720, n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746, n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754, n45755, n45756, n45757, n45758, n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782, n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790, n45791, n45792, n45793, n45794, n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802, n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810, n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832, n45833, n45834, n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842, n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864, n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890, n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899, n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954, n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962, n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972, n45973, n45974, n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026, n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043, n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058, n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078, n46079, n46080, n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106, n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150, n46151, n46152, n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202, n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211, n46212, n46213, n46214, n46215, n46216, n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224, n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274, n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296, n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322, n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331, n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363, n46364, n46365, n46366, n46367, n46368, n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403, n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430, n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438, n46439, n46440, n46441, n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466, n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474, n46475, n46476, n46477, n46478, n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502, n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510, n46511, n46512, n46513, n46514, n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538, n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553, n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562, n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570, n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578, n46579, n46580, n46581, n46582, n46583, n46584, n46585, n46586, n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610, n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626, n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634, n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642, n46643, n46644, n46645, n46646, n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654, n46655, n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682, n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706, n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714, n46715, n46716, n46717, n46718, n46719, n46720, n46721, n46722, n46723, n46724, n46725, n46726, n46727, n46728, n46729, n46730, n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754, n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762, n46763, n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778, n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786, n46787, n46788, n46789, n46790, n46791, n46792, n46793, n46794, n46795, n46796, n46797, n46798, n46799, n46800, n46801, n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810, n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826, n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834, n46835, n46836, n46837, n46838, n46839, n46840, n46841, n46842, n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850, n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858, n46859, n46860, n46861, n46862, n46863, n46864, n46865, n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873, n46874, n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882, n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890, n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898, n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906, n46907, n46908, n46909, n46910, n46911, n46912, n46913, n46914, n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922, n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930, n46931, n46932, n46933, n46934, n46935, n46936, n46937, n46938, n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946, n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954, n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962, n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970, n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978, n46979, n46980, n46981, n46982, n46983, n46984, n46985, n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994, n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002, n47003, n47004, n47005, n47006, n47007, n47008, n47009, n47010, n47011, n47012, n47013, n47014, n47015, n47016, n47017, n47018, n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026, n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042, n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057, n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066, n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074, n47075, n47076, n47077, n47078, n47079, n47080, n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089, n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138, n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146, n47147, n47148, n47149, n47150, n47151, n47152, n47153, n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161, n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186, n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201, n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210, n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218, n47219, n47220, n47221, n47222, n47223, n47224, n47225, n47226, n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47234, n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250, n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258, n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266, n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306, n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322, n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345, n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354, n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377, n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402, n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410, n47411, n47412, n47413, n47414, n47415, n47416, n47417, n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426, n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434, n47435, n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443, n47444, n47445, n47446, n47447, n47448, n47449, n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466, n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498, n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522, n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530, n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538, n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546, n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554, n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570, n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578, n47579, n47580, n47581, n47582, n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590, n47591, n47592, n47593, n47594, n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610, n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618, n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642, n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650, n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659, n47660, n47661, n47662, n47663, n47664, n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690, n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699, n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714, n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722, n47723, n47724, n47725, n47726, n47727, n47728, n47729, n47730, n47731, n47732, n47733, n47734, n47735, n47736, n47737, n47738, n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746, n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771, n47772, n47773, n47774, n47775, n47776, n47777, n47778, n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786, n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794, n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802, n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810, n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818, n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826, n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834, n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842, n47843, n47844, n47845, n47846, n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882, n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890, n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898, n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914, n47915, n47916, n47917, n47918, n47919, n47920, n47921, n47922, n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930, n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938, n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946, n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954, n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962, n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970, n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978, n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987, n47988, n47989, n47990, n47991, n47992, n47993, n47994, n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002, n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026, n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058, n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48066, n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074, n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082, n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090, n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098, n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106, n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114, n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122, n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130, n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162, n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170, n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178, n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186, n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194, n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202, n48203, n48204, n48205, n48206, n48207, n48208, n48209, n48210, n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218, n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226, n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234, n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242, n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250, n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258, n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266, n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274, n48275, n48276, n48277, n48278, n48279, n48280, n48281, n48282, n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290, n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298, n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306, n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322, n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330, n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338, n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346, n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354, n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362, n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370, n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378, n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386, n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394, n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410, n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418, n48419, n48420, n48421, n48422, n48423, n48424, n48425, n48426, n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434, n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442, n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450, n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458, n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466, n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474, n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482, n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490, n48491, n48492, n48493, n48494, n48495, n48496, n48497, n48498, n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506, n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514, n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530, n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554, n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570, n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578, n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602, n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610, n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618, n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626, n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634, n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642, n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650, n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658, n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666, n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674, n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682, n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690, n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698, n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706, n48707, n48708, n48709, n48710, n48711, n48712, n48713, n48714, n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722, n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746, n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754, n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762, n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770, n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778, n48779, n48780, n48781, n48782, n48783, n48784, n48785, n48786, n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794, n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818, n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826, n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834, n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842, n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850, n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858, n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866, n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882, n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890, n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898, n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906, n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914, n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922, n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930, n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938, n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946, n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962, n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970, n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978, n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986, n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994, n48995, n48996, n48997, n48998, n48999, n49000, n49001, n49002, n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010, n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018, n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026, n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042, n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050, n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058, n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066, n49067, n49068, n49069, n49070, n49071, n49072, n49073, n49074, n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082, n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090, n49091, n49092, n49093, n49094, n49095, n49096, n49097, n49098, n49099, n49100, n49101, n49102, n49103, n49104, n49105, n49106, n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114, n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122, n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130, n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138, n49139, n49140, n49141, n49142, n49143, n49144, n49145, n49146, n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154, n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168, n49169, n49170, n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178, n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186, n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194, n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202, n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210, n49211, n49212, n49213, n49214, n49215, n49216, n49217, n49218, n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226, n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234, n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242, n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250, n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258, n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266, n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274, n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282, n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290, n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298, n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306, n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314, n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322, n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330, n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338, n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346, n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360, n49361, n49362, n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370, n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378, n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386, n49387, n49388, n49389, n49390, n49391, n49392, n49393, n49394, n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402, n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410, n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418, n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442, n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458, n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466, n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474, n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482, n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490, n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498, n49499, n49500, n49501, n49502, n49503, n49504, n49505, n49506, n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514, n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522, n49523, n49524, n49525, n49526, n49527, n49528, n49529, n49530, n49531, n49532, n49533, n49534, n49535, n49536, n49537, n49538, n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554, n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562, n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570, n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578, n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586, n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594, n49595, n49596, n49597, n49598, n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606, n49607, n49608, n49609, n49610, n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618, n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626, n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634, n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642, n49643, n49644, n49645, n49646, n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658, n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666, n49667, n49668, n49669, n49670, n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678, n49679, n49680, n49681, n49682, n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698, n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706, n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714, n49715, n49716, n49717, n49718, n49719, n49720, n49721, n49722, n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742, n49743, n49744, n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752, n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762, n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770, n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778, n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786, n49787, n49788, n49789, n49790, n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810, n49811, n49812, n49813, n49814, n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834, n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842, n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850, n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858, n49859, n49860, n49861, n49862, n49863, n49864, n49865, n49866, n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874, n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882, n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890, n49891, n49892, n49893, n49894, n49895, n49896, n49897, n49898, n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906, n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922, n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930, n49931, n49932, n49933, n49934, n49935, n49936, n49937, n49938, n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946, n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954, n49955, n49956, n49957, n49958, n49959, n49960, n49961, n49962, n49963, n49964, n49965, n49966, n49967, n49968, n49969, n49970, n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986, n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994, n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002, n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030, n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040, n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058, n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066, n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074, n50075, n50076, n50077, n50078, n50079, n50080, n50081, n50082, n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090, n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098, n50099, n50100, n50101, n50102, n50103, n50104, n50105, n50106, n50107, n50108, n50109, n50110, n50111, n50112, n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122, n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130, n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138, n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146, n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154, n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162, n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176, n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184, n50185, n50186, n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194, n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202, n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210, n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218, n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226, n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234, n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242, n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258, n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274, n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282, n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290, n50291, n50292, n50293, n50294, n50295, n50296, n50297, n50298, n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306, n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322, n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338, n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346, n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354, n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362, n50363, n50364, n50365, n50366, n50367, n50368, n50369, n50370, n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378, n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392, n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400, n50401, n50402, n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410, n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418, n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426, n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442, n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450, n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466, n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474, n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490, n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498, n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507, n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522, n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531, n50532, n50533, n50534, n50535, n50536, n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544, n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554, n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578, n50579, n50580, n50581, n50582, n50583, n50584, n50585, n50586, n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594, n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608, n50609, n50610, n50611, n50612, n50613, n50614, n50615, n50616, n50617, n50618, n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626, n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634, n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642, n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650, n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666, n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674, n50675, n50676, n50677, n50678, n50679, n50680, n50681, n50682, n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690, n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698, n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714, n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722, n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730, n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738, n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746, n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754, n50755, n50756, n50757, n50758, n50759, n50760, n50761, n50762, n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770, n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778, n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786, n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794, n50795, n50796, n50797, n50798, n50799, n50800, n50801, n50802, n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810, n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818, n50819, n50820, n50821, n50822, n50823, n50824, n50825, n50826, n50827, n50828, n50829, n50830, n50831, n50832, n50833, n50834, n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842, n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850, n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858, n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866, n50867, n50868, n50869, n50870, n50871, n50872, n50873, n50874, n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882, n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890, n50891, n50892, n50893, n50894, n50895, n50896, n50897, n50898, n50899, n50900, n50901, n50902, n50903, n50904, n50905, n50906, n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914, n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922, n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930, n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938, n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954, n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962, n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970, n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978, n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986, n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994, n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002, n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010, n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018, n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026, n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034, n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050, n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058, n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066, n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074, n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082, n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090, n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098, n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106, n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114, n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122, n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130, n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138, n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146, n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154, n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162, n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186, n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194, n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202, n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210, n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218, n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226, n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234, n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242, n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250, n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258, n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266, n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274, n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282, n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290, n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298, n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306, n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314, n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322, n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330, n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338, n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346, n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354, n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362, n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370, n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386, n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394, n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402, n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410, n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418, n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426, n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434, n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442, n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450, n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458, n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474, n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482, n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490, n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498, n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506, n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514, n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522, n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530, n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538, n51539, n51540, n51541, n51542, n51543, n51544, n51545, n51546, n51547, n51548, n51549, n51550, n51551, n51552, n51553, n51554, n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562, n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570, n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594, n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602, n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616, n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624, n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634, n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642, n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650, n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658, n51659, n51660, n51661, n51662, n51663, n51664, n51665, n51666, n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674, n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696, n51697, n51698, n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706, n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714, n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732, n51733, n51734, n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746, n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760, n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768, n51769, n51770, n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778, n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786, n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802, n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810, n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826, n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834, n51835, n51836, n51837, n51838, n51839, n51840, n51841, n51842, n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850, n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858, n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866, n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874, n51875, n51876, n51877, n51878, n51879, n51880, n51881, n51882, n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890, n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898, n51899, n51900, n51901, n51902, n51903, n51904, n51905, n51906, n51907, n51908, n51909, n51910, n51911, n51912, n51913, n51914, n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922, n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930, n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938, n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946, n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954, n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962, n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976, n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984, n51985, n51986, n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994, n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002, n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010, n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018, n52019, n52020, n52021, n52022, n52023, n52024, n52025, n52026, n52027, n52028, n52029, n52030, n52031, n52032, n52033, n52034, n52035, n52036, n52037, n52038, n52039, n52040, n52041, n52042, n52043, n52044, n52045, n52046, n52047, n52048, n52049, n52050, n52051, n52052, n52053, n52054, n52055, n52056, n52057, n52058, n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066, n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074, n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084, n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092, n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100, n52101, n52102, n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110, n52111, n52112, n52113, n52114, n52115, n52116, n52117, n52118, n52119, n52120, n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128, n52129, n52130, n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138, n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156, n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164, n52165, n52166, n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178, n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192, n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202, n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210, n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219, n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228, n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236, n52237, n52238, n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246, n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264, n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272, n52273, n52274, n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282, n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291, n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300, n52301, n52302, n52303, n52304, n52305, n52306, n52307, n52308, n52309, n52310, n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322, n52323, n52324, n52325, n52326, n52327, n52328, n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336, n52337, n52338, n52339, n52340, n52341, n52342, n52343, n52344, n52345, n52346, n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354, n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380, n52381, n52382, n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390, n52391, n52392, n52393, n52394, n52395, n52396, n52397, n52398, n52399, n52400, n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408, n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416, n52417, n52418, n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426, n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434, n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443, n52444, n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452, n52453, n52454, n52455, n52456, n52457, n52458, n52459, n52460, n52461, n52462, n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470, n52471, n52472, n52473, n52474, n52475, n52476, n52477, n52478, n52479, n52480, n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488, n52489, n52490, n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498, n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506, n52507, n52508, n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516, n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524, n52525, n52526, n52527, n52528, n52529, n52530, n52531, n52532, n52533, n52534, n52535, n52536, n52537, n52538, n52539, n52540, n52541, n52542, n52543, n52544, n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562, n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570, n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579, n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588, n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596, n52597, n52598, n52599, n52600, n52601, n52602, n52603, n52604, n52605, n52606, n52607, n52608, n52609, n52610, n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618, n52619, n52620, n52621, n52622, n52623, n52624, n52625, n52626, n52627, n52628, n52629, n52630, n52631, n52632, n52633, n52634, n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642, n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650, n52651, n52652, n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660, n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668, n52669, n52670, n52671, n52672, n52673, n52674, n52675, n52676, n52677, n52678, n52679, n52680, n52681, n52682, n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696, n52697, n52698, n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706, n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714, n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722, n52723, n52724, n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732, n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740, n52741, n52742, n52743, n52744, n52745, n52746, n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754, n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762, n52763, n52764, n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772, n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786, n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794, n52795, n52796, n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812, n52813, n52814, n52815, n52816, n52817, n52818, n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826, n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840, n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848, n52849, n52850, n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858, n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866, n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876, n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884, n52885, n52886, n52887, n52888, n52889, n52890, n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898, n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906, n52907, n52908, n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916, n52917, n52918, n52919, n52920, n52921, n52922, n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930, n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938, n52939, n52940, n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956, n52957, n52958, n52959, n52960, n52961, n52962, n52963, n52964, n52965, n52966, n52967, n52968, n52969, n52970, n52971, n52972, n52973, n52974, n52975, n52976, n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984, n52985, n52986, n52987, n52988, n52989, n52990, n52991, n52992, n52993, n52994, n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002, n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010, n53011, n53012, n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028, n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050, n53051, n53052, n53053, n53054, n53055, n53056, n53057, n53058, n53059, n53060, n53061, n53062, n53063, n53064, n53065, n53066, n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074, n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082, n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100, n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108, n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116, n53117, n53118, n53119, n53120, n53121, n53122, n53123, n53124, n53125, n53126, n53127, n53128, n53129, n53130, n53131, n53132, n53133, n53134, n53135, n53136, n53137, n53138, n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146, n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154, n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172, n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180, n53181, n53182, n53183, n53184, n53185, n53186, n53187, n53188, n53189, n53190, n53191, n53192, n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200, n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209, n53210, n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218, n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227, n53228, n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236, n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244, n53245, n53246, n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254, n53255, n53256, n53257, n53258, n53259, n53260, n53261, n53262, n53263, n53264, n53265, n53266, n53267, n53268, n53269, n53270, n53271, n53272, n53273, n53274, n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282, n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290, n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298, n53299, n53300, n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308, n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316, n53317, n53318, n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326, n53327, n53328, n53329, n53330, n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338, n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346, n53347, n53348, n53349, n53350, n53351, n53352, n53353, n53354, n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362, n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370, n53371, n53372, n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380, n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388, n53389, n53390, n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398, n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410, n53411, n53412, n53413, n53414, n53415, n53416, n53417, n53418, n53419, n53420, n53421, n53422, n53423, n53424, n53425, n53426, n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434, n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442, n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450, n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458, n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466, n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474, n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482, n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490, n53491, n53492, n53493, n53494, n53495, n53496, n53497, n53498, n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506, n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514, n53515, n53516, n53517, n53518, n53519, n53520, n53521, n53522, n53523, n53524, n53525, n53526, n53527, n53528, n53529, n53530, n53531, n53532, n53533, n53534, n53535, n53536, n53537, n53538, n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546, n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554, n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562, n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570, n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578, n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586, n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594, n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602, n53603, n53604, n53605, n53606, n53607, n53608, n53609, n53610, n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618, n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626, n53627, n53628, n53629, n53630, n53631, n53632, n53633, n53634, n53635, n53636, n53637, n53638, n53639, n53640, n53641, n53642, n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650, n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658, n53659, n53660, n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676, n53677, n53678, n53679, n53680, n53681, n53682, n53683, n53684, n53685, n53686, n53687, n53688, n53689, n53690, n53691, n53692, n53693, n53694, n53695, n53696, n53697, n53698, n53699, n53700, n53701, n53702, n53703, n53704, n53705, n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713, n53714, n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722, n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730, n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738, n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746, n53747, n53748, n53749, n53750, n53751, n53752, n53753, n53754, n53755, n53756, n53757, n53758, n53759, n53760, n53761, n53762, n53763, n53764, n53765, n53766, n53767, n53768, n53769, n53770, n53771, n53772, n53773, n53774, n53775, n53776, n53777, n53778, n53779, n53780, n53781, n53782, n53783, n53784, n53785, n53786, n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794, n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802, n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810, n53811, n53812, n53813, n53814, n53815, n53816, n53817, n53818, n53819, n53820, n53821, n53822, n53823, n53824, n53825, n53826, n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834, n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842, n53843, n53844, n53845, n53846, n53847, n53848, n53849, n53850, n53851, n53852, n53853, n53854, n53855, n53856, n53857, n53858, n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866, n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874, n53875, n53876, n53877, n53878, n53879, n53880, n53881, n53882, n53883, n53884, n53885, n53886, n53887, n53888, n53889, n53890, n53891, n53892, n53893, n53894, n53895, n53896, n53897, n53898, n53899, n53900, n53901, n53902, n53903, n53904, n53905, n53906, n53907, n53908, n53909, n53910, n53911, n53912, n53913, n53914, n53915, n53916, n53917, n53918, n53919, n53920, n53921, n53922, n53923, n53924, n53925, n53926, n53927, n53928, n53929, n53930, n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938, n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946, n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954, n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962, n53963, n53964, n53965, n53966, n53967, n53968, n53969, n53970, n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53978, n53979, n53980, n53981, n53982, n53983, n53984, n53985, n53986, n53987, n53988, n53989, n53990, n53991, n53992, n53993, n53994, n53995, n53996, n53997, n53998, n53999, n54000, n54001, n54002, n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010, n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018, n54019, n54020, n54021, n54022, n54023, n54024, n54025, n54026, n54027, n54028, n54029, n54030, n54031, n54032, n54033, n54034, n54035, n54036, n54037, n54038, n54039, n54040, n54041, n54042, n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050, n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058, n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066, n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074, n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082, n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090, n54091, n54092, n54093, n54094, n54095, n54096, n54097, n54098, n54099, n54100, n54101, n54102, n54103, n54104, n54105, n54106, n54107, n54108, n54109, n54110, n54111, n54112, n54113, n54114, n54115, n54116, n54117, n54118, n54119, n54120, n54121, n54122, n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130, n54131, n54132, n54133, n54134, n54135, n54136, n54137, n54138, n54139, n54140, n54141, n54142, n54143, n54144, n54145, n54146, n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154, n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162, n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170, n54171, n54172, n54173, n54174, n54175, n54176, n54177, n54178, n54179, n54180, n54181, n54182, n54183, n54184, n54185, n54186, n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194, n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202, n54203, n54204, n54205, n54206, n54207, n54208, n54209, n54210, n54211, n54212, n54213, n54214, n54215, n54216, n54217, n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226, n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234, n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242, n54243, n54244, n54245, n54246, n54247, n54248, n54249, n54250, n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258, n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266, n54267, n54268, n54269, n54270, n54271, n54272, n54273, n54274, n54275, n54276, n54277, n54278, n54279, n54280, n54281, n54282, n54283, n54284, n54285, n54286, n54287, n54288, n54289, n54290, n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298, n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306, n54307, n54308, n54309, n54310, n54311, n54312, n54313, n54314, n54315, n54316, n54317, n54318, n54319, n54320, n54321, n54322, n54323, n54324, n54325, n54326, n54327, n54328, n54329, n54330, n54331, n54332, n54333, n54334, n54335, n54336, n54337, n54338, n54339, n54340, n54341, n54342, n54343, n54344, n54345, n54346, n54347, n54348, n54349, n54350, n54351, n54352, n54353, n54354, n54355, n54356, n54357, n54358, n54359, n54360, n54361, n54362, n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370, n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378, n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386, n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394, n54395, n54396, n54397, n54398, n54399, n54400, n54401, n54402, n54403, n54404, n54405, n54406, n54407, n54408, n54409, n54410, n54411, n54412, n54413, n54414, n54415, n54416, n54417, n54418, n54419, n54420, n54421, n54422, n54423, n54424, n54425, n54426, n54427, n54428, n54429, n54430, n54431, n54432, n54433, n54434, n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442, n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450, n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458, n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466, n54467, n54468, n54469, n54470, n54471, n54472, n54473, n54474, n54475, n54476, n54477, n54478, n54479, n54480, n54481, n54482, n54483, n54484, n54485, n54486, n54487, n54488, n54489, n54490, n54491, n54492, n54493, n54494, n54495, n54496, n54497, n54498, n54499, n54500, n54501, n54502, n54503, n54504, n54505, n54506, n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514, n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522, n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530, n54531, n54532, n54533, n54534, n54535, n54536, n54537, n54538, n54539, n54540, n54541, n54542, n54543, n54544, n54545, n54546, n54547, n54548, n54549, n54550, n54551, n54552, n54553, n54554, n54555, n54556, n54557, n54558, n54559, n54560, n54561, n54562, n54563, n54564, n54565, n54566, n54567, n54568, n54569, n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577, n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586, n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594, n54595, n54596, n54597, n54598, n54599, n54600, n54601, n54602, n54603, n54604, n54605, n54606, n54607, n54608, n54609, n54610, n54611, n54612, n54613, n54614, n54615, n54616, n54617, n54618, n54619, n54620, n54621, n54622, n54623, n54624, n54625, n54626, n54627, n54628, n54629, n54630, n54631, n54632, n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640, n54641, n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658, n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666, n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674, n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682, n54683, n54684, n54685, n54686, n54687, n54688, n54689, n54690, n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698, n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706, n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714, n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722, n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730, n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738, n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746, n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754, n54755, n54756, n54757, n54758, n54759, n54760, n54761, n54762, n54763, n54764, n54765, n54766, n54767, n54768, n54769, n54770, n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778, n54779, n54780, n54781, n54782, n54783, n54784, n54785, n54786, n54787, n54788, n54789, n54790, n54791, n54792, n54793, n54794, n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802, n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810, n54811, n54812, n54813, n54814, n54815, n54816, n54817, n54818, n54819, n54820, n54821, n54822, n54823, n54824, n54825, n54826, n54827, n54828, n54829, n54830, n54831, n54832, n54833, n54834, n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842, n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850, n54851, n54852, n54853, n54854, n54855, n54856, n54857, n54858, n54859, n54860, n54861, n54862, n54863, n54864, n54865, n54866, n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874, n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882, n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890, n54891, n54892, n54893, n54894, n54895, n54896, n54897, n54898, n54899, n54900, n54901, n54902, n54903, n54904, n54905, n54906, n54907, n54908, n54909, n54910, n54911, n54912, n54913, n54914, n54915, n54916, n54917, n54918, n54919, n54920, n54921, n54922, n54923, n54924, n54925, n54926, n54927, n54928, n54929, n54930, n54931, n54932, n54933, n54934, n54935, n54936, n54937, n54938, n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946, n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954, n54955, n54956, n54957, n54958, n54959, n54960, n54961, n54962, n54963, n54964, n54965, n54966, n54967, n54968, n54969, n54970, n54971, n54972, n54973, n54974, n54975, n54976, n54977, n54978, n54979, n54980, n54981, n54982, n54983, n54984, n54985, n54986, n54987, n54988, n54989, n54990, n54991, n54992, n54993, n54994, n54995, n54996, n54997, n54998, n54999, n55000, n55001, n55002, n55003, n55004, n55005, n55006, n55007, n55008, n55009, n55010, n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018, n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026, n55027, n55028, n55029, n55030, n55031, n55032, n55033, n55034, n55035, n55036, n55037, n55038, n55039, n55040, n55041, n55042, n55043, n55044, n55045, n55046, n55047, n55048, n55049, n55050, n55051, n55052, n55053, n55054, n55055, n55056, n55057, n55058, n55059, n55060, n55061, n55062, n55063, n55064, n55065, n55066, n55067, n55068, n55069, n55070, n55071, n55072, n55073, n55074, n55075, n55076, n55077, n55078, n55079, n55080, n55081, n55082, n55083, n55084, n55085, n55086, n55087, n55088, n55089, n55090, n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098, n55099, n55100, n55101, n55102, n55103, n55104, n55105, n55106, n55107, n55108, n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116, n55117, n55118, n55119, n55120, n55121, n55122, n55123, n55124, n55125, n55126, n55127, n55128, n55129, n55130, n55131, n55132, n55133, n55134, n55135, n55136, n55137, n55138, n55139, n55140, n55141, n55142, n55143, n55144, n55145, n55146, n55147, n55148, n55149, n55150, n55151, n55152, n55153, n55154, n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162, n55163, n55164, n55165, n55166, n55167, n55168, n55169, n55170, n55171, n55172, n55173, n55174, n55175, n55176, n55177, n55178, n55179, n55180, n55181, n55182, n55183, n55184, n55185, n55186, n55187, n55188, n55189, n55190, n55191, n55192, n55193, n55194, n55195, n55196, n55197, n55198, n55199, n55200, n55201, n55202, n55203, n55204, n55205, n55206, n55207, n55208, n55209, n55210, n55211, n55212, n55213, n55214, n55215, n55216, n55217, n55218, n55219, n55220, n55221, n55222, n55223, n55224, n55225, n55226, n55227, n55228, n55229, n55230, n55231, n55232, n55233, n55234, n55235, n55236, n55237, n55238, n55239, n55240, n55241, n55242, n55243, n55244, n55245, n55246, n55247, n55248, n55249, n55250, n55251, n55252, n55253, n55254, n55255, n55256, n55257, n55258, n55259, n55260, n55261, n55262, n55263, n55264, n55265, n55266, n55267, n55268, n55269, n55270, n55271, n55272, n55273, n55274, n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55282, n55283, n55284, n55285, n55286, n55287, n55288, n55289, n55290, n55291, n55292, n55293, n55294, n55295, n55296, n55297, n55298, n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306, n55307, n55308, n55309, n55310, n55311, n55312, n55313, n55314, n55315, n55316, n55317, n55318, n55319, n55320, n55321, n55322, n55323, n55324, n55325, n55326, n55327, n55328, n55329, n55330, n55331, n55332, n55333, n55334, n55335, n55336, n55337, n55338, n55339, n55340, n55341, n55342, n55343, n55344, n55345, n55346, n55347, n55348, n55349, n55350, n55351, n55352, n55353, n55354, n55355, n55356, n55357, n55358, n55359, n55360, n55361, n55362, n55363, n55364, n55365, n55366, n55367, n55368, n55369, n55370, n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378, n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386, n55387, n55388, n55389, n55390, n55391, n55392, n55393, n55394, n55395, n55396, n55397, n55398, n55399, n55400, n55401, n55402, n55403, n55404, n55405, n55406, n55407, n55408, n55409, n55410, n55411, n55412, n55413, n55414, n55415, n55416, n55417, n55418, n55419, n55420, n55421, n55422, n55423, n55424, n55425, n55426, n55427, n55428, n55429, n55430, n55431, n55432, n55433, n55434, n55435, n55436, n55437, n55438, n55439, n55440, n55441, n55442, n55443, n55444, n55445, n55446, n55447, n55448, n55449, n55450, n55451, n55452, n55453, n55454, n55455, n55456, n55457, n55458, n55459, n55460, n55461, n55462, n55463, n55464, n55465, n55466, n55467, n55468, n55469, n55470, n55471, n55472, n55473, n55474, n55475, n55476, n55477, n55478, n55479, n55480, n55481, n55482, n55483, n55484, n55485, n55486, n55487, n55488, n55489, n55490, n55491, n55492, n55493, n55494, n55495, n55496, n55497, n55498, n55499, n55500, n55501, n55502, n55503, n55504, n55505, n55506, n55507, n55508, n55509, n55510, n55511, n55512, n55513, n55514, n55515, n55516, n55517, n55518, n55519, n55520, n55521, n55522, n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530, n55531, n55532, n55533, n55534, n55535, n55536, n55537, n55538, n55539, n55540, n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548, n55549, n55550, n55551, n55552, n55553, n55554, n55555, n55556, n55557, n55558, n55559, n55560, n55561, n55562, n55563, n55564, n55565, n55566, n55567, n55568, n55569, n55570, n55571, n55572, n55573, n55574, n55575, n55576, n55577, n55578, n55579, n55580, n55581, n55582, n55583, n55584, n55585, n55586, n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594, n55595, n55596, n55597, n55598, n55599, n55600, n55601, n55602, n55603, n55604, n55605, n55606, n55607, n55608, n55609, n55610, n55611, n55612, n55613, n55614, n55615, n55616, n55617, n55618, n55619, n55620, n55621, n55622, n55623, n55624, n55625, n55626, n55627, n55628, n55629, n55630, n55631, n55632, n55633, n55634, n55635, n55636, n55637, n55638, n55639, n55640, n55641, n55642, n55643, n55644, n55645, n55646, n55647, n55648, n55649, n55650, n55651, n55652, n55653, n55654, n55655, n55656, n55657, n55658, n55659, n55660, n55661, n55662, n55663, n55664, n55665, n55666, n55667, n55668, n55669, n55670, n55671, n55672, n55673, n55674, n55675, n55676, n55677, n55678, n55679, n55680, n55681, n55682, n55683, n55684, n55685, n55686, n55687, n55688, n55689, n55690, n55691, n55692, n55693, n55694, n55695, n55696, n55697, n55698, n55699, n55700, n55701, n55702, n55703, n55704, n55705, n55706, n55707, n55708, n55709, n55710, n55711, n55712, n55713, n55714, n55715, n55716, n55717, n55718, n55719, n55720, n55721, n55722, n55723, n55724, n55725, n55726, n55727, n55728, n55729, n55730, n55731, n55732, n55733, n55734, n55735, n55736, n55737, n55738, n55739, n55740, n55741, n55742, n55743, n55744, n55745, n55746, n55747, n55748, n55749, n55750, n55751, n55752, n55753, n55754, n55755, n55756, n55757, n55758, n55759, n55760, n55761, n55762, n55763, n55764, n55765, n55766, n55767, n55768, n55769, n55770, n55771, n55772, n55773, n55774, n55775, n55776, n55777, n55778, n55779, n55780, n55781, n55782, n55783, n55784, n55785, n55786, n55787, n55788, n55789, n55790, n55791, n55792, n55793, n55794, n55795, n55796, n55797, n55798, n55799, n55800, n55801, n55802, n55803, n55804, n55805, n55806, n55807, n55808, n55809, n55810, n55811, n55812, n55813, n55814, n55815, n55816, n55817, n55818, n55819, n55820, n55821, n55822, n55823, n55824, n55825, n55826, n55827, n55828, n55829, n55830, n55831, n55832, n55833, n55834, n55835, n55836, n55837, n55838, n55839, n55840, n55841, n55842, n55843, n55844, n55845, n55846, n55847, n55848, n55849, n55850, n55851, n55852, n55853, n55854, n55855, n55856, n55857, n55858, n55859, n55860, n55861, n55862, n55863, n55864, n55865, n55866, n55867, n55868, n55869, n55870, n55871, n55872, n55873, n55874, n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882, n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890, n55891, n55892, n55893, n55894, n55895, n55896, n55897, n55898, n55899, n55900, n55901, n55902, n55903, n55904, n55905, n55906, n55907, n55908, n55909, n55910, n55911, n55912, n55913, n55914, n55915, n55916, n55917, n55918, n55919, n55920, n55921, n55922, n55923, n55924, n55925, n55926, n55927, n55928, n55929, n55930, n55931, n55932, n55933, n55934, n55935, n55936, n55937, n55938, n55939, n55940, n55941, n55942, n55943, n55944, n55945, n55946, n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55954, n55955, n55956, n55957, n55958, n55959, n55960, n55961, n55962, n55963, n55964, n55965, n55966, n55967, n55968, n55969, n55970, n55971, n55972, n55973, n55974, n55975, n55976, n55977, n55978, n55979, n55980, n55981, n55982, n55983, n55984, n55985, n55986, n55987, n55988, n55989, n55990, n55991, n55992, n55993, n55994, n55995, n55996, n55997, n55998, n55999, n56000, n56001, n56002, n56003, n56004, n56005, n56006, n56007, n56008, n56009, n56010, n56011, n56012, n56013, n56014, n56015, n56016, n56017, n56018, n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026, n56027, n56028, n56029, n56030, n56031, n56032, n56033, n56034, n56035, n56036, n56037, n56038, n56039, n56040, n56041, n56042, n56043, n56044, n56045, n56046, n56047, n56048, n56049, n56050, n56051, n56052, n56053, n56054, n56055, n56056, n56057, n56058, n56059, n56060, n56061, n56062, n56063, n56064, n56065, n56066, n56067, n56068, n56069, n56070, n56071, n56072, n56073, n56074, n56075, n56076, n56077, n56078, n56079, n56080, n56081, n56082, n56083, n56084, n56085, n56086, n56087, n56088, n56089, n56090, n56091, n56092, n56093, n56094, n56095, n56096, n56097, n56098, n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106, n56107, n56108, n56109, n56110, n56111, n56112, n56113, n56114, n56115, n56116, n56117, n56118, n56119, n56120, n56121, n56122, n56123, n56124, n56125, n56126, n56127, n56128, n56129, n56130, n56131, n56132, n56133, n56134, n56135, n56136, n56137, n56138, n56139, n56140, n56141, n56142, n56143, n56144, n56145, n56146, n56147, n56148, n56149, n56150, n56151, n56152, n56153, n56154, n56155, n56156, n56157, n56158, n56159, n56160, n56161, n56162, n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170, n56171, n56172, n56173, n56174, n56175, n56176, n56177, n56178, n56179, n56180, n56181, n56182, n56183, n56184, n56185, n56186, n56187, n56188, n56189, n56190, n56191, n56192, n56193, n56194, n56195, n56196, n56197, n56198, n56199, n56200, n56201, n56202, n56203, n56204, n56205, n56206, n56207, n56208, n56209, n56210, n56211, n56212, n56213, n56214, n56215, n56216, n56217, n56218, n56219, n56220, n56221, n56222, n56223, n56224, n56225, n56226, n56227, n56228, n56229, n56230, n56231, n56232, n56233, n56234, n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242, n56243, n56244, n56245, n56246, n56247, n56248, n56249, n56250, n56251, n56252, n56253, n56254, n56255, n56256, n56257, n56258, n56259, n56260, n56261, n56262, n56263, n56264, n56265, n56266, n56267, n56268, n56269, n56270, n56271, n56272, n56273, n56274, n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282, n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290, n56291, n56292, n56293, n56294, n56295, n56296, n56297, n56298, n56299, n56300, n56301, n56302, n56303, n56304, n56305, n56306, n56307, n56308, n56309, n56310, n56311, n56312, n56313, n56314, n56315, n56316, n56317, n56318, n56319, n56320, n56321, n56322, n56323, n56324, n56325, n56326, n56327, n56328, n56329, n56330, n56331, n56332, n56333, n56334, n56335, n56336, n56337, n56338, n56339, n56340, n56341, n56342, n56343, n56344, n56345, n56346, n56347, n56348, n56349, n56350, n56351, n56352, n56353, n56354, n56355, n56356, n56357, n56358, n56359, n56360, n56361, n56362, n56363, n56364, n56365, n56366, n56367, n56368, n56369, n56370, n56371, n56372, n56373, n56374, n56375, n56376, n56377, n56378, n56379, n56380, n56381, n56382, n56383, n56384, n56385, n56386, n56387, n56388, n56389, n56390, n56391, n56392, n56393, n56394, n56395, n56396, n56397, n56398, n56399, n56400, n56401, n56402, n56403, n56404, n56405, n56406, n56407, n56408, n56409, n56410, n56411, n56412, n56413, n56414, n56415, n56416, n56417, n56418, n56419, n56420, n56421, n56422, n56423, n56424, n56425, n56426, n56427, n56428, n56429, n56430, n56431, n56432, n56433, n56434, n56435, n56436, n56437, n56438, n56439, n56440, n56441, n56442, n56443, n56444, n56445, n56446, n56447, n56448, n56449, n56450, n56451, n56452, n56453, n56454, n56455, n56456, n56457, n56458, n56459, n56460, n56461, n56462, n56463, n56464, n56465, n56466, n56467, n56468, n56469, n56470, n56471, n56472, n56473, n56474, n56475, n56476, n56477, n56478, n56479, n56480, n56481, n56482, n56483, n56484, n56485, n56486, n56487, n56488, n56489, n56490, n56491, n56492, n56493, n56494, n56495, n56496, n56497, n56498, n56499, n56500, n56501, n56502, n56503, n56504, n56505, n56506, n56507, n56508, n56509, n56510, n56511, n56512, n56513, n56514, n56515, n56516, n56517, n56518, n56519, n56520, n56521, n56522, n56523, n56524, n56525, n56526, n56527, n56528, n56529, n56530, n56531, n56532, n56533, n56534, n56535, n56536, n56537, n56538, n56539, n56540, n56541, n56542, n56543, n56544, n56545, n56546, n56547, n56548, n56549, n56550, n56551, n56552, n56553, n56554, n56555, n56556, n56557, n56558, n56559, n56560, n56561, n56562, n56563, n56564, n56565, n56566, n56567, n56568, n56569, n56570, n56571, n56572, n56573, n56574, n56575, n56576, n56577, n56578, n56579, n56580, n56581, n56582, n56583, n56584, n56585, n56586, n56587, n56588, n56589, n56590, n56591, n56592, n56593, n56594, n56595, n56596, n56597, n56598, n56599, n56600, n56601, n56602, n56603, n56604, n56605, n56606, n56607, n56608, n56609, n56610, n56611, n56612, n56613, n56614, n56615, n56616, n56617, n56618, n56619, n56620, n56621, n56622, n56623, n56624, n56625, n56626, n56627, n56628, n56629, n56630, n56631, n56632, n56633, n56634, n56635, n56636, n56637, n56638, n56639, n56640, n56641, n56642, n56643, n56644, n56645, n56646, n56647, n56648, n56649, n56650, n56651, n56652, n56653, n56654, n56655, n56656, n56657, n56658, n56659, n56660, n56661, n56662, n56663, n56664, n56665, n56666, n56667, n56668, n56669, n56670, n56671, n56672, n56673, n56674, n56675, n56676, n56677, n56678, n56679, n56680, n56681, n56682, n56683, n56684, n56685, n56686, n56687, n56688, n56689, n56690, n56691, n56692, n56693, n56694, n56695, n56696, n56697, n56698, n56699, n56700, n56701, n56702, n56703, n56704, n56705, n56706, n56707, n56708, n56709, n56710, n56711, n56712, n56713, n56714, n56715, n56716, n56717, n56718, n56719, n56720, n56721, n56722, n56723, n56724, n56725, n56726, n56727, n56728, n56729, n56730, n56731, n56732, n56733, n56734, n56735, n56736, n56737, n56738, n56739, n56740, n56741, n56742, n56743, n56744, n56745, n56746, n56747, n56748, n56749, n56750, n56751, n56752, n56753, n56754, n56755, n56756, n56757, n56758, n56759, n56760, n56761, n56762, n56763, n56764, n56765, n56766, n56767, n56768, n56769, n56770, n56771, n56772, n56773, n56774, n56775, n56776, n56777, n56778, n56779, n56780, n56781, n56782, n56783, n56784, n56785, n56786, n56787, n56788, n56789, n56790, n56791, n56792, n56793, n56794, n56795, n56796, n56797, n56798, n56799, n56800, n56801, n56802, n56803, n56804, n56805, n56806, n56807, n56808, n56809, n56810, n56811, n56812, n56813, n56814, n56815, n56816, n56817, n56818, n56819, n56820, n56821, n56822, n56823, n56824, n56825, n56826, n56827, n56828, n56829, n56830, n56831, n56832, n56833, n56834, n56835, n56836, n56837, n56838, n56839, n56840, n56841, n56842, n56843, n56844, n56845, n56846, n56847, n56848, n56849, n56850, n56851, n56852, n56853, n56854, n56855, n56856, n56857, n56858, n56859, n56860, n56861, n56862, n56863, n56864, n56865, n56866, n56867, n56868, n56869, n56870, n56871, n56872, n56873, n56874, n56875, n56876, n56877, n56878, n56879, n56880, n56881, n56882, n56883, n56884, n56885, n56886, n56887, n56888, n56889, n56890, n56891, n56892, n56893, n56894, n56895, n56896, n56897, n56898, n56899, n56900, n56901, n56902, n56903, n56904, n56905, n56906, n56907, n56908, n56909, n56910, n56911, n56912, n56913, n56914, n56915, n56916, n56917, n56918, n56919, n56920, n56921, n56922, n56923, n56924, n56925, n56926, n56927, n56928, n56929, n56930, n56931, n56932, n56933, n56934, n56935, n56936, n56937, n56938, n56939, n56940, n56941, n56942, n56943, n56944, n56945, n56946, n56947, n56948, n56949, n56950, n56951, n56952, n56953, n56954, n56955, n56956, n56957, n56958, n56959, n56960, n56961, n56962, n56963, n56964, n56965, n56966, n56967, n56968, n56969, n56970, n56971, n56972, n56973, n56974, n56975, n56976, n56977, n56978, n56979, n56980, n56981, n56982, n56983, n56984, n56985, n56986, n56987, n56988, n56989, n56990, n56991, n56992, n56993, n56994, n56995, n56996, n56997, n56998, n56999, n57000, n57001, n57002, n57003, n57004, n57005, n57006, n57007, n57008, n57009, n57010, n57011, n57012, n57013, n57014, n57015, n57016, n57017, n57018, n57019, n57020, n57021, n57022, n57023, n57024, n57025, n57026, n57027, n57028, n57029, n57030, n57031, n57032, n57033, n57034, n57035, n57036, n57037, n57038, n57039, n57040, n57041, n57042, n57043, n57044, n57045, n57046, n57047, n57048, n57049, n57050, n57051, n57052, n57053, n57054, n57055, n57056, n57057, n57058, n57059, n57060, n57061, n57062, n57063, n57064, n57065, n57066, n57067, n57068, n57069, n57070, n57071, n57072, n57073, n57074, n57075, n57076, n57077, n57078, n57079, n57080, n57081, n57082, n57083, n57084, n57085, n57086, n57087, n57088, n57089, n57090, n57091, n57092, n57093, n57094, n57095, n57096, n57097, n57098, n57099, n57100, n57101, n57102, n57103, n57104, n57105, n57106, n57107, n57108, n57109, n57110, n57111, n57112, n57113, n57114, n57115, n57116, n57117, n57118, n57119, n57120, n57121, n57122, n57123, n57124, n57125, n57126, n57127, n57128, n57129, n57130, n57131, n57132, n57133, n57134, n57135, n57136, n57137, n57138, n57139, n57140, n57141, n57142, n57143, n57144, n57145, n57146, n57147, n57148, n57149, n57150, n57151, n57152, n57153, n57154, n57155, n57156, n57157, n57158, n57159, n57160, n57161, n57162, n57163, n57164, n57165, n57166, n57167, n57168, n57169, n57170, n57171, n57172, n57173, n57174, n57175, n57176, n57177, n57178, n57179, n57180, n57181, n57182, n57183, n57184, n57185, n57186, n57187, n57188, n57189, n57190, n57191, n57192, n57193, n57194, n57195, n57196, n57197, n57198, n57199, n57200, n57201, n57202, n57203, n57204, n57205, n57206, n57207, n57208, n57209, n57210, n57211, n57212, n57213, n57214, n57215, n57216, n57217, n57218, n57219, n57220, n57221, n57222, n57223, n57224, n57225, n57226, n57227, n57228, n57229, n57230, n57231, n57232, n57233, n57234, n57235, n57236, n57237, n57238, n57239, n57240, n57241, n57242, n57243, n57244, n57245, n57246, n57247, n57248, n57249, n57250, n57251, n57252, n57253, n57254, n57255, n57256, n57257, n57258, n57259, n57260, n57261, n57262, n57263, n57264, n57265, n57266, n57267, n57268, n57269, n57270, n57271, n57272, n57273, n57274, n57275, n57276, n57277, n57278, n57279, n57280, n57281, n57282, n57283, n57284, n57285, n57286, n57287, n57288, n57289, n57290, n57291, n57292, n57293, n57294, n57295, n57296, n57297, n57298, n57299, n57300, n57301, n57302, n57303, n57304, n57305, n57306, n57307, n57308, n57309, n57310, n57311, n57312, n57313, n57314, n57315, n57316, n57317, n57318, n57319, n57320, n57321, n57322, n57323, n57324, n57325, n57326, n57327, n57328, n57329, n57330, n57331, n57332, n57333, n57334, n57335, n57336, n57337, n57338, n57339, n57340, n57341, n57342, n57343, n57344, n57345, n57346, n57347, n57348, n57349, n57350, n57351, n57352, n57353, n57354, n57355, n57356, n57357, n57358, n57359, n57360, n57361, n57362, n57363, n57364, n57365, n57366, n57367, n57368, n57369, n57370, n57371, n57372, n57373, n57374, n57375, n57376, n57377, n57378, n57379, n57380, n57381, n57382, n57383, n57384, n57385, n57386, n57387, n57388, n57389, n57390, n57391, n57392, n57393, n57394, n57395, n57396, n57397, n57398, n57399, n57400, n57401, n57402, n57403, n57404, n57405, n57406, n57407, n57408, n57409, n57410, n57411, n57412, n57413, n57414, n57415, n57416, n57417, n57418, n57419, n57420, n57421, n57422, n57423, n57424, n57425, n57426, n57427, n57428, n57429, n57430, n57431, n57432, n57433, n57434, n57435, n57436, n57437, n57438, n57439, n57440, n57441, n57442, n57443, n57444, n57445, n57446, n57447, n57448, n57449, n57450, n57451, n57452, n57453, n57454, n57455, n57456, n57457, n57458, n57459, n57460, n57461, n57462, n57463, n57464, n57465, n57466, n57467, n57468, n57469, n57470, n57471, n57472, n57473, n57474, n57475, n57476, n57477, n57478, n57479, n57480, n57481, n57482, n57483, n57484, n57485, n57486, n57487, n57488, n57489, n57490, n57491, n57492, n57493, n57494, n57495, n57496, n57497, n57498, n57499, n57500, n57501, n57502, n57503, n57504, n57505, n57506, n57507, n57508, n57509, n57510, n57511, n57512, n57513, n57514, n57515, n57516, n57517, n57518, n57519, n57520, n57521, n57522, n57523, n57524, n57525, n57526, n57527, n57528, n57529, n57530, n57531, n57532, n57533, n57534, n57535, n57536, n57537, n57538, n57539, n57540, n57541, n57542, n57543, n57544, n57545, n57546, n57547, n57548, n57549, n57550, n57551, n57552, n57553, n57554, n57555, n57556, n57557, n57558, n57559, n57560, n57561, n57562, n57563, n57564, n57565, n57566, n57567, n57568, n57569, n57570, n57571, n57572, n57573, n57574, n57575, n57576, n57577, n57578, n57579, n57580, n57581, n57582, n57583, n57584, n57585, n57586, n57587, n57588, n57589, n57590, n57591, n57592, n57593, n57594, n57595, n57596, n57597, n57598, n57599, n57600, n57601, n57602, n57603, n57604, n57605, n57606, n57607, n57608, n57609, n57610, n57611, n57612, n57613, n57614, n57615, n57616, n57617, n57618, n57619, n57620, n57621, n57622, n57623, n57624, n57625, n57626, n57627, n57628, n57629, n57630, n57631, n57632, n57633, n57634, n57635, n57636, n57637, n57638, n57639, n57640, n57641, n57642, n57643, n57644, n57645, n57646, n57647, n57648, n57649, n57650, n57651, n57652, n57653, n57654, n57655, n57656, n57657, n57658, n57659, n57660, n57661, n57662, n57663, n57664, n57665, n57666, n57667, n57668, n57669, n57670, n57671, n57672, n57673, n57674, n57675, n57676, n57677, n57678, n57679, n57680, n57681, n57682, n57683, n57684, n57685, n57686, n57687, n57688, n57689, n57690, n57691, n57692, n57693, n57694, n57695, n57696, n57697, n57698, n57699, n57700, n57701, n57702, n57703, n57704, n57705, n57706, n57707, n57708, n57709, n57710, n57711, n57712, n57713, n57714, n57715, n57716, n57717, n57718, n57719, n57720, n57721, n57722, n57723, n57724, n57725, n57726, n57727, n57728, n57729, n57730, n57731, n57732, n57733, n57734, n57735, n57736, n57737, n57738, n57739, n57740, n57741, n57742, n57743, n57744, n57745, n57746, n57747, n57748, n57749, n57750, n57751, n57752, n57753, n57754, n57755, n57756, n57757, n57758, n57759, n57760, n57761, n57762, n57763, n57764, n57765, n57766, n57767, n57768, n57769, n57770, n57771, n57772, n57773, n57774, n57775, n57776, n57777, n57778, n57779, n57780, n57781, n57782, n57783, n57784, n57785, n57786, n57787, n57788, n57789, n57790, n57791, n57792, n57793, n57794, n57795, n57796, n57797, n57798, n57799, n57800, n57801, n57802, n57803, n57804, n57805, n57806, n57807, n57808, n57809, n57810, n57811, n57812, n57813, n57814, n57815, n57816, n57817, n57818, n57819, n57820, n57821, n57822, n57823, n57824, n57825, n57826, n57827, n57828, n57829, n57830, n57831, n57832, n57833, n57834, n57835, n57836, n57837, n57838, n57839, n57840, n57841, n57842, n57843, n57844, n57845, n57846, n57847, n57848, n57849, n57850, n57851, n57852, n57853, n57854, n57855, n57856, n57857, n57858, n57859, n57860, n57861, n57862, n57863, n57864, n57865, n57866, n57867, n57868, n57869, n57870, n57871, n57872, n57873, n57874, n57875, n57876, n57877, n57878, n57879, n57880, n57881, n57882, n57883, n57884, n57885, n57886, n57887, n57888, n57889, n57890, n57891, n57892, n57893, n57894, n57895, n57896, n57897, n57898, n57899, n57900, n57901, n57902, n57903, n57904, n57905, n57906, n57907, n57908, n57909, n57910, n57911, n57912, n57913, n57914, n57915, n57916, n57917, n57918, n57919, n57920, n57921, n57922, n57923, n57924, n57925, n57926, n57927, n57928, n57929, n57930, n57931, n57932, n57933, n57934, n57935, n57936, n57937, n57938, n57939, n57940, n57941, n57942, n57943, n57944, n57945, n57946, n57947, n57948, n57949, n57950, n57951, n57952, n57953, n57954, n57955, n57956, n57957, n57958, n57959, n57960, n57961, n57962, n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970, n57971, n57972, n57973, n57974, n57975, n57976, n57977, n57978, n57979, n57980, n57981, n57982, n57983, n57984, n57985, n57986, n57987, n57988, n57989, n57990, n57991, n57992, n57993, n57994, n57995, n57996, n57997, n57998, n57999, n58000, n58001, n58002, n58003, n58004, n58005, n58006, n58007, n58008, n58009, n58010, n58011, n58012, n58013, n58014, n58015, n58016, n58017, n58018, n58019, n58020, n58021, n58022, n58023, n58024, n58025, n58026, n58027, n58028, n58029, n58030, n58031, n58032, n58033, n58034, n58035, n58036, n58037, n58038, n58039, n58040, n58041, n58042, n58043, n58044, n58045, n58046, n58047, n58048, n58049, n58050, n58051, n58052, n58053, n58054, n58055, n58056, n58057, n58058, n58059, n58060, n58061, n58062, n58063, n58064, n58065, n58066, n58067, n58068, n58069, n58070, n58071, n58072, n58073, n58074, n58075, n58076, n58077, n58078, n58079, n58080, n58081, n58082, n58083, n58084, n58085, n58086, n58087, n58088, n58089, n58090, n58091, n58092, n58093, n58094, n58095, n58096, n58097, n58098, n58099, n58100, n58101, n58102, n58103, n58104, n58105, n58106, n58107, n58108, n58109, n58110, n58111, n58112, n58113, n58114, n58115, n58116, n58117, n58118, n58119, n58120, n58121, n58122, n58123, n58124, n58125, n58126, n58127, n58128, n58129, n58130, n58131, n58132, n58133, n58134, n58135, n58136, n58137, n58138, n58139, n58140, n58141, n58142, n58143, n58144, n58145, n58146, n58147, n58148, n58149, n58150, n58151, n58152, n58153, n58154, n58155, n58156, n58157, n58158, n58159, n58160, n58161, n58162, n58163, n58164, n58165, n58166, n58167, n58168, n58169, n58170, n58171, n58172, n58173, n58174, n58175, n58176, n58177, n58178, n58179, n58180, n58181, n58182, n58183, n58184, n58185, n58186, n58187, n58188, n58189, n58190, n58191, n58192, n58193, n58194, n58195, n58196, n58197, n58198, n58199, n58200, n58201, n58202, n58203, n58204, n58205, n58206, n58207, n58208, n58209, n58210, n58211, n58212, n58213, n58214, n58215, n58216, n58217, n58218, n58219, n58220, n58221, n58222, n58223, n58224, n58225, n58226, n58227, n58228, n58229, n58230, n58231, n58232, n58233, n58234, n58235, n58236, n58237, n58238, n58239, n58240, n58241, n58242, n58243, n58244, n58245, n58246, n58247, n58248, n58249, n58250, n58251, n58252, n58253, n58254, n58255, n58256, n58257, n58258, n58259, n58260, n58261, n58262, n58263, n58264, n58265, n58266, n58267, n58268, n58269, n58270, n58271, n58272, n58273, n58274, n58275, n58276, n58277, n58278, n58279, n58280, n58281, n58282, n58283, n58284, n58285, n58286, n58287, n58288, n58289, n58290, n58291, n58292, n58293, n58294, n58295, n58296, n58297, n58298, n58299, n58300, n58301, n58302, n58303, n58304, n58305, n58306, n58307, n58308, n58309, n58310, n58311, n58312, n58313, n58314, n58315, n58316, n58317, n58318, n58319, n58320, n58321, n58322, n58323, n58324, n58325, n58326, n58327, n58328, n58329, n58330, n58331, n58332, n58333, n58334, n58335, n58336, n58337, n58338, n58339, n58340, n58341, n58342, n58343, n58344, n58345, n58346, n58347, n58348, n58349, n58350, n58351, n58352, n58353, n58354, n58355, n58356, n58357, n58358, n58359, n58360, n58361, n58362, n58363, n58364, n58365, n58366, n58367, n58368, n58369, n58370, n58371, n58372, n58373, n58374, n58375, n58376, n58377, n58378, n58379, n58380, n58381, n58382, n58383, n58384, n58385, n58386, n58387, n58388, n58389, n58390, n58391, n58392, n58393, n58394, n58395, n58396, n58397, n58398, n58399, n58400, n58401, n58402, n58403, n58404, n58405, n58406, n58407, n58408, n58409, n58410, n58411, n58412, n58413, n58414, n58415, n58416, n58417, n58418, n58419, n58420, n58421, n58422, n58423, n58424, n58425, n58426, n58427, n58428, n58429, n58430, n58431, n58432, n58433, n58434, n58435, n58436, n58437, n58438, n58439, n58440, n58441, n58442, n58443, n58444, n58445, n58446, n58447, n58448, n58449, n58450, n58451, n58452, n58453, n58454, n58455, n58456, n58457, n58458, n58459, n58460, n58461, n58462, n58463, n58464, n58465, n58466, n58467, n58468, n58469, n58470, n58471, n58472, n58473, n58474, n58475, n58476, n58477, n58478, n58479, n58480, n58481, n58482, n58483, n58484, n58485, n58486, n58487, n58488, n58489, n58490, n58491, n58492, n58493, n58494, n58495, n58496, n58497, n58498, n58499, n58500, n58501, n58502, n58503, n58504, n58505, n58506, n58507, n58508, n58509, n58510, n58511, n58512, n58513, n58514, n58515, n58516, n58517, n58518, n58519, n58520, n58521, n58522, n58523, n58524, n58525, n58526, n58527, n58528, n58529, n58530, n58531, n58532, n58533, n58534, n58535, n58536, n58537, n58538, n58539, n58540, n58541, n58542, n58543, n58544, n58545, n58546, n58547, n58548, n58549, n58550, n58551, n58552, n58553, n58554, n58555, n58556, n58557, n58558, n58559, n58560, n58561, n58562, n58563, n58564, n58565, n58566, n58567, n58568, n58569, n58570, n58571, n58572, n58573, n58574, n58575, n58576, n58577, n58578, n58579, n58580, n58581, n58582, n58583, n58584, n58585, n58586, n58587, n58588, n58589, n58590, n58591, n58592, n58593, n58594, n58595, n58596, n58597, n58598, n58599, n58600, n58601, n58602, n58603, n58604, n58605, n58606, n58607, n58608, n58609, n58610, n58611, n58612, n58613, n58614, n58615, n58616, n58617, n58618, n58619, n58620, n58621, n58622, n58623, n58624, n58625, n58626, n58627, n58628, n58629, n58630, n58631, n58632, n58633, n58634, n58635, n58636, n58637, n58638, n58639, n58640, n58641, n58642, n58643, n58644, n58645, n58646, n58647, n58648, n58649, n58650, n58651, n58652, n58653, n58654, n58655, n58656, n58657, n58658, n58659, n58660, n58661, n58662, n58663, n58664, n58665, n58666, n58667, n58668, n58669, n58670, n58671, n58672, n58673, n58674, n58675, n58676, n58677, n58678, n58679, n58680, n58681, n58682, n58683, n58684, n58685, n58686, n58687, n58688, n58689, n58690, n58691, n58692, n58693, n58694, n58695, n58696, n58697, n58698, n58699, n58700, n58701, n58702, n58703, n58704, n58705, n58706, n58707, n58708, n58709, n58710, n58711, n58712, n58713, n58714, n58715, n58716, n58717, n58718, n58719, n58720, n58721, n58722, n58723, n58724, n58725, n58726, n58727, n58728, n58729, n58730, n58731, n58732, n58733, n58734, n58735, n58736, n58737, n58738, n58739, n58740, n58741, n58742, n58743, n58744, n58745, n58746, n58747, n58748, n58749, n58750, n58751, n58752, n58753, n58754, n58755, n58756, n58757, n58758, n58759, n58760, n58761, n58762, n58763, n58764, n58765, n58766, n58767, n58768, n58769, n58770, n58771, n58772, n58773, n58774, n58775, n58776, n58777, n58778, n58779, n58780, n58781, n58782, n58783, n58784, n58785, n58786, n58787, n58788, n58789, n58790, n58791, n58792, n58793, n58794, n58795, n58796, n58797, n58798, n58799, n58800, n58801, n58802, n58803, n58804, n58805, n58806, n58807, n58808, n58809, n58810, n58811, n58812, n58813, n58814, n58815, n58816, n58817, n58818, n58819, n58820, n58821, n58822, n58823, n58824, n58825, n58826, n58827, n58828, n58829, n58830, n58831, n58832, n58833, n58834, n58835, n58836, n58837, n58838, n58839, n58840, n58841, n58842, n58843, n58844, n58845, n58846, n58847, n58848, n58849, n58850, n58851, n58852, n58853, n58854, n58855, n58856, n58857, n58858, n58859, n58860, n58861, n58862, n58863, n58864, n58865, n58866, n58867, n58868, n58869, n58870, n58871, n58872, n58873, n58874, n58875, n58876, n58877, n58878, n58879, n58880, n58881, n58882, n58883, n58884, n58885, n58886, n58887, n58888, n58889, n58890, n58891, n58892, n58893, n58894, n58895, n58896, n58897, n58898, n58899, n58900, n58901, n58902, n58903, n58904, n58905, n58906, n58907, n58908, n58909, n58910, n58911, n58912, n58913, n58914, n58915, n58916, n58917, n58918, n58919, n58920, n58921, n58922, n58923, n58924, n58925, n58926, n58927, n58928, n58929, n58930, n58931, n58932, n58933, n58934, n58935, n58936, n58937, n58938, n58939, n58940, n58941, n58942, n58943, n58944, n58945, n58946, n58947, n58948, n58949, n58950, n58951, n58952, n58953, n58954, n58955, n58956, n58957, n58958, n58959, n58960, n58961, n58962, n58963, n58964, n58965, n58966, n58967, n58968, n58969, n58970, n58971, n58972, n58973, n58974, n58975, n58976, n58977, n58978, n58979, n58980, n58981, n58982, n58983, n58984, n58985, n58986, n58987, n58988, n58989, n58990, n58991, n58992, n58993, n58994, n58995, n58996, n58997, n58998, n58999, n59000, n59001, n59002, n59003, n59004, n59005, n59006, n59007, n59008, n59009, n59010, n59011, n59012, n59013, n59014, n59015, n59016, n59017, n59018, n59019, n59020, n59021, n59022, n59023, n59024, n59025, n59026, n59027, n59028, n59029, n59030, n59031, n59032, n59033, n59034, n59035, n59036, n59037, n59038, n59039, n59040, n59041, n59042, n59043, n59044, n59045, n59046, n59047, n59048, n59049, n59050, n59051, n59052, n59053, n59054, n59055, n59056, n59057, n59058, n59059, n59060, n59061, n59062, n59063, n59064, n59065, n59066, n59067, n59068, n59069, n59070, n59071, n59072, n59073, n59074, n59075, n59076, n59077, n59078, n59079, n59080, n59081, n59082, n59083, n59084, n59085, n59086, n59087, n59088, n59089, n59090, n59091, n59092, n59093, n59094, n59095, n59096, n59097, n59098, n59099, n59100, n59101, n59102, n59103, n59104, n59105, n59106, n59107, n59108, n59109, n59110, n59111, n59112, n59113, n59114, n59115, n59116, n59117, n59118, n59119, n59120, n59121, n59122, n59123, n59124, n59125, n59126, n59127, n59128, n59129, n59130, n59131, n59132, n59133, n59134, n59135, n59136, n59137, n59138, n59139, n59140, n59141, n59142, n59143, n59144, n59145, n59146, n59147, n59148, n59149, n59150, n59151, n59152, n59153, n59154, n59155, n59156, n59157, n59158, n59159, n59160, n59161, n59162, n59163, n59164, n59165, n59166, n59167, n59168, n59169, n59170, n59171, n59172, n59173, n59174, n59175, n59176, n59177, n59178, n59179, n59180, n59181, n59182, n59183, n59184, n59185, n59186, n59187, n59188, n59189, n59190, n59191, n59192, n59193, n59194, n59195, n59196, n59197, n59198, n59199, n59200, n59201, n59202, n59203, n59204, n59205, n59206, n59207, n59208, n59209, n59210, n59211, n59212, n59213, n59214, n59215, n59216, n59217, n59218, n59219, n59220, n59221, n59222, n59223, n59224, n59225, n59226, n59227, n59228, n59229, n59230, n59231, n59232, n59233, n59234, n59235, n59236, n59237, n59238, n59239, n59240, n59241, n59242, n59243, n59244, n59245, n59246, n59247, n59248, n59249, n59250, n59251, n59252, n59253, n59254, n59255, n59256, n59257, n59258, n59259, n59260, n59261, n59262, n59263, n59264, n59265, n59266, n59267, n59268, n59269, n59270, n59271, n59272, n59273, n59274, n59275, n59276, n59277, n59278, n59279, n59280, n59281, n59282, n59283, n59284, n59285, n59286, n59287, n59288, n59289, n59290, n59291, n59292, n59293, n59294, n59295, n59296, n59297, n59298, n59299, n59300, n59301, n59302, n59303, n59304, n59305, n59306, n59307, n59308, n59309, n59310, n59311, n59312, n59313, n59314, n59315, n59316, n59317, n59318, n59319, n59320, n59321, n59322, n59323, n59324, n59325, n59326, n59327, n59328, n59329, n59330, n59331, n59332, n59333, n59334, n59335, n59336, n59337, n59338, n59339, n59340, n59341, n59342, n59343, n59344, n59345, n59346, n59347, n59348, n59349, n59350, n59351, n59352, n59353, n59354, n59355, n59356, n59357, n59358, n59359, n59360, n59361, n59362, n59363, n59364, n59365, n59366, n59367, n59368, n59369, n59370, n59371, n59372, n59373, n59374, n59375, n59376, n59377, n59378, n59379, n59380, n59381, n59382, n59383, n59384, n59385, n59386, n59387, n59388, n59389, n59390, n59391, n59392, n59393, n59394, n59395, n59396, n59397, n59398, n59399, n59400, n59401, n59402, n59403, n59404, n59405, n59406, n59407, n59408, n59409, n59410, n59411, n59412, n59413, n59414, n59415, n59416, n59417, n59418, n59419, n59420, n59421, n59422, n59423, n59424, n59425, n59426, n59427, n59428, n59429, n59430, n59431, n59432, n59433, n59434, n59435, n59436, n59437, n59438, n59439, n59440, n59441, n59442, n59443, n59444, n59445, n59446, n59447, n59448, n59449, n59450, n59451, n59452, n59453, n59454, n59455, n59456, n59457, n59458, n59459, n59460, n59461, n59462, n59463, n59464, n59465, n59466, n59467, n59468, n59469, n59470, n59471, n59472, n59473, n59474, n59475, n59476, n59477, n59478, n59479, n59480, n59481, n59482, n59483, n59484, n59485, n59486, n59487, n59488, n59489, n59490, n59491, n59492, n59493, n59494, n59495, n59496, n59497, n59498, n59499, n59500, n59501, n59502, n59503, n59504, n59505, n59506, n59507, n59508, n59509, n59510, n59511, n59512, n59513, n59514, n59515, n59516, n59517, n59518, n59519, n59520, n59521, n59522, n59523, n59524, n59525, n59526, n59527, n59528, n59529, n59530, n59531, n59532, n59533, n59534, n59535, n59536, n59537, n59538, n59539, n59540, n59541, n59542, n59543, n59544, n59545, n59546, n59547, n59548, n59549, n59550, n59551, n59552, n59553, n59554, n59555, n59556, n59557, n59558, n59559, n59560, n59561, n59562, n59563, n59564, n59565, n59566, n59567, n59568, n59569, n59570, n59571, n59572, n59573, n59574, n59575, n59576, n59577, n59578, n59579, n59580, n59581, n59582, n59583, n59584, n59585, n59586, n59587, n59588, n59589, n59590, n59591, n59592, n59593, n59594, n59595, n59596, n59597, n59598, n59599, n59600, n59601, n59602, n59603, n59604, n59605, n59606, n59607, n59608, n59609, n59610, n59611, n59612, n59613, n59614, n59615, n59616, n59617, n59618, n59619, n59620, n59621, n59622, n59623, n59624, n59625, n59626, n59627, n59628, n59629, n59630, n59631, n59632, n59633, n59634, n59635, n59636, n59637, n59638, n59639, n59640, n59641, n59642, n59643, n59644, n59645, n59646, n59647, n59648, n59649, n59650, n59651, n59652, n59653, n59654, n59655, n59656, n59657, n59658, n59659, n59660, n59661, n59662, n59663, n59664, n59665, n59666, n59667, n59668, n59669, n59670, n59671, n59672, n59673, n59674, n59675, n59676, n59677, n59678, n59679, n59680, n59681, n59682, n59683, n59684, n59685, n59686, n59687, n59688, n59689, n59690, n59691, n59692, n59693, n59694, n59695, n59696, n59697, n59698, n59699, n59700, n59701, n59702, n59703, n59704, n59705, n59706, n59707, n59708, n59709, n59710, n59711, n59712, n59713, n59714, n59715, n59716, n59717, n59718, n59719, n59720, n59721, n59722, n59723, n59724, n59725, n59726, n59727, n59728, n59729, n59730, n59731, n59732, n59733, n59734, n59735, n59736, n59737, n59738, n59739, n59740, n59741, n59742, n59743, n59744, n59745, n59746, n59747, n59748, n59749, n59750, n59751, n59752, n59753, n59754, n59755, n59756, n59757, n59758, n59759, n59760, n59761, n59762, n59763, n59764, n59765, n59766, n59767, n59768, n59769, n59770, n59771, n59772, n59773, n59774, n59775, n59776, n59777, n59778, n59779, n59780, n59781, n59782, n59783, n59784, n59785, n59786, n59787, n59788, n59789, n59790, n59791, n59792, n59793, n59794, n59795, n59796, n59797, n59798, n59799, n59800, n59801, n59802, n59803, n59804, n59805, n59806, n59807, n59808, n59809, n59810, n59811, n59812, n59813, n59814, n59815, n59816, n59817, n59818, n59819, n59820, n59821, n59822, n59823, n59824, n59825, n59826, n59827, n59828, n59829, n59830, n59831, n59832, n59833, n59834, n59835, n59836, n59837, n59838, n59839, n59840, n59841, n59842, n59843, n59844, n59845, n59846, n59847, n59848, n59849, n59850, n59851, n59852, n59853, n59854, n59855, n59856, n59857, n59858, n59859, n59860, n59861, n59862, n59863, n59864, n59865, n59866, n59867, n59868, n59869, n59870, n59871, n59872, n59873, n59874, n59875, n59876, n59877, n59878, n59879, n59880, n59881, n59882, n59883, n59884, n59885, n59886, n59887, n59888, n59889, n59890, n59891, n59892, n59893, n59894, n59895, n59896, n59897, n59898, n59899, n59900, n59901, n59902, n59903, n59904, n59905, n59906, n59907, n59908, n59909, n59910, n59911, n59912, n59913, n59914, n59915, n59916, n59917, n59918, n59919, n59920, n59921, n59922, n59923, n59924, n59925, n59926, n59927, n59928, n59929, n59930, n59931, n59932, n59933, n59934, n59935, n59936, n59937, n59938, n59939, n59940, n59941, n59942, n59943, n59944, n59945, n59946, n59947, n59948, n59949, n59950, n59951, n59952, n59953, n59954, n59955, n59956, n59957, n59958, n59959, n59960, n59961, n59962, n59963, n59964, n59965, n59966, n59967, n59968, n59969, n59970, n59971, n59972, n59973, n59974, n59975, n59976, n59977, n59978, n59979, n59980, n59981, n59982, n59983, n59984, n59985, n59986, n59987, n59988, n59989, n59990, n59991, n59992, n59993, n59994, n59995, n59996, n59997, n59998, n59999, n60000, n60001, n60002, n60003, n60004, n60005, n60006, n60007, n60008, n60009, n60010, n60011, n60012, n60013, n60014, n60015, n60016, n60017, n60018, n60019, n60020, n60021, n60022, n60023, n60024, n60025, n60026, n60027, n60028, n60029, n60030, n60031, n60032, n60033, n60034, n60035, n60036, n60037, n60038, n60039, n60040, n60041, n60042, n60043, n60044, n60045, n60046, n60047, n60048, n60049, n60050, n60051, n60052, n60053, n60054, n60055, n60056, n60057, n60058, n60059, n60060, n60061, n60062, n60063, n60064, n60065, n60066, n60067, n60068, n60069, n60070, n60071, n60072, n60073, n60074, n60075, n60076, n60077, n60078, n60079, n60080, n60081, n60082, n60083, n60084, n60085, n60086, n60087, n60088, n60089, n60090, n60091, n60092, n60093, n60094, n60095, n60096, n60097, n60098, n60099, n60100, n60101, n60102, n60103, n60104, n60105, n60106, n60107, n60108, n60109, n60110, n60111, n60112, n60113, n60114, n60115, n60116, n60117, n60118, n60119, n60120, n60121, n60122, n60123, n60124, n60125, n60126, n60127, n60128, n60129, n60130, n60131, n60132, n60133, n60134, n60135, n60136, n60137, n60138, n60139, n60140, n60141, n60142, n60143, n60144, n60145, n60146, n60147, n60148, n60149, n60150, n60151, n60152, n60153, n60154, n60155, n60156, n60157, n60158, n60159, n60160, n60161, n60162, n60163, n60164, n60165, n60166, n60167, n60168, n60169, n60170, n60171, n60172, n60173, n60174, n60175, n60176, n60177, n60178, n60179, n60180, n60181, n60182, n60183, n60184, n60185, n60186, n60187, n60188, n60189, n60190, n60191, n60192, n60193, n60194, n60195, n60196, n60197, n60198, n60199, n60200, n60201, n60202, n60203, n60204, n60205, n60206, n60207, n60208, n60209, n60210, n60211, n60212, n60213, n60214, n60215, n60216, n60217, n60218, n60219, n60220, n60221, n60222, n60223, n60224, n60225, n60226, n60227, n60228, n60229, n60230, n60231, n60232, n60233, n60234, n60235, n60236, n60237, n60238, n60239, n60240, n60241, n60242, n60243, n60244, n60245, n60246, n60247, n60248, n60249, n60250, n60251, n60252, n60253, n60254, n60255, n60256, n60257, n60258, n60259, n60260, n60261, n60262, n60263, n60264, n60265, n60266, n60267, n60268, n60269, n60270, n60271, n60272, n60273, n60274, n60275, n60276, n60277, n60278, n60279, n60280, n60281, n60282, n60283, n60284, n60285, n60286, n60287, n60288, n60289, n60290, n60291, n60292, n60293, n60294, n60295, n60296, n60297, n60298, n60299, n60300, n60301, n60302, n60303, n60304, n60305, n60306, n60307, n60308, n60309, n60310, n60311, n60312, n60313, n60314, n60315, n60316, n60317, n60318, n60319, n60320, n60321, n60322, n60323, n60324, n60325, n60326, n60327, n60328, n60329, n60330, n60331, n60332, n60333, n60334, n60335, n60336, n60337, n60338, n60339, n60340, n60341, n60342, n60343, n60344, n60345, n60346, n60347, n60348, n60349, n60350, n60351, n60352, n60353, n60354, n60355, n60356, n60357, n60358, n60359, n60360, n60361, n60362, n60363, n60364, n60365, n60366, n60367, n60368, n60369, n60370, n60371, n60372, n60373, n60374, n60375, n60376, n60377, n60378, n60379, n60380, n60381, n60382, n60383, n60384, n60385, n60386, n60387, n60388, n60389, n60390, n60391, n60392, n60393, n60394, n60395, n60396, n60397, n60398, n60399, n60400, n60401, n60402, n60403, n60404, n60405, n60406, n60407, n60408, n60409, n60410, n60411, n60412, n60413, n60414, n60415, n60416, n60417, n60418, n60419, n60420, n60421, n60422, n60423, n60424, n60425, n60426, n60427, n60428, n60429, n60430, n60431, n60432, n60433, n60434, n60435, n60436, n60437, n60438, n60439, n60440, n60441, n60442, n60443, n60444, n60445, n60446, n60447, n60448, n60449, n60450, n60451, n60452, n60453, n60454, n60455, n60456, n60457, n60458, n60459, n60460, n60461, n60462, n60463, n60464, n60465, n60466, n60467, n60468, n60469, n60470, n60471, n60472, n60473, n60474, n60475, n60476, n60477, n60478, n60479, n60480, n60481, n60482, n60483, n60484, n60485, n60486, n60487, n60488, n60489, n60490, n60491, n60492, n60493, n60494, n60495, n60496, n60497, n60498, n60499, n60500, n60501, n60502, n60503, n60504, n60505, n60506, n60507, n60508, n60509, n60510, n60511, n60512, n60513, n60514, n60515, n60516, n60517, n60518, n60519, n60520, n60521, n60522, n60523, n60524, n60525, n60526, n60527, n60528, n60529, n60530, n60531, n60532, n60533, n60534, n60535, n60536, n60537, n60538, n60539, n60540, n60541, n60542, n60543, n60544, n60545, n60546, n60547, n60548, n60549, n60550, n60551, n60552, n60553, n60554, n60555, n60556, n60557, n60558, n60559, n60560, n60561, n60562, n60563, n60564, n60565, n60566, n60567, n60568, n60569, n60570, n60571, n60572, n60573, n60574, n60575, n60576, n60577, n60578, n60579, n60580, n60581, n60582, n60583, n60584, n60585, n60586, n60587, n60588, n60589, n60590, n60591, n60592, n60593, n60594, n60595, n60596, n60597, n60598, n60599, n60600, n60601, n60602, n60603, n60604, n60605, n60606, n60607, n60608, n60609, n60610, n60611, n60612, n60613, n60614, n60615, n60616, n60617, n60618, n60619, n60620, n60621, n60622, n60623, n60624, n60625, n60626, n60627, n60628, n60629, n60630, n60631, n60632, n60633, n60634, n60635, n60636, n60637, n60638, n60639, n60640, n60641, n60642, n60643, n60644, n60645, n60646, n60647, n60648, n60649, n60650, n60651, n60652, n60653, n60654, n60655, n60656, n60657, n60658, n60659, n60660, n60661, n60662, n60663, n60664, n60665, n60666, n60667, n60668, n60669, n60670, n60671, n60672, n60673, n60674, n60675, n60676, n60677, n60678, n60679, n60680, n60681, n60682, n60683, n60684, n60685, n60686, n60687, n60688, n60689, n60690, n60691, n60692, n60693, n60694, n60695, n60696, n60697, n60698, n60699, n60700, n60701, n60702, n60703, n60704, n60705, n60706, n60707, n60708, n60709, n60710, n60711, n60712, n60713, n60714, n60715, n60716, n60717, n60718, n60719, n60720, n60721, n60722, n60723, n60724, n60725, n60726, n60727, n60728, n60729, n60730, n60731, n60732, n60733, n60734, n60735, n60736, n60737, n60738, n60739, n60740, n60741, n60742, n60743, n60744, n60745, n60746, n60747, n60748, n60749, n60750, n60751, n60752, n60753, n60754, n60755, n60756, n60757, n60758, n60759, n60760, n60761, n60762, n60763, n60764, n60765, n60766, n60767, n60768, n60769, n60770, n60771, n60772, n60773, n60774, n60775, n60776, n60777, n60778, n60779, n60780, n60781, n60782, n60783, n60784, n60785, n60786, n60787, n60788, n60789, n60790, n60791, n60792, n60793, n60794, n60795, n60796, n60797, n60798, n60799, n60800, n60801, n60802, n60803, n60804, n60805, n60806, n60807, n60808, n60809, n60810, n60811, n60812, n60813, n60814, n60815, n60816, n60817, n60818, n60819, n60820, n60821, n60822, n60823, n60824, n60825, n60826, n60827, n60828, n60829, n60830, n60831, n60832, n60833, n60834, n60835, n60836, n60837, n60838, n60839, n60840, n60841, n60842, n60843, n60844, n60845, n60846, n60847, n60848, n60849, n60850, n60851, n60852, n60853, n60854, n60855, n60856, n60857, n60858, n60859, n60860, n60861, n60862, n60863, n60864, n60865, n60866, n60867, n60868, n60869, n60870, n60871, n60872, n60873, n60874, n60875, n60876, n60877, n60878, n60879, n60880, n60881, n60882, n60883, n60884, n60885, n60886, n60887, n60888, n60889, n60890, n60891, n60892, n60893, n60894, n60895, n60896, n60897, n60898, n60899, n60900, n60901, n60902, n60903, n60904, n60905, n60906, n60907, n60908, n60909, n60910, n60911, n60912, n60913, n60914, n60915, n60916, n60917, n60918, n60919, n60920, n60921, n60922, n60923, n60924, n60925, n60926, n60927, n60928, n60929, n60930, n60931, n60932, n60933, n60934, n60935, n60936, n60937, n60938, n60939, n60940, n60941, n60942, n60943, n60944, n60945, n60946, n60947, n60948, n60949, n60950, n60951, n60952, n60953, n60954, n60955, n60956, n60957, n60958, n60959, n60960, n60961, n60962, n60963, n60964, n60965, n60966, n60967, n60968, n60969, n60970, n60971, n60972, n60973, n60974, n60975, n60976, n60977, n60978, n60979, n60980, n60981, n60982, n60983, n60984, n60985, n60986, n60987, n60988, n60989, n60990, n60991, n60992, n60993, n60994, n60995, n60996, n60997, n60998, n60999, n61000, n61001, n61002, n61003, n61004, n61005, n61006, n61007, n61008, n61009, n61010, n61011, n61012, n61013, n61014, n61015, n61016, n61017, n61018, n61019, n61020, n61021, n61022, n61023, n61024, n61025, n61026, n61027, n61028, n61029, n61030, n61031, n61032, n61033, n61034, n61035, n61036, n61037, n61038, n61039, n61040, n61041, n61042, n61043, n61044, n61045, n61046, n61047, n61048, n61049, n61050, n61051, n61052, n61053, n61054, n61055, n61056, n61057, n61058, n61059, n61060, n61061, n61062, n61063, n61064, n61065, n61066, n61067, n61068, n61069, n61070, n61071, n61072, n61073, n61074, n61075, n61076, n61077, n61078, n61079, n61080, n61081, n61082, n61083, n61084, n61085, n61086, n61087, n61088, n61089, n61090, n61091, n61092, n61093, n61094, n61095, n61096, n61097, n61098, n61099, n61100, n61101, n61102, n61103, n61104, n61105, n61106, n61107, n61108, n61109, n61110, n61111, n61112, n61113, n61114, n61115, n61116, n61117, n61118, n61119, n61120, n61121, n61122, n61123, n61124, n61125, n61126, n61127, n61128, n61129, n61130, n61131, n61132, n61133, n61134, n61135, n61136, n61137, n61138, n61139, n61140, n61141, n61142, n61143, n61144, n61145, n61146, n61147, n61148, n61149, n61150, n61151, n61152, n61153, n61154, n61155, n61156, n61157, n61158, n61159, n61160, n61161, n61162, n61163, n61164, n61165, n61166, n61167, n61168, n61169, n61170, n61171, n61172, n61173, n61174, n61175, n61176, n61177, n61178, n61179, n61180, n61181, n61182, n61183, n61184, n61185, n61186, n61187, n61188, n61189, n61190, n61191, n61192, n61193, n61194, n61195, n61196, n61197, n61198, n61199, n61200, n61201, n61202, n61203, n61204, n61205, n61206, n61207, n61208, n61209, n61210, n61211, n61212, n61213, n61214, n61215, n61216, n61217, n61218, n61219, n61220, n61221, n61222, n61223, n61224, n61225, n61226, n61227, n61228, n61229, n61230, n61231, n61232, n61233, n61234, n61235, n61236, n61237, n61238, n61239, n61240, n61241, n61242, n61243, n61244, n61245, n61246, n61247, n61248, n61249, n61250, n61251, n61252, n61253, n61254, n61255, n61256, n61257, n61258, n61259, n61260, n61261, n61262, n61263, n61264, n61265, n61266, n61267, n61268, n61269, n61270, n61271, n61272, n61273, n61274, n61275, n61276, n61277, n61278, n61279, n61280, n61281, n61282, n61283, n61284, n61285, n61286, n61287, n61288, n61289, n61290, n61291, n61292, n61293, n61294, n61295, n61296, n61297, n61298, n61299, n61300, n61301, n61302, n61303, n61304, n61305, n61306, n61307, n61308, n61309, n61310, n61311, n61312, n61313, n61314, n61315, n61316, n61317, n61318, n61319, n61320, n61321, n61322, n61323, n61324, n61325, n61326, n61327, n61328, n61329, n61330, n61331, n61332, n61333, n61334, n61335, n61336, n61337, n61338, n61339, n61340, n61341, n61342, n61343, n61344, n61345, n61346, n61347, n61348, n61349, n61350, n61351, n61352, n61353, n61354, n61355, n61356, n61357, n61358, n61359, n61360, n61361, n61362, n61363, n61364, n61365, n61366, n61367, n61368, n61369, n61370, n61371, n61372, n61373, n61374, n61375, n61376, n61377, n61378, n61379, n61380, n61381, n61382, n61383, n61384, n61385, n61386, n61387, n61388, n61389, n61390, n61391, n61392, n61393, n61394, n61395, n61396, n61397, n61398, n61399, n61400, n61401, n61402, n61403, n61404, n61405, n61406, n61407, n61408, n61409, n61410, n61411, n61412, n61413, n61414, n61415, n61416, n61417, n61418, n61419, n61420, n61421, n61422, n61423, n61424, n61425, n61426, n61427, n61428, n61429, n61430, n61431, n61432, n61433, n61434, n61435, n61436, n61437, n61438, n61439, n61440, n61441, n61442, n61443, n61444, n61445, n61446, n61447, n61448, n61449, n61450, n61451, n61452, n61453, n61454, n61455, n61456, n61457, n61458, n61459, n61460, n61461, n61462, n61463, n61464, n61465, n61466, n61467, n61468, n61469, n61470, n61471, n61472, n61473, n61474, n61475, n61476, n61477, n61478, n61479, n61480, n61481, n61482, n61483, n61484, n61485, n61486, n61487, n61488, n61489, n61490, n61491, n61492, n61493, n61494, n61495, n61496, n61497, n61498, n61499, n61500, n61501, n61502, n61503, n61504, n61505, n61506, n61507, n61508, n61509, n61510, n61511, n61512, n61513, n61514, n61515, n61516, n61517, n61518, n61519, n61520, n61521, n61522, n61523, n61524, n61525, n61526, n61527, n61528, n61529, n61530, n61531, n61532, n61533, n61534, n61535, n61536, n61537, n61538, n61539, n61540, n61541, n61542, n61543, n61544, n61545, n61546, n61547, n61548, n61549, n61550, n61551, n61552, n61553, n61554, n61555, n61556, n61557, n61558, n61559, n61560, n61561, n61562, n61563, n61564, n61565, n61566, n61567, n61568, n61569, n61570, n61571, n61572, n61573, n61574, n61575, n61576, n61577, n61578, n61579, n61580, n61581, n61582, n61583, n61584, n61585, n61586, n61587, n61588, n61589, n61590, n61591, n61592, n61593, n61594, n61595, n61596, n61597, n61598, n61599, n61600, n61601, n61602, n61603, n61604, n61605, n61606, n61607, n61608, n61609, n61610, n61611, n61612, n61613, n61614, n61615, n61616, n61617, n61618, n61619, n61620, n61621, n61622, n61623, n61624, n61625, n61626, n61627, n61628, n61629, n61630, n61631, n61632, n61633, n61634, n61635, n61636, n61637, n61638, n61639, n61640, n61641, n61642, n61643, n61644, n61645, n61646, n61647, n61648, n61649, n61650, n61651, n61652, n61653, n61654, n61655, n61656, n61657, n61658, n61659, n61660, n61661, n61662, n61663, n61664, n61665, n61666, n61667, n61668, n61669, n61670, n61671, n61672, n61673, n61674, n61675, n61676, n61677, n61678, n61679, n61680, n61681, n61682, n61683, n61684, n61685, n61686, n61687, n61688, n61689, n61690, n61691, n61692, n61693, n61694, n61695, n61696, n61697, n61698, n61699, n61700, n61701, n61702, n61703, n61704, n61705, n61706, n61707, n61708, n61709, n61710, n61711, n61712, n61713, n61714, n61715, n61716, n61717, n61718, n61719, n61720, n61721, n61722, n61723, n61724, n61725, n61726, n61727, n61728, n61729, n61730, n61731, n61732, n61733, n61734, n61735, n61736, n61737, n61738, n61739, n61740, n61741, n61742, n61743, n61744, n61745, n61746, n61747, n61748, n61749, n61750, n61751, n61752, n61753, n61754, n61755, n61756, n61757, n61758, n61759, n61760, n61761, n61762, n61763, n61764, n61765, n61766, n61767, n61768, n61769, n61770, n61771, n61772, n61773, n61774, n61775, n61776, n61777, n61778, n61779, n61780, n61781, n61782, n61783, n61784, n61785, n61786, n61787, n61788, n61789, n61790, n61791, n61792, n61793, n61794, n61795, n61796, n61797, n61798, n61799, n61800, n61801, n61802, n61803, n61804, n61805, n61806, n61807, n61808, n61809, n61810, n61811, n61812, n61813, n61814, n61815, n61816, n61817, n61818, n61819, n61820, n61821, n61822, n61823, n61824, n61825, n61826, n61827, n61828, n61829, n61830, n61831, n61832, n61833, n61834, n61835, n61836, n61837, n61838, n61839, n61840, n61841, n61842, n61843, n61844, n61845, n61846, n61847, n61848, n61849, n61850, n61851, n61852, n61853, n61854, n61855, n61856, n61857, n61858, n61859, n61860, n61861, n61862, n61863, n61864, n61865, n61866, n61867, n61868, n61869, n61870, n61871, n61872, n61873, n61874, n61875, n61876, n61877, n61878, n61879, n61880, n61881, n61882, n61883, n61884, n61885, n61886, n61887, n61888, n61889, n61890, n61891, n61892, n61893, n61894, n61895, n61896, n61897, n61898, n61899, n61900, n61901, n61902, n61903, n61904, n61905, n61906, n61907, n61908, n61909, n61910, n61911, n61912, n61913, n61914, n61915, n61916, n61917, n61918, n61919, n61920, n61921, n61922, n61923, n61924, n61925, n61926, n61927, n61928, n61929, n61930, n61931, n61932, n61933, n61934, n61935, n61936, n61937, n61938, n61939, n61940, n61941, n61942, n61943, n61944, n61945, n61946, n61947, n61948, n61949, n61950, n61951, n61952, n61953, n61954, n61955, n61956, n61957, n61958, n61959, n61960, n61961, n61962, n61963, n61964, n61965, n61966, n61967, n61968, n61969, n61970, n61971, n61972, n61973, n61974, n61975, n61976, n61977, n61978, n61979, n61980, n61981, n61982, n61983, n61984, n61985, n61986, n61987, n61988, n61989, n61990, n61991, n61992, n61993, n61994, n61995, n61996, n61997, n61998, n61999, n62000, n62001, n62002, n62003, n62004, n62005, n62006, n62007, n62008, n62009, n62010, n62011, n62012, n62013, n62014, n62015, n62016, n62017, n62018, n62019, n62020, n62021, n62022, n62023, n62024, n62025, n62026, n62027, n62028, n62029, n62030, n62031, n62032, n62033, n62034, n62035, n62036, n62037, n62038, n62039, n62040, n62041, n62042, n62043, n62044, n62045, n62046, n62047, n62048, n62049, n62050, n62051, n62052, n62053, n62054, n62055, n62056, n62057, n62058, n62059, n62060, n62061, n62062, n62063, n62064, n62065, n62066, n62067, n62068, n62069, n62070, n62071, n62072, n62073, n62074, n62075, n62076, n62077, n62078, n62079, n62080, n62081, n62082, n62083, n62084, n62085, n62086, n62087, n62088, n62089, n62090, n62091, n62092, n62093, n62094, n62095, n62096, n62097, n62098, n62099, n62100, n62101, n62102, n62103, n62104, n62105, n62106, n62107, n62108, n62109, n62110, n62111, n62112, n62113, n62114, n62115, n62116, n62117, n62118, n62119, n62120, n62121, n62122, n62123, n62124, n62125, n62126, n62127, n62128, n62129, n62130, n62131, n62132, n62133, n62134, n62135, n62136, n62137, n62138, n62139, n62140, n62141, n62142, n62143, n62144, n62145, n62146, n62147, n62148, n62149, n62150, n62151, n62152, n62153, n62154, n62155, n62156, n62157, n62158, n62159, n62160, n62161, n62162, n62163, n62164, n62165, n62166, n62167, n62168, n62169, n62170, n62171, n62172, n62173, n62174, n62175, n62176, n62177, n62178, n62179, n62180, n62181, n62182, n62183, n62184, n62185, n62186, n62187, n62188, n62189, n62190, n62191, n62192, n62193, n62194, n62195, n62196, n62197, n62198, n62199, n62200, n62201, n62202, n62203, n62204, n62205, n62206, n62207, n62208, n62209, n62210, n62211, n62212, n62213, n62214, n62215, n62216, n62217, n62218, n62219, n62220, n62221, n62222, n62223, n62224, n62225, n62226, n62227, n62228, n62229, n62230, n62231, n62232, n62233, n62234, n62235, n62236, n62237, n62238, n62239, n62240, n62241, n62242, n62243, n62244, n62245, n62246, n62247, n62248, n62249, n62250, n62251, n62252, n62253, n62254, n62255, n62256, n62257, n62258, n62259, n62260, n62261, n62262, n62263, n62264, n62265, n62266, n62267, n62268, n62269, n62270, n62271, n62272, n62273, n62274, n62275, n62276, n62277, n62278, n62279, n62280, n62281, n62282, n62283, n62284, n62285, n62286, n62287, n62288, n62289, n62290, n62291, n62292, n62293, n62294, n62295, n62296, n62297, n62298, n62299, n62300, n62301, n62302, n62303, n62304, n62305, n62306, n62307, n62308, n62309, n62310, n62311, n62312, n62313, n62314, n62315, n62316, n62317, n62318, n62319, n62320, n62321, n62322, n62323, n62324, n62325, n62326, n62327, n62328, n62329, n62330, n62331, n62332, n62333, n62334, n62335, n62336, n62337, n62338, n62339, n62340, n62341, n62342, n62343, n62344, n62345, n62346, n62347, n62348, n62349, n62350, n62351, n62352, n62353, n62354, n62355, n62356, n62357, n62358, n62359, n62360, n62361, n62362, n62363, n62364, n62365, n62366, n62367, n62368, n62369, n62370, n62371, n62372, n62373, n62374, n62375, n62376, n62377, n62378, n62379, n62380, n62381, n62382, n62383, n62384, n62385, n62386, n62387, n62388, n62389, n62390, n62391, n62392, n62393, n62394, n62395, n62396, n62397, n62398, n62399, n62400, n62401, n62402, n62403, n62404, n62405, n62406, n62407, n62408, n62409, n62410, n62411, n62412, n62413, n62414, n62415, n62416, n62417, n62418, n62419, n62420, n62421, n62422, n62423, n62424, n62425, n62426, n62427, n62428, n62429, n62430, n62431, n62432, n62433, n62434, n62435, n62436, n62437, n62438, n62439, n62440, n62441, n62442, n62443, n62444, n62445, n62446, n62447, n62448, n62449, n62450, n62451, n62452, n62453, n62454, n62455, n62456, n62457, n62458, n62459, n62460, n62461, n62462, n62463, n62464, n62465, n62466, n62467, n62468, n62469, n62470, n62471, n62472, n62473, n62474, n62475, n62476, n62477, n62478, n62479, n62480, n62481, n62482, n62483, n62484, n62485, n62486, n62487, n62488, n62489, n62490, n62491, n62492, n62493, n62494, n62495, n62496, n62497, n62498, n62499, n62500, n62501, n62502, n62503, n62504, n62505, n62506, n62507, n62508, n62509, n62510, n62511, n62512, n62513, n62514, n62515, n62516, n62517, n62518, n62519, n62520, n62521, n62522, n62523, n62524, n62525, n62526, n62527, n62528, n62529, n62530, n62531, n62532, n62533, n62534, n62535, n62536, n62537, n62538, n62539, n62540, n62541, n62542, n62543, n62544, n62545, n62546, n62547, n62548, n62549, n62550, n62551, n62552, n62553, n62554, n62555, n62556, n62557, n62558, n62559, n62560, n62561, n62562, n62563, n62564, n62565, n62566, n62567, n62568, n62569, n62570, n62571, n62572, n62573, n62574, n62575, n62576, n62577, n62578, n62579, n62580, n62581, n62582, n62583, n62584, n62585, n62586, n62587, n62588, n62589, n62590, n62591, n62592, n62593, n62594, n62595, n62596, n62597, n62598, n62599, n62600, n62601, n62602, n62603, n62604, n62605, n62606, n62607, n62608, n62609, n62610, n62611, n62612, n62613, n62614, n62615, n62616, n62617, n62618, n62619, n62620, n62621, n62622, n62623, n62624, n62625, n62626, n62627, n62628, n62629, n62630, n62631, n62632, n62633, n62634, n62635, n62636, n62637, n62638, n62639, n62640, n62641, n62642, n62643, n62644, n62645, n62646, n62647, n62648, n62649, n62650, n62651, n62652, n62653, n62654, n62655, n62656, n62657, n62658, n62659, n62660, n62661, n62662, n62663, n62664, n62665, n62666, n62667, n62668, n62669, n62670, n62671, n62672, n62673, n62674, n62675, n62676, n62677, n62678, n62679, n62680, n62681, n62682, n62683, n62684, n62685, n62686, n62687, n62688, n62689, n62690, n62691, n62692, n62693, n62694, n62695, n62696, n62697, n62698, n62699, n62700, n62701, n62702, n62703, n62704, n62705, n62706, n62707, n62708, n62709, n62710, n62711, n62712, n62713, n62714, n62715, n62716, n62717, n62718, n62719, n62720, n62721, n62722, n62723, n62724, n62725, n62726, n62727, n62728, n62729, n62730, n62731, n62732, n62733, n62734, n62735, n62736, n62737, n62738, n62739, n62740, n62741, n62742, n62743, n62744, n62745, n62746, n62747, n62748, n62749, n62750, n62751, n62752, n62753, n62754, n62755, n62756, n62757, n62758, n62759, n62760, n62761, n62762, n62763, n62764, n62765, n62766, n62767, n62768, n62769, n62770, n62771, n62772, n62773, n62774, n62775, n62776, n62777, n62778, n62779, n62780, n62781, n62782, n62783, n62784, n62785, n62786, n62787, n62788, n62789, n62790, n62791, n62792, n62793, n62794, n62795, n62796, n62797, n62798, n62799, n62800, n62801, n62802, n62803, n62804, n62805, n62806, n62807, n62808, n62809, n62810, n62811, n62812, n62813, n62814, n62815, n62816, n62817, n62818, n62819, n62820, n62821, n62822, n62823, n62824, n62825, n62826, n62827, n62828, n62829, n62830, n62831, n62832, n62833, n62834, n62835, n62836, n62837, n62838, n62839, n62840, n62841, n62842, n62843, n62844, n62845, n62846, n62847, n62848, n62849, n62850, n62851, n62852, n62853, n62854, n62855, n62856, n62857, n62858, n62859, n62860, n62861, n62862, n62863, n62864, n62865, n62866, n62867, n62868, n62869, n62870, n62871, n62872, n62873, n62874, n62875, n62876, n62877, n62878, n62879, n62880, n62881, n62882, n62883, n62884, n62885, n62886, n62887, n62888, n62889, n62890, n62891, n62892, n62893, n62894, n62895, n62896, n62897, n62898, n62899, n62900, n62901, n62902, n62903, n62904, n62905, n62906, n62907, n62908, n62909, n62910, n62911, n62912, n62913, n62914, n62915, n62916, n62917, n62918, n62919, n62920, n62921, n62922, n62923, n62924, n62925, n62926, n62927, n62928, n62929, n62930, n62931, n62932, n62933, n62934, n62935, n62936, n62937, n62938, n62939, n62940, n62941, n62942, n62943, n62944, n62945, n62946, n62947, n62948, n62949, n62950, n62951, n62952, n62953, n62954, n62955, n62956, n62957, n62958, n62959, n62960, n62961, n62962, n62963, n62964, n62965, n62966, n62967, n62968, n62969, n62970, n62971, n62972, n62973, n62974, n62975, n62976, n62977, n62978, n62979, n62980, n62981, n62982, n62983, n62984, n62985, n62986, n62987, n62988, n62989, n62990, n62991, n62992, n62993, n62994, n62995, n62996, n62997, n62998, n62999, n63000, n63001, n63002, n63003, n63004, n63005, n63006, n63007, n63008, n63009, n63010, n63011, n63012, n63013, n63014, n63015, n63016, n63017, n63018, n63019, n63020, n63021, n63022, n63023, n63024, n63025, n63026, n63027, n63028, n63029, n63030, n63031, n63032, n63033, n63034, n63035, n63036, n63037, n63038, n63039, n63040, n63041, n63042, n63043, n63044, n63045, n63046, n63047, n63048, n63049, n63050, n63051, n63052, n63053, n63054, n63055, n63056, n63057, n63058, n63059, n63060, n63061, n63062, n63063, n63064, n63065, n63066, n63067, n63068, n63069, n63070, n63071, n63072, n63073, n63074, n63075, n63076, n63077, n63078, n63079, n63080, n63081, n63082, n63083, n63084, n63085, n63086, n63087, n63088, n63089, n63090, n63091, n63092, n63093, n63094, n63095, n63096, n63097, n63098, n63099, n63100, n63101, n63102, n63103, n63104, n63105, n63106, n63107, n63108, n63109, n63110, n63111, n63112, n63113, n63114, n63115, n63116, n63117, n63118, n63119, n63120, n63121, n63122, n63123, n63124, n63125, n63126, n63127, n63128, n63129, n63130, n63131, n63132, n63133, n63134, n63135, n63136, n63137, n63138, n63139, n63140, n63141, n63142, n63143, n63144, n63145, n63146, n63147, n63148, n63149, n63150, n63151, n63152, n63153, n63154, n63155, n63156, n63157, n63158, n63159, n63160, n63161, n63162, n63163, n63164, n63165, n63166, n63167, n63168, n63169, n63170, n63171, n63172, n63173, n63174, n63175, n63176, n63177, n63178, n63179, n63180, n63181, n63182, n63183, n63184, n63185, n63186, n63187, n63188, n63189, n63190, n63191, n63192, n63193, n63194, n63195, n63196, n63197, n63198, n63199, n63200, n63201, n63202, n63203, n63204, n63205, n63206, n63207, n63208, n63209, n63210, n63211, n63212, n63213, n63214, n63215, n63216, n63217, n63218, n63219, n63220, n63221, n63222, n63223, n63224, n63225, n63226, n63227, n63228, n63229, n63230, n63231, n63232, n63233, n63234, n63235, n63236, n63237, n63238, n63239, n63240, n63241, n63242, n63243, n63244, n63245, n63246, n63247, n63248, n63249, n63250, n63251, n63252, n63253, n63254, n63255, n63256, n63257, n63258, n63259, n63260, n63261, n63262, n63263, n63264, n63265, n63266, n63267, n63268, n63269, n63270, n63271, n63272, n63273, n63274, n63275, n63276, n63277, n63278, n63279, n63280, n63281, n63282, n63283, n63284, n63285, n63286, n63287, n63288, n63289, n63290, n63291, n63292, n63293, n63294, n63295, n63296, n63297, n63298, n63299, n63300, n63301, n63302, n63303, n63304, n63305, n63306, n63307, n63308, n63309, n63310, n63311, n63312, n63313, n63314, n63315, n63316, n63317, n63318, n63319, n63320, n63321, n63322, n63323, n63324, n63325, n63326, n63327, n63328, n63329, n63330, n63331, n63332, n63333, n63334, n63335, n63336, n63337, n63338, n63339, n63340, n63341, n63342, n63343, n63344, n63345, n63346, n63347, n63348, n63349, n63350, n63351, n63352, n63353, n63354, n63355, n63356, n63357, n63358, n63359, n63360, n63361, n63362, n63363, n63364, n63365, n63366, n63367, n63368, n63369, n63370, n63371, n63372, n63373, n63374, n63375, n63376, n63377, n63378, n63379, n63380, n63381, n63382, n63383, n63384, n63385, n63386, n63387, n63388, n63389, n63390, n63391, n63392, n63393, n63394, n63395, n63396, n63397, n63398, n63399, n63400, n63401, n63402, n63403, n63404, n63405, n63406, n63407, n63408, n63409, n63410, n63411, n63412, n63413, n63414, n63415, n63416, n63417, n63418, n63419, n63420, n63421, n63422, n63423, n63424, n63425, n63426, n63427, n63428, n63429, n63430, n63431, n63432, n63433, n63434, n63435, n63436, n63437, n63438, n63439, n63440, n63441, n63442, n63443, n63444, n63445, n63446, n63447, n63448, n63449, n63450, n63451, n63452, n63453, n63454, n63455, n63456, n63457, n63458, n63459, n63460, n63461, n63462, n63463, n63464, n63465, n63466, n63467, n63468, n63469, n63470, n63471, n63472, n63473, n63474, n63475, n63476, n63477, n63478, n63479, n63480, n63481, n63482, n63483, n63484, n63485, n63486, n63487, n63488, n63489, n63490, n63491, n63492, n63493, n63494, n63495, n63496, n63497, n63498, n63499, n63500, n63501, n63502, n63503, n63504, n63505, n63506, n63507, n63508, n63509, n63510, n63511, n63512, n63513, n63514, n63515, n63516, n63517, n63518, n63519, n63520, n63521, n63522, n63523, n63524, n63525, n63526, n63527, n63528, n63529, n63530, n63531, n63532, n63533, n63534, n63535, n63536, n63537, n63538, n63539, n63540, n63541, n63542, n63543, n63544, n63545, n63546, n63547, n63548, n63549, n63550, n63551, n63552, n63553, n63554, n63555, n63556, n63557, n63558, n63559, n63560, n63561, n63562, n63563, n63564, n63565, n63566, n63567, n63568, n63569, n63570, n63571, n63572, n63573, n63574, n63575, n63576, n63577, n63578, n63579, n63580, n63581, n63582, n63583, n63584, n63585, n63586, n63587, n63588, n63589, n63590, n63591, n63592, n63593, n63594, n63595, n63596, n63597, n63598, n63599, n63600, n63601, n63602, n63603, n63604, n63605, n63606, n63607, n63608, n63609, n63610, n63611, n63612, n63613, n63614, n63615, n63616, n63617, n63618, n63619, n63620, n63621, n63622, n63623, n63624, n63625, n63626, n63627, n63628, n63629, n63630, n63631, n63632, n63633, n63634, n63635, n63636, n63637, n63638, n63639, n63640, n63641, n63642, n63643, n63644, n63645, n63646, n63647, n63648, n63649, n63650, n63651, n63652, n63653, n63654, n63655, n63656, n63657, n63658, n63659, n63660, n63661, n63662, n63663, n63664, n63665, n63666, n63667, n63668, n63669, n63670, n63671, n63672, n63673, n63674, n63675, n63676, n63677, n63678, n63679, n63680, n63681, n63682, n63683, n63684, n63685, n63686, n63687, n63688, n63689, n63690, n63691, n63692, n63693, n63694, n63695, n63696, n63697, n63698, n63699, n63700, n63701, n63702, n63703, n63704, n63705, n63706, n63707, n63708, n63709, n63710, n63711, n63712, n63713, n63714, n63715, n63716, n63717, n63718, n63719, n63720, n63721, n63722, n63723, n63724, n63725, n63726, n63727, n63728, n63729, n63730, n63731, n63732, n63733, n63734, n63735, n63736, n63737, n63738, n63739, n63740, n63741, n63742, n63743, n63744, n63745, n63746, n63747, n63748, n63749, n63750, n63751, n63752, n63753, n63754, n63755, n63756, n63757, n63758, n63759, n63760, n63761, n63762, n63763, n63764, n63765, n63766, n63767, n63768, n63769, n63770, n63771, n63772, n63773, n63774, n63775, n63776, n63777, n63778, n63779, n63780, n63781, n63782, n63783, n63784, n63785, n63786, n63787, n63788, n63789, n63790, n63791, n63792, n63793, n63794, n63795, n63796, n63797, n63798, n63799, n63800, n63801, n63802, n63803, n63804, n63805, n63806, n63807, n63808, n63809, n63810, n63811, n63812, n63813, n63814, n63815, n63816, n63817, n63818, n63819, n63820, n63821, n63822, n63823, n63824, n63825, n63826, n63827, n63828, n63829, n63830, n63831, n63832, n63833, n63834, n63835, n63836, n63837, n63838, n63839, n63840, n63841, n63842, n63843, n63844, n63845, n63846, n63847, n63848, n63849, n63850, n63851, n63852, n63853, n63854, n63855, n63856, n63857, n63858, n63859, n63860, n63861, n63862, n63863, n63864, n63865, n63866, n63867, n63868, n63869, n63870, n63871, n63872, n63873, n63874, n63875, n63876, n63877, n63878, n63879, n63880, n63881, n63882, n63883, n63884, n63885, n63886, n63887, n63888, n63889, n63890, n63891, n63892, n63893, n63894, n63895, n63896, n63897, n63898, n63899, n63900, n63901, n63902, n63903, n63904, n63905, n63906, n63907, n63908, n63909, n63910, n63911, n63912, n63913, n63914, n63915, n63916, n63917, n63918, n63919, n63920, n63921, n63922, n63923, n63924, n63925, n63926, n63927, n63928, n63929, n63930, n63931, n63932, n63933, n63934, n63935, n63936, n63937, n63938, n63939, n63940, n63941, n63942, n63943, n63944, n63945, n63946, n63947, n63948, n63949, n63950, n63951, n63952, n63953, n63954, n63955, n63956, n63957, n63958, n63959, n63960, n63961, n63962, n63963, n63964, n63965, n63966, n63967, n63968, n63969, n63970, n63971, n63972, n63973, n63974, n63975, n63976, n63977, n63978, n63979, n63980, n63981, n63982, n63983, n63984, n63985, n63986, n63987, n63988, n63989, n63990, n63991, n63992, n63993, n63994, n63995, n63996, n63997, n63998, n63999, n64000, n64001, n64002, n64003, n64004, n64005, n64006, n64007, n64008, n64009, n64010, n64011, n64012, n64013, n64014, n64015, n64016, n64017, n64018, n64019, n64020, n64021, n64022, n64023, n64024, n64025, n64026, n64027, n64028, n64029, n64030, n64031, n64032, n64033, n64034, n64035, n64036, n64037, n64038, n64039, n64040, n64041, n64042, n64043, n64044, n64045, n64046, n64047, n64048, n64049, n64050, n64051, n64052, n64053, n64054, n64055, n64056, n64057, n64058, n64059, n64060, n64061, n64062, n64063, n64064, n64065, n64066, n64067, n64068, n64069, n64070, n64071, n64072, n64073, n64074, n64075, n64076, n64077, n64078, n64079, n64080, n64081, n64082, n64083, n64084, n64085, n64086, n64087, n64088, n64089, n64090, n64091, n64092, n64093, n64094, n64095, n64096, n64097, n64098, n64099, n64100, n64101, n64102, n64103, n64104, n64105, n64106, n64107, n64108, n64109, n64110, n64111, n64112, n64113, n64114, n64115, n64116, n64117, n64118, n64119, n64120, n64121, n64122, n64123, n64124, n64125, n64126, n64127, n64128, n64129, n64130, n64131, n64132, n64133, n64134, n64135, n64136, n64137, n64138, n64139, n64140, n64141, n64142, n64143, n64144, n64145, n64146, n64147, n64148, n64149, n64150, n64151, n64152, n64153, n64154, n64155, n64156, n64157, n64158, n64159, n64160, n64161, n64162, n64163, n64164, n64165, n64166, n64167, n64168, n64169, n64170, n64171, n64172, n64173, n64174, n64175, n64176, n64177, n64178, n64179, n64180, n64181, n64182, n64183, n64184, n64185, n64186, n64187, n64188, n64189, n64190, n64191, n64192, n64193, n64194, n64195, n64196, n64197, n64198, n64199, n64200, n64201, n64202, n64203, n64204, n64205, n64206, n64207, n64208, n64209, n64210, n64211, n64212, n64213, n64214, n64215, n64216, n64217, n64218, n64219, n64220, n64221, n64222, n64223, n64224, n64225, n64226, n64227, n64228, n64229, n64230, n64231, n64232, n64233, n64234, n64235, n64236, n64237, n64238, n64239, n64240, n64241, n64242, n64243, n64244, n64245, n64246, n64247, n64248, n64249, n64250, n64251, n64252, n64253, n64254, n64255, n64256, n64257, n64258, n64259, n64260, n64261, n64262, n64263, n64264, n64265, n64266, n64267, n64268, n64269, n64270, n64271, n64272, n64273, n64274, n64275, n64276, n64277, n64278, n64279, n64280, n64281, n64282, n64283, n64284, n64285, n64286, n64287, n64288, n64289, n64290, n64291, n64292, n64293, n64294, n64295, n64296, n64297, n64298, n64299, n64300, n64301, n64302, n64303, n64304, n64305, n64306, n64307, n64308, n64309, n64310, n64311, n64312, n64313, n64314, n64315, n64316, n64317, n64318, n64319, n64320, n64321, n64322, n64323, n64324, n64325, n64326, n64327, n64328, n64329, n64330, n64331, n64332, n64333, n64334, n64335, n64336, n64337, n64338, n64339, n64340, n64341, n64342, n64343, n64344, n64345, n64346, n64347, n64348, n64349, n64350, n64351, n64352, n64353, n64354, n64355, n64356, n64357, n64358, n64359, n64360, n64361, n64362, n64363, n64364, n64365, n64366, n64367, n64368, n64369, n64370, n64371, n64372, n64373, n64374, n64375, n64376, n64377, n64378, n64379, n64380, n64381, n64382, n64383, n64384, n64385, n64386, n64387, n64388, n64389, n64390, n64391, n64392, n64393, n64394, n64395, n64396, n64397, n64398, n64399, n64400, n64401, n64402, n64403, n64404, n64405, n64406, n64407, n64408, n64409, n64410, n64411, n64412, n64413, n64414, n64415, n64416, n64417, n64418, n64419, n64420, n64421, n64422, n64423, n64424, n64425, n64426, n64427, n64428, n64429, n64430, n64431, n64432, n64433, n64434, n64435, n64436, n64437, n64438, n64439, n64440, n64441, n64442, n64443, n64444, n64445, n64446, n64447, n64448, n64449, n64450, n64451, n64452, n64453, n64454, n64455, n64456, n64457, n64458, n64459, n64460, n64461, n64462, n64463, n64464, n64465, n64466, n64467, n64468, n64469, n64470, n64471, n64472, n64473, n64474, n64475, n64476, n64477, n64478, n64479, n64480, n64481, n64482, n64483, n64484, n64485, n64486, n64487, n64488, n64489, n64490, n64491, n64492, n64493, n64494, n64495, n64496, n64497, n64498, n64499, n64500, n64501, n64502, n64503, n64504, n64505, n64506, n64507, n64508, n64509, n64510, n64511, n64512, n64513, n64514, n64515, n64516, n64517, n64518, n64519, n64520, n64521, n64522, n64523, n64524, n64525, n64526, n64527, n64528, n64529, n64530, n64531, n64532, n64533, n64534, n64535, n64536, n64537, n64538, n64539, n64540, n64541, n64542, n64543, n64544, n64545, n64546, n64547, n64548, n64549, n64550, n64551, n64552, n64553, n64554, n64555, n64556, n64557, n64558, n64559, n64560, n64561, n64562, n64563, n64564, n64565, n64566, n64567, n64568, n64569, n64570, n64571, n64572, n64573, n64574, n64575, n64576, n64577, n64578, n64579, n64580, n64581, n64582, n64583, n64584, n64585, n64586, n64587, n64588, n64589, n64590, n64591, n64592, n64593, n64594, n64595, n64596, n64597, n64598, n64599, n64600, n64601, n64602, n64603, n64604, n64605, n64606, n64607, n64608, n64609, n64610, n64611, n64612, n64613, n64614, n64615, n64616, n64617, n64618, n64619, n64620, n64621, n64622, n64623, n64624, n64625, n64626, n64627, n64628, n64629, n64630, n64631, n64632, n64633, n64634, n64635, n64636, n64637, n64638, n64639, n64640, n64641, n64642, n64643, n64644, n64645, n64646, n64647, n64648, n64649, n64650, n64651, n64652, n64653, n64654, n64655, n64656, n64657, n64658, n64659, n64660, n64661, n64662, n64663, n64664, n64665, n64666, n64667, n64668, n64669, n64670, n64671, n64672, n64673, n64674, n64675, n64676, n64677, n64678, n64679, n64680, n64681, n64682, n64683, n64684, n64685, n64686, n64687, n64688, n64689, n64690, n64691, n64692, n64693, n64694, n64695, n64696, n64697, n64698, n64699, n64700, n64701, n64702, n64703, n64704, n64705, n64706, n64707, n64708, n64709, n64710, n64711, n64712, n64713, n64714, n64715, n64716, n64717, n64718, n64719, n64720, n64721, n64722, n64723, n64724, n64725, n64726, n64727, n64728, n64729, n64730, n64731, n64732, n64733, n64734, n64735, n64736, n64737, n64738, n64739, n64740, n64741, n64742, n64743, n64744, n64745, n64746, n64747, n64748, n64749, n64750, n64751, n64752, n64753, n64754, n64755, n64756, n64757, n64758, n64759, n64760, n64761, n64762, n64763, n64764, n64765, n64766, n64767, n64768, n64769, n64770, n64771, n64772, n64773, n64774, n64775, n64776, n64777, n64778, n64779, n64780, n64781, n64782, n64783, n64784, n64785, n64786, n64787, n64788, n64789, n64790, n64791, n64792, n64793, n64794, n64795, n64796, n64797, n64798, n64799, n64800, n64801, n64802, n64803, n64804, n64805, n64806, n64807, n64808, n64809, n64810, n64811, n64812, n64813, n64814, n64815, n64816, n64817, n64818, n64819, n64820, n64821, n64822, n64823, n64824, n64825, n64826, n64827, n64828, n64829, n64830, n64831, n64832, n64833, n64834, n64835, n64836, n64837, n64838, n64839, n64840, n64841, n64842, n64843, n64844, n64845, n64846, n64847, n64848, n64849, n64850, n64851, n64852, n64853, n64854, n64855, n64856, n64857, n64858, n64859, n64860, n64861, n64862, n64863, n64864, n64865, n64866, n64867, n64868, n64869, n64870, n64871, n64872, n64873, n64874, n64875, n64876, n64877, n64878, n64879, n64880, n64881, n64882, n64883, n64884, n64885, n64886, n64887, n64888, n64889, n64890, n64891, n64892, n64893, n64894, n64895, n64896, n64897, n64898, n64899, n64900, n64901, n64902, n64903, n64904, n64905, n64906, n64907, n64908, n64909, n64910, n64911, n64912, n64913, n64914, n64915, n64916, n64917, n64918, n64919, n64920, n64921, n64922, n64923, n64924, n64925, n64926, n64927, n64928, n64929, n64930, n64931, n64932, n64933, n64934, n64935, n64936, n64937, n64938, n64939, n64940, n64941, n64942, n64943, n64944, n64945, n64946, n64947, n64948, n64949, n64950, n64951, n64952, n64953, n64954, n64955, n64956, n64957, n64958, n64959, n64960, n64961, n64962, n64963, n64964, n64965, n64966, n64967, n64968, n64969, n64970, n64971, n64972, n64973, n64974, n64975, n64976, n64977, n64978, n64979, n64980, n64981, n64982, n64983, n64984, n64985, n64986, n64987, n64988, n64989, n64990, n64991, n64992, n64993, n64994, n64995, n64996, n64997, n64998, n64999, n65000, n65001, n65002, n65003, n65004, n65005, n65006, n65007, n65008, n65009, n65010, n65011, n65012, n65013, n65014, n65015, n65016, n65017, n65018, n65019, n65020, n65021, n65022, n65023, n65024, n65025, n65026, n65027, n65028, n65029, n65030, n65031, n65032, n65033, n65034, n65035, n65036, n65037, n65038, n65039, n65040, n65041, n65042, n65043, n65044, n65045, n65046, n65047, n65048, n65049, n65050, n65051, n65052, n65053, n65054, n65055, n65056, n65057, n65058, n65059, n65060, n65061, n65062, n65063, n65064, n65065, n65066, n65067, n65068, n65069, n65070, n65071, n65072, n65073, n65074, n65075, n65076, n65077, n65078, n65079, n65080, n65081, n65082, n65083, n65084, n65085, n65086, n65087, n65088, n65089, n65090, n65091, n65092, n65093, n65094, n65095, n65096, n65097, n65098, n65099, n65100, n65101, n65102, n65103, n65104, n65105, n65106, n65107, n65108, n65109, n65110, n65111, n65112, n65113, n65114, n65115, n65116, n65117, n65118, n65119, n65120, n65121, n65122, n65123, n65124, n65125, n65126, n65127, n65128, n65129, n65130, n65131, n65132, n65133, n65134, n65135, n65136, n65137, n65138, n65139, n65140, n65141, n65142, n65143, n65144, n65145, n65146, n65147, n65148, n65149, n65150, n65151, n65152, n65153, n65154, n65155, n65156, n65157, n65158, n65159, n65160, n65161, n65162, n65163, n65164, n65165, n65166, n65167, n65168, n65169, n65170, n65171, n65172, n65173, n65174, n65175, n65176, n65177, n65178, n65179, n65180, n65181, n65182, n65183, n65184, n65185, n65186, n65187, n65188, n65189, n65190, n65191, n65192, n65193, n65194, n65195, n65196, n65197, n65198, n65199, n65200, n65201, n65202, n65203, n65204, n65205, n65206, n65207, n65208, n65209, n65210, n65211, n65212, n65213, n65214, n65215, n65216, n65217, n65218, n65219, n65220, n65221, n65222, n65223, n65224, n65225, n65226, n65227, n65228, n65229, n65230, n65231, n65232, n65233, n65234, n65235, n65236, n65237, n65238, n65239, n65240, n65241, n65242, n65243, n65244, n65245, n65246, n65247, n65248, n65249, n65250, n65251, n65252, n65253, n65254, n65255, n65256, n65257, n65258, n65259, n65260, n65261, n65262, n65263, n65264, n65265, n65266, n65267, n65268, n65269, n65270, n65271, n65272, n65273, n65274, n65275, n65276, n65277, n65278, n65279, n65280, n65281, n65282, n65283, n65284, n65285, n65286, n65287, n65288, n65289, n65290, n65291, n65292, n65293, n65294, n65295, n65296, n65297, n65298, n65299, n65300, n65301, n65302, n65303, n65304, n65305, n65306, n65307, n65308, n65309, n65310, n65311, n65312, n65313, n65314, n65315, n65316, n65317, n65318, n65319, n65320, n65321, n65322, n65323, n65324, n65325, n65326, n65327, n65328, n65329, n65330, n65331, n65332, n65333, n65334, n65335, n65336, n65337, n65338, n65339, n65340, n65341, n65342, n65343, n65344, n65345, n65346, n65347, n65348, n65349, n65350, n65351, n65352, n65353, n65354, n65355, n65356, n65357, n65358, n65359, n65360, n65361, n65362, n65363, n65364, n65365, n65366, n65367, n65368, n65369, n65370, n65371, n65372, n65373, n65374, n65375, n65376, n65377, n65378, n65379, n65380, n65381, n65382, n65383, n65384, n65385, n65386, n65387, n65388, n65389, n65390, n65391, n65392, n65393, n65394, n65395, n65396, n65397, n65398, n65399, n65400, n65401, n65402, n65403, n65404, n65405, n65406, n65407, n65408, n65409, n65410, n65411, n65412, n65413, n65414, n65415, n65416, n65417, n65418, n65419, n65420, n65421, n65422, n65423, n65424, n65425, n65426, n65427, n65428, n65429, n65430, n65431, n65432, n65433, n65434, n65435, n65436, n65437, n65438, n65439, n65440, n65441, n65442, n65443, n65444, n65445, n65446, n65447, n65448, n65449, n65450, n65451, n65452, n65453, n65454, n65455, n65456, n65457, n65458, n65459, n65460, n65461, n65462, n65463, n65464, n65465, n65466, n65467, n65468, n65469, n65470, n65471, n65472, n65473, n65474, n65475, n65476, n65477, n65478, n65479, n65480, n65481, n65482, n65483, n65484, n65485, n65486, n65487, n65488, n65489, n65490, n65491, n65492, n65493, n65494, n65495, n65496, n65497, n65498, n65499, n65500, n65501, n65502, n65503, n65504, n65505, n65506, n65507, n65508, n65509, n65510, n65511, n65512, n65513, n65514, n65515, n65516, n65517, n65518, n65519, n65520, n65521, n65522, n65523, n65524, n65525, n65526, n65527, n65528, n65529, n65530, n65531, n65532, n65533, n65534, n65535, n65536, n65537, n65538, n65539, n65540, n65541, n65542, n65543, n65544, n65545, n65546, n65547, n65548, n65549, n65550, n65551, n65552, n65553, n65554, n65555, n65556, n65557, n65558, n65559, n65560, n65561, n65562, n65563, n65564, n65565, n65566, n65567, n65568, n65569, n65570, n65571, n65572, n65573, n65574, n65575, n65576, n65577, n65578, n65579, n65580, n65581, n65582, n65583, n65584, n65585, n65586, n65587, n65588, n65589, n65590, n65591, n65592, n65593, n65594, n65595, n65596, n65597, n65598, n65599, n65600, n65601, n65602, n65603, n65604, n65605, n65606, n65607, n65608, n65609, n65610, n65611, n65612, n65613, n65614, n65615, n65616, n65617, n65618, n65619, n65620, n65621, n65622, n65623, n65624, n65625, n65626, n65627, n65628, n65629, n65630, n65631, n65632, n65633, n65634, n65635, n65636, n65637, n65638, n65639, n65640, n65641, n65642, n65643, n65644, n65645, n65646, n65647, n65648, n65649, n65650, n65651, n65652, n65653, n65654, n65655, n65656, n65657, n65658, n65659, n65660, n65661, n65662, n65663, n65664, n65665, n65666, n65667, n65668, n65669, n65670, n65671, n65672, n65673, n65674, n65675, n65676, n65677, n65678, n65679, n65680, n65681, n65682, n65683, n65684, n65685, n65686, n65687, n65688, n65689, n65690, n65691, n65692, n65693, n65694, n65695, n65696, n65697, n65698, n65699, n65700, n65701, n65702, n65703, n65704, n65705, n65706, n65707, n65708, n65709, n65710, n65711, n65712, n65713, n65714, n65715, n65716, n65717, n65718, n65719, n65720, n65721, n65722, n65723, n65724, n65725, n65726, n65727, n65728, n65729, n65730, n65731, n65732, n65733, n65734, n65735, n65736, n65737, n65738, n65739, n65740, n65741, n65742, n65743, n65744, n65745, n65746, n65747, n65748, n65749, n65750, n65751, n65752, n65753, n65754, n65755, n65756, n65757, n65758, n65759, n65760, n65761, n65762, n65763, n65764, n65765, n65766, n65767, n65768, n65769, n65770, n65771, n65772, n65773, n65774, n65775, n65776, n65777, n65778, n65779, n65780, n65781, n65782, n65783, n65784, n65785, n65786, n65787, n65788, n65789, n65790, n65791, n65792, n65793, n65794, n65795, n65796, n65797, n65798, n65799, n65800, n65801, n65802, n65803, n65804, n65805, n65806, n65807, n65808, n65809, n65810, n65811, n65812, n65813, n65814, n65815, n65816, n65817, n65818, n65819, n65820, n65821, n65822, n65823, n65824, n65825, n65826, n65827, n65828, n65829, n65830, n65831, n65832, n65833, n65834, n65835, n65836, n65837, n65838, n65839, n65840, n65841, n65842, n65843, n65844, n65845, n65846, n65847, n65848, n65849, n65850, n65851, n65852, n65853, n65854, n65855, n65856, n65857, n65858, n65859, n65860, n65861, n65862, n65863, n65864, n65865, n65866, n65867, n65868, n65869, n65870, n65871, n65872, n65873, n65874, n65875, n65876, n65877, n65878, n65879, n65880, n65881, n65882, n65883, n65884, n65885, n65886, n65887, n65888, n65889, n65890, n65891, n65892, n65893, n65894, n65895, n65896, n65897, n65898, n65899, n65900, n65901, n65902, n65903, n65904, n65905, n65906, n65907, n65908, n65909, n65910, n65911, n65912, n65913, n65914, n65915, n65916, n65917, n65918, n65919, n65920, n65921, n65922, n65923, n65924, n65925, n65926, n65927, n65928, n65929, n65930, n65931, n65932, n65933, n65934, n65935, n65936, n65937, n65938, n65939, n65940, n65941, n65942, n65943, n65944, n65945, n65946, n65947, n65948, n65949, n65950, n65951, n65952, n65953, n65954, n65955, n65956, n65957, n65958, n65959, n65960, n65961, n65962, n65963, n65964, n65965, n65966, n65967, n65968, n65969, n65970, n65971, n65972, n65973, n65974, n65975, n65976, n65977, n65978, n65979, n65980, n65981, n65982, n65983, n65984, n65985, n65986, n65987, n65988, n65989, n65990, n65991, n65992, n65993, n65994, n65995, n65996, n65997, n65998, n65999, n66000, n66001, n66002, n66003, n66004, n66005, n66006, n66007, n66008, n66009, n66010, n66011, n66012, n66013, n66014, n66015, n66016, n66017, n66018, n66019, n66020, n66021, n66022, n66023, n66024, n66025, n66026, n66027, n66028, n66029, n66030, n66031, n66032, n66033, n66034, n66035, n66036, n66037, n66038, n66039, n66040, n66041, n66042, n66043, n66044, n66045, n66046, n66047, n66048, n66049, n66050, n66051, n66052, n66053, n66054, n66055, n66056, n66057, n66058, n66059, n66060, n66061, n66062, n66063, n66064, n66065, n66066, n66067, n66068, n66069, n66070, n66071, n66072, n66073, n66074, n66075, n66076, n66077, n66078, n66079, n66080, n66081, n66082, n66083, n66084, n66085, n66086, n66087, n66088, n66089, n66090, n66091, n66092, n66093, n66094, n66095, n66096, n66097, n66098, n66099, n66100, n66101, n66102, n66103, n66104, n66105, n66106, n66107, n66108, n66109, n66110, n66111, n66112, n66113, n66114, n66115, n66116, n66117, n66118, n66119, n66120, n66121, n66122, n66123, n66124, n66125, n66126, n66127, n66128, n66129, n66130, n66131, n66132, n66133, n66134, n66135, n66136, n66137, n66138, n66139, n66140, n66141, n66142, n66143, n66144, n66145, n66146, n66147, n66148, n66149, n66150, n66151, n66152, n66153, n66154, n66155, n66156, n66157, n66158, n66159, n66160, n66161, n66162, n66163, n66164, n66165, n66166, n66167, n66168, n66169, n66170, n66171, n66172, n66173, n66174, n66175, n66176, n66177, n66178, n66179, n66180, n66181, n66182, n66183, n66184, n66185, n66186, n66187, n66188, n66189, n66190, n66191, n66192, n66193, n66194, n66195, n66196, n66197, n66198, n66199, n66200, n66201, n66202, n66203, n66204, n66205, n66206, n66207, n66208, n66209, n66210, n66211, n66212, n66213, n66214, n66215, n66216, n66217, n66218, n66219, n66220, n66221, n66222, n66223, n66224, n66225, n66226, n66227, n66228, n66229, n66230, n66231, n66232, n66233, n66234, n66235, n66236, n66237, n66238, n66239, n66240, n66241, n66242, n66243, n66244, n66245, n66246, n66247, n66248, n66249, n66250, n66251, n66252, n66253, n66254, n66255, n66256, n66257, n66258, n66259, n66260, n66261, n66262, n66263, n66264, n66265, n66266, n66267, n66268, n66269, n66270, n66271, n66272, n66273, n66274, n66275, n66276, n66277, n66278, n66279, n66280, n66281, n66282, n66283, n66284, n66285, n66286, n66287, n66288, n66289, n66290, n66291, n66292, n66293, n66294, n66295, n66296, n66297, n66298, n66299, n66300, n66301, n66302, n66303, n66304, n66305, n66306, n66307, n66308, n66309, n66310, n66311, n66312, n66313, n66314, n66315, n66316, n66317, n66318, n66319, n66320, n66321, n66322, n66323, n66324, n66325, n66326, n66327, n66328, n66329, n66330, n66331, n66332, n66333, n66334, n66335, n66336, n66337, n66338, n66339, n66340, n66341, n66342, n66343, n66344, n66345, n66346, n66347, n66348, n66349, n66350, n66351, n66352, n66353, n66354, n66355, n66356, n66357, n66358, n66359, n66360, n66361, n66362, n66363, n66364, n66365, n66366, n66367, n66368, n66369, n66370, n66371, n66372, n66373, n66374, n66375, n66376, n66377, n66378, n66379, n66380, n66381, n66382, n66383, n66384, n66385, n66386, n66387, n66388, n66389, n66390, n66391, n66392, n66393, n66394, n66395, n66396, n66397, n66398, n66399, n66400, n66401, n66402, n66403, n66404, n66405, n66406, n66407, n66408, n66409, n66410, n66411, n66412, n66413, n66414, n66415, n66416, n66417, n66418, n66419, n66420, n66421, n66422, n66423, n66424, n66425, n66426, n66427, n66428, n66429, n66430, n66431, n66432, n66433, n66434, n66435, n66436, n66437, n66438, n66439, n66440, n66441, n66442, n66443, n66444, n66445, n66446, n66447, n66448, n66449, n66450, n66451, n66452, n66453, n66454, n66455, n66456, n66457, n66458, n66459, n66460, n66461, n66462, n66463, n66464, n66465, n66466, n66467, n66468, n66469, n66470, n66471, n66472, n66473, n66474, n66475, n66476, n66477, n66478, n66479, n66480, n66481, n66482, n66483, n66484, n66485, n66486, n66487, n66488, n66489, n66490, n66491, n66492, n66493, n66494, n66495, n66496, n66497, n66498, n66499, n66500, n66501, n66502, n66503, n66504, n66505, n66506, n66507, n66508, n66509, n66510, n66511, n66512, n66513, n66514, n66515, n66516, n66517, n66518, n66519, n66520, n66521, n66522, n66523, n66524, n66525, n66526, n66527, n66528, n66529, n66530, n66531, n66532, n66533, n66534, n66535, n66536, n66537, n66538, n66539, n66540, n66541, n66542, n66543, n66544, n66545, n66546, n66547, n66548, n66549, n66550, n66551, n66552, n66553, n66554, n66555, n66556, n66557, n66558, n66559, n66560, n66561, n66562, n66563, n66564, n66565, n66566, n66567, n66568, n66569, n66570, n66571, n66572, n66573, n66574, n66575, n66576, n66577, n66578, n66579, n66580, n66581, n66582, n66583, n66584, n66585, n66586, n66587, n66588, n66589, n66590, n66591, n66592, n66593, n66594, n66595, n66596, n66597, n66598, n66599, n66600, n66601, n66602, n66603, n66604, n66605, n66606, n66607, n66608, n66609, n66610, n66611, n66612, n66613, n66614, n66615, n66616, n66617, n66618, n66619, n66620, n66621, n66622, n66623, n66624, n66625, n66626, n66627, n66628, n66629, n66630, n66631, n66632, n66633, n66634, n66635, n66636, n66637, n66638, n66639, n66640, n66641, n66642, n66643, n66644, n66645, n66646, n66647, n66648, n66649, n66650, n66651, n66652, n66653, n66654, n66655, n66656, n66657, n66658, n66659, n66660, n66661, n66662, n66663, n66664, n66665, n66666, n66667, n66668, n66669, n66670, n66671, n66672, n66673, n66674, n66675, n66676, n66677, n66678, n66679, n66680, n66681, n66682, n66683, n66684, n66685, n66686, n66687, n66688, n66689, n66690, n66691, n66692, n66693, n66694, n66695, n66696, n66697, n66698, n66699, n66700, n66701, n66702, n66703, n66704, n66705, n66706, n66707, n66708, n66709, n66710, n66711, n66712, n66713, n66714, n66715, n66716, n66717, n66718, n66719, n66720, n66721, n66722, n66723, n66724, n66725, n66726, n66727, n66728, n66729, n66730, n66731, n66732, n66733, n66734, n66735, n66736, n66737, n66738, n66739, n66740, n66741, n66742, n66743, n66744, n66745, n66746, n66747, n66748, n66749, n66750, n66751, n66752, n66753, n66754, n66755, n66756, n66757, n66758, n66759, n66760, n66761, n66762, n66763, n66764, n66765, n66766, n66767, n66768, n66769, n66770, n66771, n66772, n66773, n66774, n66775, n66776, n66777, n66778, n66779, n66780, n66781, n66782, n66783, n66784, n66785, n66786, n66787, n66788, n66789, n66790, n66791, n66792, n66793, n66794, n66795, n66796, n66797, n66798, n66799, n66800, n66801, n66802, n66803, n66804, n66805, n66806, n66807, n66808, n66809, n66810, n66811, n66812, n66813, n66814, n66815, n66816, n66817, n66818, n66819, n66820, n66821, n66822, n66823, n66824, n66825, n66826, n66827, n66828, n66829, n66830, n66831, n66832, n66833, n66834, n66835, n66836, n66837, n66838, n66839, n66840, n66841, n66842, n66843, n66844, n66845, n66846, n66847, n66848, n66849, n66850, n66851, n66852, n66853, n66854, n66855, n66856, n66857, n66858, n66859, n66860, n66861, n66862, n66863, n66864, n66865, n66866, n66867, n66868, n66869, n66870, n66871, n66872, n66873, n66874, n66875, n66876, n66877, n66878, n66879, n66880, n66881, n66882, n66883, n66884, n66885, n66886, n66887, n66888, n66889, n66890, n66891, n66892, n66893, n66894, n66895, n66896, n66897, n66898, n66899, n66900, n66901, n66902, n66903, n66904, n66905, n66906, n66907, n66908, n66909, n66910, n66911, n66912, n66913, n66914, n66915, n66916, n66917, n66918, n66919, n66920, n66921, n66922, n66923, n66924, n66925, n66926, n66927, n66928, n66929, n66930, n66931, n66932, n66933, n66934, n66935, n66936, n66937, n66938, n66939, n66940, n66941, n66942, n66943, n66944, n66945, n66946, n66947, n66948, n66949, n66950, n66951, n66952, n66953, n66954, n66955, n66956, n66957, n66958, n66959, n66960, n66961, n66962, n66963, n66964, n66965, n66966, n66967, n66968, n66969, n66970, n66971, n66972, n66973, n66974, n66975, n66976, n66977, n66978, n66979, n66980, n66981, n66982, n66983, n66984, n66985, n66986, n66987, n66988, n66989, n66990, n66991, n66992, n66993, n66994, n66995, n66996, n66997, n66998, n66999, n67000, n67001, n67002, n67003, n67004, n67005, n67006, n67007, n67008, n67009, n67010, n67011, n67012, n67013, n67014, n67015, n67016, n67017, n67018, n67019, n67020, n67021, n67022, n67023, n67024, n67025, n67026, n67027, n67028, n67029, n67030, n67031, n67032, n67033, n67034, n67035, n67036, n67037, n67038, n67039, n67040, n67041, n67042, n67043, n67044, n67045, n67046, n67047, n67048, n67049, n67050, n67051, n67052, n67053, n67054, n67055, n67056, n67057, n67058, n67059, n67060, n67061, n67062, n67063, n67064, n67065, n67066, n67067, n67068, n67069, n67070, n67071, n67072, n67073, n67074, n67075, n67076, n67077, n67078, n67079, n67080, n67081, n67082, n67083, n67084, n67085, n67086, n67087, n67088, n67089, n67090, n67091, n67092, n67093, n67094, n67095, n67096, n67097, n67098, n67099, n67100, n67101, n67102, n67103, n67104, n67105, n67106, n67107, n67108, n67109, n67110, n67111, n67112, n67113, n67114, n67115, n67116, n67117, n67118, n67119, n67120, n67121, n67122, n67123, n67124, n67125, n67126, n67127, n67128, n67129, n67130, n67131, n67132, n67133, n67134, n67135, n67136, n67137, n67138, n67139, n67140, n67141, n67142, n67143, n67144, n67145, n67146, n67147, n67148, n67149, n67150, n67151, n67152, n67153, n67154, n67155, n67156, n67157, n67158, n67159, n67160, n67161, n67162, n67163, n67164, n67165, n67166, n67167, n67168, n67169, n67170, n67171, n67172, n67173, n67174, n67175, n67176, n67177, n67178, n67179, n67180, n67181, n67182, n67183, n67184, n67185, n67186, n67187, n67188, n67189, n67190, n67191, n67192, n67193, n67194, n67195, n67196, n67197, n67198, n67199, n67200, n67201, n67202, n67203, n67204, n67205, n67206, n67207, n67208, n67209, n67210, n67211, n67212, n67213, n67214, n67215, n67216, n67217, n67218, n67219, n67220, n67221, n67222, n67223, n67224, n67225, n67226, n67227, n67228, n67229, n67230, n67231, n67232, n67233, n67234, n67235, n67236, n67237, n67238, n67239, n67240, n67241, n67242, n67243, n67244, n67245, n67246, n67247, n67248, n67249, n67250, n67251, n67252, n67253, n67254, n67255, n67256, n67257, n67258, n67259, n67260, n67261, n67262, n67263, n67264, n67265, n67266, n67267, n67268, n67269, n67270, n67271, n67272, n67273, n67274, n67275, n67276, n67277, n67278, n67279, n67280, n67281, n67282, n67283, n67284, n67285, n67286, n67287, n67288, n67289, n67290, n67291, n67292, n67293, n67294, n67295, n67296, n67297, n67298, n67299, n67300, n67301, n67302, n67303, n67304, n67305, n67306, n67307, n67308, n67309, n67310, n67311, n67312, n67313, n67314, n67315, n67316, n67317, n67318, n67319, n67320, n67321, n67322, n67323, n67324, n67325, n67326, n67327, n67328, n67329, n67330, n67331, n67332, n67333, n67334, n67335, n67336, n67337, n67338, n67339, n67340, n67341, n67342, n67343, n67344, n67345, n67346, n67347, n67348, n67349, n67350, n67351, n67352, n67353, n67354, n67355, n67356, n67357, n67358, n67359, n67360, n67361, n67362, n67363, n67364, n67365, n67366, n67367, n67368, n67369, n67370, n67371, n67372, n67373, n67374, n67375, n67376, n67377, n67378, n67379, n67380, n67381, n67382, n67383, n67384, n67385, n67386, n67387, n67388, n67389, n67390, n67391, n67392, n67393, n67394, n67395, n67396, n67397, n67398, n67399, n67400, n67401, n67402, n67403, n67404, n67405, n67406, n67407, n67408, n67409, n67410, n67411, n67412, n67413, n67414, n67415, n67416, n67417, n67418, n67419, n67420, n67421, n67422, n67423, n67424, n67425, n67426, n67427, n67428, n67429, n67430, n67431, n67432, n67433, n67434, n67435, n67436, n67437, n67438, n67439, n67440, n67441, n67442, n67443, n67444, n67445, n67446, n67447, n67448, n67449, n67450, n67451, n67452, n67453, n67454, n67455, n67456, n67457, n67458, n67459, n67460, n67461, n67462, n67463, n67464, n67465, n67466, n67467, n67468, n67469, n67470, n67471, n67472, n67473, n67474, n67475, n67476, n67477, n67478, n67479, n67480, n67481, n67482, n67483, n67484, n67485, n67486, n67487, n67488, n67489, n67490, n67491, n67492, n67493, n67494, n67495, n67496, n67497, n67498, n67499, n67500, n67501, n67502, n67503, n67504, n67505, n67506, n67507, n67508, n67509, n67510, n67511, n67512, n67513, n67514, n67515, n67516, n67517, n67518, n67519, n67520, n67521, n67522, n67523, n67524, n67525, n67526, n67527, n67528, n67529, n67530, n67531, n67532, n67533, n67534, n67535, n67536, n67537, n67538, n67539, n67540, n67541, n67542, n67543, n67544, n67545, n67546, n67547, n67548, n67549, n67550, n67551, n67552, n67553, n67554, n67555, n67556, n67557, n67558, n67559, n67560, n67561, n67562, n67563, n67564, n67565, n67566, n67567, n67568, n67569, n67570, n67571, n67572, n67573, n67574, n67575, n67576, n67577, n67578, n67579, n67580, n67581, n67582, n67583, n67584, n67585, n67586, n67587, n67588, n67589, n67590, n67591, n67592, n67593, n67594, n67595, n67596, n67597, n67598, n67599, n67600, n67601, n67602, n67603, n67604, n67605, n67606, n67607, n67608, n67609, n67610, n67611, n67612, n67613, n67614, n67615, n67616, n67617, n67618, n67619, n67620, n67621, n67622, n67623, n67624, n67625, n67626, n67627, n67628, n67629, n67630, n67631, n67632, n67633, n67634, n67635, n67636, n67637, n67638, n67639, n67640, n67641, n67642, n67643, n67644, n67645, n67646, n67647, n67648, n67649, n67650, n67651, n67652, n67653, n67654, n67655, n67656, n67657, n67658, n67659, n67660, n67661, n67662, n67663, n67664, n67665, n67666, n67667, n67668, n67669, n67670, n67671, n67672, n67673, n67674, n67675, n67676, n67677, n67678, n67679, n67680, n67681, n67682, n67683, n67684, n67685, n67686, n67687, n67688, n67689, n67690, n67691, n67692, n67693, n67694, n67695, n67696, n67697, n67698, n67699, n67700, n67701, n67702, n67703, n67704, n67705, n67706, n67707, n67708, n67709, n67710, n67711, n67712, n67713, n67714, n67715, n67716, n67717, n67718, n67719, n67720, n67721, n67722, n67723, n67724, n67725, n67726, n67727, n67728, n67729, n67730, n67731, n67732, n67733, n67734, n67735, n67736, n67737, n67738, n67739, n67740, n67741, n67742, n67743, n67744, n67745, n67746, n67747, n67748, n67749, n67750, n67751, n67752, n67753, n67754, n67755, n67756, n67757, n67758, n67759, n67760, n67761, n67762, n67763, n67764, n67765, n67766, n67767, n67768, n67769, n67770, n67771, n67772, n67773, n67774, n67775, n67776, n67777, n67778, n67779, n67780, n67781, n67782, n67783, n67784, n67785, n67786, n67787, n67788, n67789, n67790, n67791, n67792, n67793, n67794, n67795, n67796, n67797, n67798, n67799, n67800, n67801, n67802, n67803, n67804, n67805, n67806, n67807, n67808, n67809, n67810, n67811, n67812, n67813, n67814, n67815, n67816, n67817, n67818, n67819, n67820, n67821, n67822, n67823, n67824, n67825, n67826, n67827, n67828, n67829, n67830, n67831, n67832, n67833, n67834, n67835, n67836, n67837, n67838, n67839, n67840, n67841, n67842, n67843, n67844, n67845, n67846, n67847, n67848, n67849, n67850, n67851, n67852, n67853, n67854, n67855, n67856, n67857, n67858, n67859, n67860, n67861, n67862, n67863, n67864, n67865, n67866, n67867, n67868, n67869, n67870, n67871, n67872, n67873, n67874, n67875, n67876, n67877, n67878, n67879, n67880, n67881, n67882, n67883, n67884, n67885, n67886, n67887, n67888, n67889, n67890, n67891, n67892, n67893, n67894, n67895, n67896, n67897, n67898, n67899, n67900, n67901, n67902, n67903, n67904, n67905, n67906, n67907, n67908, n67909, n67910, n67911, n67912, n67913, n67914, n67915, n67916, n67917, n67918, n67919, n67920, n67921, n67922, n67923, n67924, n67925, n67926, n67927, n67928, n67929, n67930, n67931, n67932, n67933, n67934, n67935, n67936, n67937, n67938, n67939, n67940, n67941, n67942, n67943, n67944, n67945, n67946, n67947, n67948, n67949, n67950, n67951, n67952, n67953, n67954, n67955, n67956, n67957, n67958, n67959, n67960, n67961, n67962, n67963, n67964, n67965, n67966, n67967, n67968, n67969, n67970, n67971, n67972, n67973, n67974, n67975, n67976, n67977, n67978, n67979, n67980, n67981, n67982, n67983, n67984, n67985, n67986, n67987, n67988, n67989, n67990, n67991, n67992, n67993, n67994, n67995, n67996, n67997, n67998, n67999, n68000, n68001, n68002, n68003, n68004, n68005, n68006, n68007, n68008, n68009, n68010, n68011, n68012, n68013, n68014, n68015, n68016, n68017, n68018, n68019, n68020, n68021, n68022, n68023, n68024, n68025, n68026, n68027, n68028, n68029, n68030, n68031, n68032, n68033, n68034, n68035, n68036, n68037, n68038, n68039, n68040, n68041, n68042, n68043, n68044, n68045, n68046, n68047, n68048, n68049, n68050, n68051, n68052, n68053, n68054, n68055, n68056, n68057, n68058, n68059, n68060, n68061, n68062, n68063, n68064, n68065, n68066, n68067, n68068, n68069, n68070, n68071, n68072, n68073, n68074, n68075, n68076, n68077, n68078, n68079, n68080, n68081, n68082, n68083, n68084, n68085, n68086, n68087, n68088, n68089, n68090, n68091, n68092, n68093, n68094, n68095, n68096, n68097, n68098, n68099, n68100, n68101, n68102, n68103, n68104, n68105, n68106, n68107, n68108, n68109, n68110, n68111, n68112, n68113, n68114, n68115, n68116, n68117, n68118, n68119, n68120, n68121, n68122, n68123, n68124, n68125, n68126, n68127, n68128, n68129, n68130, n68131, n68132, n68133, n68134, n68135, n68136, n68137, n68138, n68139, n68140, n68141, n68142, n68143, n68144, n68145, n68146, n68147, n68148, n68149, n68150, n68151, n68152, n68153, n68154, n68155, n68156, n68157, n68158, n68159, n68160, n68161, n68162, n68163, n68164, n68165, n68166, n68167, n68168, n68169, n68170, n68171, n68172, n68173, n68174, n68175, n68176, n68177, n68178, n68179, n68180, n68181, n68182, n68183, n68184, n68185, n68186, n68187, n68188, n68189, n68190, n68191, n68192, n68193, n68194, n68195, n68196, n68197, n68198, n68199, n68200, n68201, n68202, n68203, n68204, n68205, n68206, n68207, n68208, n68209, n68210, n68211, n68212, n68213, n68214, n68215, n68216, n68217, n68218, n68219, n68220, n68221, n68222, n68223, n68224, n68225, n68226, n68227, n68228, n68229, n68230, n68231, n68232, n68233, n68234, n68235, n68236, n68237, n68238, n68239, n68240, n68241, n68242, n68243, n68244, n68245, n68246, n68247, n68248, n68249, n68250, n68251, n68252, n68253, n68254, n68255, n68256, n68257, n68258, n68259, n68260, n68261, n68262, n68263, n68264, n68265, n68266, n68267, n68268, n68269, n68270, n68271, n68272, n68273, n68274, n68275, n68276, n68277, n68278, n68279, n68280, n68281, n68282, n68283, n68284, n68285, n68286, n68287, n68288, n68289, n68290, n68291, n68292, n68293, n68294, n68295, n68296, n68297, n68298, n68299, n68300, n68301, n68302, n68303, n68304, n68305, n68306, n68307, n68308, n68309, n68310, n68311, n68312, n68313, n68314, n68315, n68316, n68317, n68318, n68319, n68320, n68321, n68322, n68323, n68324, n68325, n68326, n68327, n68328, n68329, n68330, n68331, n68332, n68333, n68334, n68335, n68336, n68337, n68338, n68339, n68340, n68341, n68342, n68343, n68344, n68345, n68346, n68347, n68348, n68349, n68350, n68351, n68352, n68353, n68354, n68355, n68356, n68357, n68358, n68359, n68360, n68361, n68362, n68363, n68364, n68365, n68366, n68367, n68368, n68369, n68370, n68371, n68372, n68373, n68374, n68375, n68376, n68377, n68378, n68379, n68380, n68381, n68382, n68383, n68384, n68385, n68386, n68387, n68388, n68389, n68390, n68391, n68392, n68393, n68394, n68395, n68396, n68397, n68398, n68399, n68400, n68401, n68402, n68403, n68404, n68405, n68406, n68407, n68408, n68409, n68410, n68411, n68412, n68413, n68414, n68415, n68416, n68417, n68418, n68419, n68420, n68421, n68422, n68423, n68424, n68425, n68426, n68427, n68428, n68429, n68430, n68431, n68432, n68433, n68434, n68435, n68436, n68437, n68438, n68439, n68440, n68441, n68442, n68443, n68444, n68445, n68446, n68447, n68448, n68449, n68450, n68451, n68452, n68453, n68454, n68455, n68456, n68457, n68458, n68459, n68460, n68461, n68462, n68463, n68464, n68465, n68466, n68467, n68468, n68469, n68470, n68471, n68472, n68473, n68474, n68475, n68476, n68477, n68478, n68479, n68480, n68481, n68482, n68483, n68484, n68485, n68486, n68487, n68488, n68489, n68490, n68491, n68492, n68493, n68494, n68495, n68496, n68497, n68498, n68499, n68500, n68501, n68502, n68503, n68504, n68505, n68506, n68507, n68508, n68509, n68510, n68511, n68512, n68513, n68514, n68515, n68516, n68517, n68518, n68519, n68520, n68521, n68522, n68523, n68524, n68525, n68526, n68527, n68528, n68529, n68530, n68531, n68532, n68533, n68534, n68535, n68536, n68537, n68538, n68539, n68540, n68541, n68542, n68543, n68544, n68545, n68546, n68547, n68548, n68549, n68550, n68551, n68552, n68553, n68554, n68555, n68556, n68557, n68558, n68559, n68560, n68561, n68562, n68563, n68564, n68565, n68566, n68567, n68568, n68569, n68570, n68571, n68572, n68573, n68574, n68575, n68576, n68577, n68578, n68579, n68580, n68581, n68582, n68583, n68584, n68585, n68586, n68587, n68588, n68589, n68590, n68591, n68592, n68593, n68594, n68595, n68596, n68597, n68598, n68599, n68600, n68601, n68602, n68603, n68604, n68605, n68606, n68607, n68608, n68609, n68610, n68611, n68612, n68613, n68614, n68615, n68616, n68617, n68618, n68619, n68620, n68621, n68622, n68623, n68624, n68625, n68626, n68627, n68628, n68629, n68630, n68631, n68632, n68633, n68634, n68635, n68636, n68637, n68638, n68639, n68640, n68641, n68642, n68643, n68644, n68645, n68646, n68647, n68648, n68649, n68650, n68651, n68652, n68653, n68654, n68655, n68656, n68657, n68658, n68659, n68660, n68661, n68662, n68663, n68664, n68665, n68666, n68667, n68668, n68669, n68670, n68671, n68672, n68673, n68674, n68675, n68676, n68677, n68678, n68679, n68680, n68681, n68682, n68683, n68684, n68685, n68686, n68687, n68688, n68689, n68690, n68691, n68692, n68693, n68694, n68695, n68696, n68697, n68698, n68699, n68700, n68701, n68702, n68703, n68704, n68705, n68706, n68707, n68708, n68709, n68710, n68711, n68712, n68713, n68714, n68715, n68716, n68717, n68718, n68719, n68720, n68721, n68722, n68723, n68724, n68725, n68726, n68727, n68728, n68729, n68730, n68731, n68732, n68733, n68734, n68735, n68736, n68737, n68738, n68739, n68740, n68741, n68742, n68743, n68744, n68745, n68746, n68747, n68748, n68749, n68750, n68751, n68752, n68753, n68754, n68755, n68756, n68757, n68758, n68759, n68760, n68761, n68762, n68763, n68764, n68765, n68766, n68767, n68768, n68769, n68770, n68771, n68772, n68773, n68774, n68775, n68776, n68777, n68778, n68779, n68780, n68781, n68782, n68783, n68784, n68785, n68786, n68787, n68788, n68789, n68790, n68791, n68792, n68793, n68794, n68795, n68796, n68797, n68798, n68799, n68800, n68801, n68802, n68803, n68804, n68805, n68806, n68807, n68808, n68809, n68810, n68811, n68812, n68813, n68814, n68815, n68816, n68817, n68818, n68819, n68820, n68821, n68822, n68823, n68824, n68825, n68826, n68827, n68828, n68829, n68830, n68831, n68832, n68833, n68834, n68835, n68836, n68837, n68838, n68839, n68840, n68841, n68842, n68843, n68844, n68845, n68846, n68847, n68848, n68849, n68850, n68851, n68852, n68853, n68854, n68855, n68856, n68857, n68858, n68859, n68860, n68861, n68862, n68863, n68864, n68865, n68866, n68867, n68868, n68869, n68870, n68871, n68872, n68873, n68874, n68875, n68876, n68877, n68878, n68879, n68880, n68881, n68882, n68883, n68884, n68885, n68886, n68887, n68888, n68889, n68890, n68891, n68892, n68893, n68894, n68895, n68896, n68897, n68898, n68899, n68900, n68901, n68902, n68903, n68904, n68905, n68906, n68907, n68908, n68909, n68910, n68911, n68912, n68913, n68914, n68915, n68916, n68917, n68918, n68919, n68920, n68921, n68922, n68923, n68924, n68925, n68926, n68927, n68928, n68929, n68930, n68931, n68932, n68933, n68934, n68935, n68936, n68937, n68938, n68939, n68940, n68941, n68942, n68943, n68944, n68945, n68946, n68947, n68948, n68949, n68950, n68951, n68952, n68953, n68954, n68955, n68956, n68957, n68958, n68959, n68960, n68961, n68962, n68963, n68964, n68965, n68966, n68967, n68968, n68969, n68970, n68971, n68972, n68973, n68974, n68975, n68976, n68977, n68978, n68979, n68980, n68981, n68982, n68983, n68984, n68985, n68986, n68987, n68988, n68989, n68990, n68991, n68992, n68993, n68994, n68995, n68996, n68997, n68998, n68999, n69000, n69001, n69002, n69003, n69004, n69005, n69006, n69007, n69008, n69009, n69010, n69011, n69012, n69013, n69014, n69015, n69016, n69017, n69018, n69019, n69020, n69021, n69022, n69023, n69024, n69025, n69026, n69027, n69028, n69029, n69030, n69031, n69032, n69033, n69034, n69035, n69036, n69037, n69038, n69039, n69040, n69041, n69042, n69043, n69044, n69045, n69046, n69047, n69048, n69049, n69050, n69051, n69052, n69053, n69054, n69055, n69056, n69057, n69058, n69059, n69060, n69061, n69062, n69063, n69064, n69065, n69066, n69067, n69068, n69069, n69070, n69071, n69072, n69073, n69074, n69075, n69076, n69077, n69078, n69079, n69080, n69081, n69082, n69083, n69084, n69085, n69086, n69087, n69088, n69089, n69090, n69091, n69092, n69093, n69094, n69095, n69096, n69097, n69098, n69099, n69100, n69101, n69102, n69103, n69104, n69105, n69106, n69107, n69108, n69109, n69110, n69111, n69112, n69113, n69114, n69115, n69116, n69117, n69118, n69119, n69120, n69121, n69122, n69123, n69124, n69125, n69126, n69127, n69128, n69129, n69130, n69131, n69132, n69133, n69134, n69135, n69136, n69137, n69138, n69139, n69140, n69141, n69142, n69143, n69144, n69145, n69146, n69147, n69148, n69149, n69150, n69151, n69152, n69153, n69154, n69155, n69156, n69157, n69158, n69159, n69160, n69161, n69162, n69163, n69164, n69165, n69166, n69167, n69168, n69169, n69170, n69171, n69172, n69173, n69174, n69175, n69176, n69177, n69178, n69179, n69180, n69181, n69182, n69183, n69184, n69185, n69186, n69187, n69188, n69189, n69190, n69191, n69192, n69193, n69194, n69195, n69196, n69197, n69198, n69199, n69200, n69201, n69202, n69203, n69204, n69205, n69206, n69207, n69208, n69209, n69210, n69211, n69212, n69213, n69214, n69215, n69216, n69217, n69218, n69219, n69220, n69221, n69222, n69223, n69224, n69225, n69226, n69227, n69228, n69229, n69230, n69231, n69232, n69233, n69234, n69235, n69236, n69237, n69238, n69239, n69240, n69241, n69242, n69243, n69244, n69245, n69246, n69247, n69248, n69249, n69250, n69251, n69252, n69253, n69254, n69255, n69256, n69257, n69258, n69259, n69260, n69261, n69262, n69263, n69264, n69265, n69266, n69267, n69268, n69269, n69270, n69271, n69272, n69273, n69274, n69275, n69276, n69277, n69278, n69279, n69280, n69281, n69282, n69283, n69284, n69285, n69286, n69287, n69288, n69289, n69290, n69291, n69292, n69293, n69294, n69295, n69296, n69297, n69298, n69299, n69300, n69301, n69302, n69303, n69304, n69305, n69306, n69307, n69308, n69309, n69310, n69311, n69312, n69313, n69314, n69315, n69316, n69317, n69318, n69319, n69320, n69321, n69322, n69323, n69324, n69325, n69326, n69327, n69328, n69329, n69330, n69331, n69332, n69333, n69334, n69335, n69336, n69337, n69338, n69339, n69340, n69341, n69342, n69343, n69344, n69345, n69346, n69347, n69348, n69349, n69350, n69351, n69352, n69353, n69354, n69355, n69356, n69357, n69358, n69359, n69360, n69361, n69362, n69363, n69364, n69365, n69366, n69367, n69368, n69369, n69370, n69371, n69372, n69373, n69374, n69375, n69376, n69377, n69378, n69379, n69380, n69381, n69382, n69383, n69384, n69385, n69386, n69387, n69388, n69389, n69390, n69391, n69392, n69393, n69394, n69395, n69396, n69397, n69398, n69399, n69400, n69401, n69402, n69403, n69404, n69405, n69406, n69407, n69408, n69409, n69410, n69411, n69412, n69413, n69414, n69415, n69416, n69417, n69418, n69419, n69420, n69421, n69422, n69423, n69424, n69425, n69426, n69427, n69428, n69429, n69430, n69431, n69432, n69433, n69434, n69435, n69436, n69437, n69438, n69439, n69440, n69441, n69442, n69443, n69444, n69445, n69446, n69447, n69448, n69449, n69450, n69451, n69452, n69453, n69454, n69455, n69456, n69457, n69458, n69459, n69460, n69461, n69462, n69463, n69464, n69465, n69466, n69467, n69468, n69469, n69470, n69471, n69472, n69473, n69474, n69475, n69476, n69477, n69478, n69479, n69480, n69481, n69482, n69483, n69484, n69485, n69486, n69487, n69488, n69489, n69490, n69491, n69492, n69493, n69494, n69495, n69496, n69497, n69498, n69499, n69500, n69501, n69502, n69503, n69504, n69505, n69506, n69507, n69508, n69509, n69510, n69511, n69512, n69513, n69514, n69515, n69516, n69517, n69518, n69519, n69520, n69521, n69522, n69523, n69524, n69525, n69526, n69527, n69528, n69529, n69530, n69531, n69532, n69533, n69534, n69535, n69536, n69537, n69538, n69539, n69540, n69541, n69542, n69543, n69544, n69545, n69546, n69547, n69548, n69549, n69550, n69551, n69552, n69553, n69554, n69555, n69556, n69557, n69558, n69559, n69560, n69561, n69562, n69563, n69564, n69565, n69566, n69567, n69568, n69569, n69570, n69571, n69572, n69573, n69574, n69575, n69576, n69577, n69578, n69579, n69580, n69581, n69582, n69583, n69584, n69585, n69586, n69587, n69588, n69589, n69590, n69591, n69592, n69593, n69594, n69595, n69596, n69597, n69598, n69599, n69600, n69601, n69602, n69603, n69604, n69605, n69606, n69607, n69608, n69609, n69610, n69611, n69612, n69613, n69614, n69615, n69616, n69617, n69618, n69619, n69620, n69621, n69622, n69623, n69624, n69625, n69626, n69627, n69628, n69629, n69630, n69631, n69632, n69633, n69634, n69635, n69636, n69637, n69638, n69639, n69640, n69641, n69642, n69643, n69644, n69645, n69646, n69647, n69648, n69649, n69650, n69651, n69652, n69653, n69654, n69655, n69656, n69657, n69658, n69659, n69660, n69661, n69662, n69663, n69664, n69665, n69666, n69667, n69668, n69669, n69670, n69671, n69672, n69673, n69674, n69675, n69676, n69677, n69678, n69679, n69680, n69681, n69682, n69683, n69684, n69685, n69686, n69687, n69688, n69689, n69690, n69691, n69692, n69693, n69694, n69695, n69696, n69697, n69698, n69699, n69700, n69701, n69702, n69703, n69704, n69705, n69706, n69707, n69708, n69709, n69710, n69711, n69712, n69713, n69714, n69715, n69716, n69717, n69718, n69719, n69720, n69721, n69722, n69723, n69724, n69725, n69726, n69727, n69728, n69729, n69730, n69731, n69732, n69733, n69734, n69735, n69736, n69737, n69738, n69739, n69740, n69741, n69742, n69743, n69744, n69745, n69746, n69747, n69748, n69749, n69750, n69751, n69752, n69753, n69754, n69755, n69756, n69757, n69758, n69759, n69760, n69761, n69762, n69763, n69764, n69765, n69766, n69767, n69768, n69769, n69770, n69771, n69772, n69773, n69774, n69775, n69776, n69777, n69778, n69779, n69780, n69781, n69782, n69783, n69784, n69785, n69786, n69787, n69788, n69789, n69790, n69791, n69792, n69793, n69794, n69795, n69796, n69797, n69798, n69799, n69800, n69801, n69802, n69803, n69804, n69805, n69806, n69807, n69808, n69809, n69810, n69811, n69812, n69813, n69814, n69815, n69816, n69817, n69818, n69819, n69820, n69821, n69822, n69823, n69824, n69825, n69826, n69827, n69828, n69829, n69830, n69831, n69832, n69833, n69834, n69835, n69836, n69837, n69838, n69839, n69840, n69841, n69842, n69843, n69844, n69845, n69846, n69847, n69848, n69849, n69850, n69851, n69852, n69853, n69854, n69855, n69856, n69857, n69858, n69859, n69860, n69861, n69862, n69863, n69864, n69865, n69866, n69867, n69868, n69869, n69870, n69871, n69872, n69873, n69874, n69875, n69876, n69877, n69878, n69879, n69880, n69881, n69882, n69883, n69884, n69885, n69886, n69887, n69888, n69889, n69890, n69891, n69892, n69893, n69894, n69895, n69896, n69897, n69898, n69899, n69900, n69901, n69902, n69903, n69904, n69905, n69906, n69907, n69908, n69909, n69910, n69911, n69912, n69913, n69914, n69915, n69916, n69917, n69918, n69919, n69920, n69921, n69922, n69923, n69924, n69925, n69926, n69927, n69928, n69929, n69930, n69931, n69932, n69933, n69934, n69935, n69936, n69937, n69938, n69939, n69940, n69941, n69942, n69943, n69944, n69945, n69946, n69947, n69948, n69949, n69950, n69951, n69952, n69953, n69954, n69955, n69956, n69957, n69958, n69959, n69960, n69961, n69962, n69963, n69964, n69965, n69966, n69967, n69968, n69969, n69970, n69971, n69972, n69973, n69974, n69975, n69976, n69977, n69978, n69979, n69980, n69981, n69982, n69983, n69984, n69985, n69986, n69987, n69988, n69989, n69990, n69991, n69992, n69993, n69994, n69995, n69996, n69997, n69998, n69999, n70000, n70001, n70002, n70003, n70004, n70005, n70006, n70007, n70008, n70009, n70010, n70011, n70012, n70013, n70014, n70015, n70016, n70017, n70018, n70019, n70020, n70021, n70022, n70023, n70024, n70025, n70026, n70027, n70028, n70029, n70030, n70031, n70032, n70033, n70034, n70035, n70036, n70037, n70038, n70039, n70040, n70041, n70042, n70043, n70044, n70045, n70046, n70047, n70048, n70049, n70050, n70051, n70052, n70053, n70054, n70055, n70056, n70057, n70058, n70059, n70060, n70061, n70062, n70063, n70064, n70065, n70066, n70067, n70068, n70069, n70070, n70071, n70072, n70073, n70074, n70075, n70076, n70077, n70078, n70079, n70080, n70081, n70082, n70083, n70084, n70085, n70086, n70087, n70088, n70089, n70090, n70091, n70092, n70093, n70094, n70095, n70096, n70097, n70098, n70099, n70100, n70101, n70102, n70103, n70104, n70105, n70106, n70107, n70108, n70109, n70110, n70111, n70112, n70113, n70114, n70115, n70116, n70117, n70118, n70119, n70120, n70121, n70122, n70123, n70124, n70125, n70126, n70127, n70128, n70129, n70130, n70131, n70132, n70133, n70134, n70135, n70136, n70137, n70138, n70139, n70140, n70141, n70142, n70143, n70144, n70145, n70146, n70147, n70148, n70149, n70150, n70151, n70152, n70153, n70154, n70155, n70156, n70157, n70158, n70159, n70160, n70161, n70162, n70163, n70164, n70165, n70166, n70167, n70168, n70169, n70170, n70171, n70172, n70173, n70174, n70175, n70176, n70177, n70178, n70179, n70180, n70181, n70182, n70183, n70184, n70185, n70186, n70187, n70188, n70189, n70190, n70191, n70192, n70193, n70194, n70195, n70196, n70197, n70198, n70199, n70200, n70201, n70202, n70203, n70204, n70205, n70206, n70207, n70208, n70209, n70210, n70211, n70212, n70213, n70214, n70215, n70216, n70217, n70218, n70219, n70220, n70221, n70222, n70223, n70224, n70225, n70226, n70227, n70228, n70229, n70230, n70231, n70232, n70233, n70234, n70235, n70236, n70237, n70238, n70239, n70240, n70241, n70242, n70243, n70244, n70245, n70246, n70247, n70248, n70249, n70250, n70251, n70252, n70253, n70254, n70255, n70256, n70257, n70258, n70259, n70260, n70261, n70262, n70263, n70264, n70265, n70266, n70267, n70268, n70269, n70270, n70271, n70272, n70273, n70274, n70275, n70276, n70277, n70278, n70279, n70280, n70281, n70282, n70283, n70284, n70285, n70286, n70287, n70288, n70289, n70290, n70291, n70292, n70293, n70294, n70295, n70296, n70297, n70298, n70299, n70300, n70301, n70302, n70303, n70304, n70305, n70306, n70307, n70308, n70309, n70310, n70311, n70312, n70313, n70314, n70315, n70316, n70317, n70318, n70319, n70320, n70321, n70322, n70323, n70324, n70325, n70326, n70327, n70328, n70329, n70330, n70331, n70332, n70333, n70334, n70335, n70336, n70337, n70338, n70339, n70340, n70341, n70342, n70343, n70344, n70345, n70346, n70347, n70348, n70349, n70350, n70351, n70352, n70353, n70354, n70355, n70356, n70357, n70358, n70359, n70360, n70361, n70362, n70363, n70364, n70365, n70366, n70367, n70368, n70369, n70370, n70371, n70372, n70373, n70374, n70375, n70376, n70377, n70378, n70379, n70380, n70381, n70382, n70383, n70384, n70385, n70386, n70387, n70388, n70389, n70390, n70391, n70392, n70393, n70394, n70395, n70396, n70397, n70398, n70399, n70400, n70401, n70402, n70403, n70404, n70405, n70406, n70407, n70408, n70409, n70410, n70411, n70412, n70413, n70414, n70415, n70416, n70417, n70418, n70419, n70420, n70421, n70422, n70423, n70424, n70425, n70426, n70427, n70428, n70429, n70430, n70431, n70432, n70433, n70434, n70435, n70436, n70437, n70438, n70439, n70440, n70441, n70442, n70443, n70444, n70445, n70446, n70447, n70448, n70449, n70450, n70451, n70452, n70453, n70454, n70455, n70456, n70457, n70458, n70459, n70460, n70461, n70462, n70463, n70464, n70465, n70466, n70467, n70468, n70469, n70470, n70471, n70472, n70473, n70474, n70475, n70476, n70477, n70478, n70479, n70480, n70481, n70482, n70483, n70484, n70485, n70486, n70487, n70488, n70489, n70490, n70491, n70492, n70493, n70494, n70495, n70496, n70497, n70498, n70499, n70500, n70501, n70502, n70503, n70504, n70505, n70506, n70507, n70508, n70509, n70510, n70511, n70512, n70513, n70514, n70515, n70516, n70517, n70518, n70519, n70520, n70521, n70522, n70523, n70524, n70525, n70526, n70527, n70528, n70529, n70530, n70531, n70532, n70533, n70534, n70535, n70536, n70537, n70538, n70539, n70540, n70541, n70542, n70543, n70544, n70545, n70546, n70547, n70548, n70549, n70550, n70551, n70552, n70553, n70554, n70555, n70556, n70557, n70558, n70559, n70560, n70561, n70562, n70563, n70564, n70565, n70566, n70567, n70568, n70569, n70570, n70571, n70572, n70573, n70574, n70575, n70576, n70577, n70578, n70579, n70580, n70581, n70582, n70583, n70584, n70585, n70586, n70587, n70588, n70589, n70590, n70591, n70592, n70593, n70594, n70595, n70596, n70597, n70598, n70599, n70600, n70601, n70602, n70603, n70604, n70605, n70606, n70607, n70608, n70609, n70610, n70611, n70612, n70613, n70614, n70615, n70616, n70617, n70618, n70619, n70620, n70621, n70622, n70623, n70624, n70625, n70626, n70627, n70628, n70629, n70630, n70631, n70632, n70633, n70634, n70635, n70636, n70637, n70638, n70639, n70640, n70641, n70642, n70643, n70644, n70645, n70646, n70647, n70648, n70649, n70650, n70651, n70652, n70653, n70654, n70655, n70656, n70657, n70658, n70659, n70660, n70661, n70662, n70663, n70664, n70665, n70666, n70667, n70668, n70669, n70670, n70671, n70672, n70673, n70674, n70675, n70676, n70677, n70678, n70679, n70680, n70681, n70682, n70683, n70684, n70685, n70686, n70687, n70688, n70689, n70690, n70691, n70692, n70693, n70694, n70695, n70696, n70697, n70698, n70699, n70700, n70701, n70702, n70703, n70704, n70705, n70706, n70707, n70708, n70709, n70710, n70711, n70712, n70713, n70714, n70715, n70716, n70717, n70718, n70719, n70720, n70721, n70722, n70723, n70724, n70725, n70726, n70727, n70728, n70729, n70730, n70731, n70732, n70733, n70734, n70735, n70736, n70737, n70738, n70739, n70740, n70741, n70742, n70743, n70744, n70745, n70746, n70747, n70748, n70749, n70750, n70751, n70752, n70753, n70754, n70755, n70756, n70757, n70758, n70759, n70760, n70761, n70762, n70763, n70764, n70765, n70766, n70767, n70768, n70769, n70770, n70771, n70772, n70773, n70774, n70775, n70776, n70777, n70778, n70779, n70780, n70781, n70782, n70783, n70784, n70785, n70786, n70787, n70788, n70789, n70790, n70791, n70792, n70793, n70794, n70795, n70796, n70797, n70798, n70799, n70800, n70801, n70802, n70803, n70804, n70805, n70806, n70807, n70808, n70809, n70810, n70811, n70812, n70813, n70814, n70815, n70816, n70817, n70818, n70819, n70820, n70821, n70822, n70823, n70824, n70825, n70826, n70827, n70828, n70829, n70830, n70831, n70832, n70833, n70834, n70835, n70836, n70837, n70838, n70839, n70840, n70841, n70842, n70843, n70844, n70845, n70846, n70847, n70848, n70849, n70850, n70851, n70852, n70853, n70854, n70855, n70856, n70857, n70858, n70859, n70860, n70861, n70862, n70863, n70864, n70865, n70866, n70867, n70868, n70869, n70870, n70871, n70872, n70873, n70874, n70875, n70876, n70877, n70878, n70879, n70880, n70881, n70882, n70883, n70884, n70885, n70886, n70887, n70888, n70889, n70890, n70891, n70892, n70893, n70894, n70895, n70896, n70897, n70898, n70899, n70900, n70901, n70902, n70903, n70904, n70905, n70906, n70907, n70908, n70909, n70910, n70911, n70912, n70913, n70914, n70915, n70916, n70917, n70918, n70919, n70920, n70921, n70922, n70923, n70924, n70925, n70926, n70927, n70928, n70929, n70930, n70931, n70932, n70933, n70934, n70935, n70936, n70937, n70938, n70939, n70940, n70941, n70942, n70943, n70944, n70945, n70946, n70947, n70948, n70949, n70950, n70951, n70952, n70953, n70954, n70955, n70956, n70957, n70958, n70959, n70960, n70961, n70962, n70963, n70964, n70965, n70966, n70967, n70968, n70969, n70970, n70971, n70972, n70973, n70974, n70975, n70976, n70977, n70978, n70979, n70980, n70981, n70982, n70983, n70984, n70985, n70986, n70987, n70988, n70989, n70990, n70991, n70992, n70993, n70994, n70995, n70996, n70997, n70998, n70999, n71000, n71001, n71002, n71003, n71004, n71005, n71006, n71007, n71008, n71009, n71010, n71011, n71012, n71013, n71014, n71015, n71016, n71017, n71018, n71019, n71020, n71021, n71022, n71023, n71024, n71025, n71026, n71027, n71028, n71029, n71030, n71031, n71032, n71033, n71034, n71035, n71036, n71037, n71038, n71039, n71040, n71041, n71042, n71043, n71044, n71045, n71046, n71047, n71048, n71049, n71050, n71051, n71052, n71053, n71054, n71055, n71056, n71057, n71058, n71059, n71060, n71061, n71062, n71063, n71064, n71065, n71066, n71067, n71068, n71069, n71070, n71071, n71072, n71073, n71074, n71075, n71076, n71077, n71078, n71079, n71080, n71081, n71082, n71083, n71084, n71085, n71086, n71087, n71088, n71089, n71090, n71091, n71092, n71093, n71094, n71095, n71096, n71097, n71098, n71099, n71100, n71101, n71102, n71103, n71104, n71105, n71106, n71107, n71108, n71109, n71110, n71111, n71112, n71113, n71114, n71115, n71116, n71117, n71118, n71119, n71120, n71121, n71122, n71123, n71124, n71125, n71126, n71127, n71128, n71129, n71130, n71131, n71132, n71133, n71134, n71135, n71136, n71137, n71138, n71139, n71140, n71141, n71142, n71143, n71144, n71145, n71146, n71147, n71148, n71149, n71150, n71151, n71152, n71153, n71154, n71155, n71156, n71157, n71158, n71159, n71160, n71161, n71162, n71163, n71164, n71165, n71166, n71167, n71168, n71169, n71170, n71171, n71172, n71173, n71174, n71175, n71176, n71177, n71178, n71179, n71180, n71181, n71182, n71183, n71184, n71185, n71186, n71187, n71188, n71189, n71190, n71191, n71192, n71193, n71194, n71195, n71196, n71197, n71198, n71199, n71200, n71201, n71202, n71203, n71204, n71205, n71206, n71207, n71208, n71209, n71210, n71211, n71212, n71213, n71214, n71215, n71216, n71217, n71218, n71219, n71220, n71221, n71222, n71223, n71224, n71225, n71226, n71227, n71228, n71229, n71230, n71231, n71232, n71233, n71234, n71235, n71236, n71237, n71238, n71239, n71240, n71241, n71242, n71243, n71244, n71245, n71246, n71247, n71248, n71249, n71250, n71251, n71252, n71253, n71254, n71255, n71256, n71257, n71258, n71259, n71260, n71261, n71262, n71263, n71264, n71265, n71266, n71267, n71268, n71269, n71270, n71271, n71272, n71273, n71274, n71275, n71276, n71277, n71278, n71279, n71280, n71281, n71282, n71283, n71284, n71285, n71286, n71287, n71288, n71289, n71290, n71291, n71292, n71293, n71294, n71295, n71296, n71297, n71298, n71299, n71300, n71301, n71302, n71303, n71304, n71305, n71306, n71307, n71308, n71309, n71310, n71311, n71312, n71313, n71314, n71315, n71316, n71317, n71318, n71319, n71320, n71321, n71322, n71323, n71324, n71325, n71326, n71327, n71328, n71329, n71330, n71331, n71332, n71333, n71334, n71335, n71336, n71337, n71338, n71339, n71340, n71341, n71342, n71343, n71344, n71345, n71346, n71347, n71348, n71349, n71350, n71351, n71352, n71353, n71354, n71355, n71356, n71357, n71358, n71359, n71360, n71361, n71362, n71363, n71364, n71365, n71366, n71367, n71368, n71369, n71370, n71371, n71372, n71373, n71374, n71375, n71376, n71377, n71378, n71379, n71380, n71381, n71382, n71383, n71384, n71385, n71386, n71387, n71388, n71389, n71390, n71391, n71392, n71393, n71394, n71395, n71396, n71397, n71398, n71399, n71400, n71401, n71402, n71403, n71404, n71405, n71406, n71407, n71408, n71409, n71410, n71411, n71412, n71413, n71414, n71415, n71416, n71417, n71418, n71419, n71420, n71421, n71422, n71423, n71424, n71425, n71426, n71427, n71428, n71429, n71430, n71431, n71432, n71433, n71434, n71435, n71436, n71437, n71438, n71439, n71440, n71441, n71442, n71443, n71444, n71445, n71446, n71447, n71448, n71449, n71450, n71451, n71452, n71453, n71454, n71455, n71456, n71457, n71458, n71459, n71460, n71461, n71462, n71463, n71464, n71465, n71466, n71467, n71468, n71469, n71470, n71471, n71472, n71473, n71474, n71475, n71476, n71477, n71478, n71479, n71480, n71481, n71482, n71483, n71484, n71485, n71486, n71487, n71488, n71489, n71490, n71491, n71492, n71493, n71494, n71495, n71496, n71497, n71498, n71499, n71500, n71501, n71502, n71503, n71504, n71505, n71506, n71507, n71508, n71509, n71510, n71511, n71512, n71513, n71514, n71515, n71516, n71517, n71518, n71519, n71520, n71521, n71522, n71523, n71524, n71525, n71526, n71527, n71528, n71529, n71530, n71531, n71532, n71533, n71534, n71535, n71536, n71537, n71538, n71539, n71540, n71541, n71542, n71543, n71544, n71545, n71546, n71547, n71548, n71549, n71550, n71551, n71552, n71553, n71554, n71555, n71556, n71557, n71558, n71559, n71560, n71561, n71562, n71563, n71564, n71565, n71566, n71567, n71568, n71569, n71570, n71571, n71572, n71573, n71574, n71575, n71576, n71577, n71578, n71579, n71580, n71581, n71582, n71583, n71584, n71585, n71586, n71587, n71588, n71589, n71590, n71591, n71592, n71593, n71594, n71595, n71596, n71597, n71598, n71599, n71600, n71601, n71602, n71603, n71604, n71605, n71606, n71607, n71608, n71609, n71610, n71611, n71612, n71613, n71614, n71615, n71616, n71617, n71618, n71619, n71620, n71621, n71622, n71623, n71624, n71625, n71626, n71627, n71628, n71629, n71630, n71631, n71632, n71633, n71634, n71635, n71636, n71637, n71638, n71639, n71640, n71641, n71642, n71643, n71644, n71645, n71646, n71647, n71648, n71649, n71650, n71651, n71652, n71653, n71654, n71655, n71656, n71657, n71658, n71659, n71660, n71661, n71662, n71663, n71664, n71665, n71666, n71667, n71668, n71669, n71670, n71671, n71672, n71673, n71674, n71675, n71676, n71677, n71678, n71679, n71680, n71681, n71682, n71683, n71684, n71685, n71686, n71687, n71688, n71689, n71690, n71691, n71692, n71693, n71694, n71695, n71696, n71697, n71698, n71699, n71700, n71701, n71702, n71703, n71704, n71705, n71706, n71707, n71708, n71709, n71710, n71711, n71712, n71713, n71714, n71715, n71716, n71717, n71718, n71719, n71720, n71721, n71722, n71723, n71724, n71725, n71726, n71727, n71728, n71729, n71730, n71731, n71732, n71733, n71734, n71735, n71736, n71737, n71738, n71739, n71740, n71741, n71742, n71743, n71744, n71745, n71746, n71747, n71748, n71749, n71750, n71751, n71752, n71753, n71754, n71755, n71756, n71757, n71758, n71759, n71760, n71761, n71762, n71763, n71764, n71765, n71766, n71767, n71768, n71769, n71770, n71771, n71772, n71773, n71774, n71775, n71776, n71777, n71778, n71779, n71780, n71781, n71782, n71783, n71784, n71785, n71786, n71787, n71788, n71789, n71790, n71791, n71792, n71793, n71794, n71795, n71796, n71797, n71798, n71799, n71800, n71801, n71802, n71803, n71804, n71805, n71806, n71807, n71808, n71809, n71810, n71811, n71812, n71813, n71814, n71815, n71816, n71817, n71818, n71819, n71820, n71821, n71822, n71823, n71824, n71825, n71826, n71827, n71828, n71829, n71830, n71831, n71832, n71833, n71834, n71835, n71836, n71837, n71838, n71839, n71840, n71841, n71842, n71843, n71844, n71845, n71846, n71847, n71848, n71849, n71850, n71851, n71852, n71853, n71854, n71855, n71856, n71857, n71858, n71859, n71860, n71861, n71862, n71863, n71864, n71865, n71866, n71867, n71868, n71869, n71870, n71871, n71872, n71873, n71874, n71875, n71876, n71877, n71878, n71879, n71880, n71881, n71882, n71883, n71884, n71885, n71886, n71887, n71888, n71889, n71890, n71891, n71892, n71893, n71894, n71895, n71896, n71897, n71898, n71899, n71900, n71901, n71902, n71903, n71904, n71905, n71906, n71907, n71908, n71909, n71910, n71911, n71912, n71913, n71914, n71915, n71916, n71917, n71918, n71919, n71920, n71921, n71922, n71923, n71924, n71925, n71926, n71927, n71928, n71929, n71930, n71931, n71932, n71933, n71934, n71935, n71936, n71937, n71938, n71939, n71940, n71941, n71942, n71943, n71944, n71945, n71946, n71947, n71948, n71949, n71950, n71951, n71952, n71953, n71954, n71955, n71956, n71957, n71958, n71959, n71960, n71961, n71962, n71963, n71964, n71965, n71966, n71967, n71968, n71969, n71970, n71971, n71972, n71973, n71974, n71975, n71976, n71977, n71978, n71979, n71980, n71981, n71982, n71983, n71984, n71985, n71986, n71987, n71988, n71989, n71990, n71991, n71992, n71993, n71994, n71995, n71996, n71997, n71998, n71999, n72000, n72001, n72002, n72003, n72004, n72005, n72006, n72007, n72008, n72009, n72010, n72011, n72012, n72013, n72014, n72015, n72016, n72017, n72018, n72019, n72020, n72021, n72022, n72023, n72024, n72025, n72026, n72027, n72028, n72029, n72030, n72031, n72032, n72033, n72034, n72035, n72036, n72037, n72038, n72039, n72040, n72041, n72042, n72043, n72044, n72045, n72046, n72047, n72048, n72049, n72050, n72051, n72052, n72053, n72054, n72055, n72056, n72057, n72058, n72059, n72060, n72061, n72062, n72063, n72064, n72065, n72066, n72067, n72068, n72069, n72070, n72071, n72072, n72073, n72074, n72075, n72076, n72077, n72078, n72079, n72080, n72081, n72082, n72083, n72084, n72085, n72086, n72087, n72088, n72089, n72090, n72091, n72092, n72093, n72094, n72095, n72096, n72097, n72098, n72099, n72100, n72101, n72102, n72103, n72104, n72105, n72106, n72107, n72108, n72109, n72110, n72111, n72112, n72113, n72114, n72115, n72116, n72117, n72118, n72119, n72120, n72121, n72122, n72123, n72124, n72125, n72126, n72127, n72128, n72129, n72130, n72131, n72132, n72133, n72134, n72135, n72136, n72137, n72138, n72139, n72140, n72141, n72142, n72143, n72144, n72145, n72146, n72147, n72148, n72149, n72150, n72151, n72152, n72153, n72154, n72155, n72156, n72157, n72158, n72159, n72160, n72161, n72162, n72163, n72164, n72165, n72166, n72167, n72168, n72169, n72170, n72171, n72172, n72173, n72174, n72175, n72176, n72177, n72178, n72179, n72180, n72181, n72182, n72183, n72184, n72185, n72186, n72187, n72188, n72189, n72190, n72191, n72192, n72193, n72194, n72195, n72196, n72197, n72198, n72199, n72200, n72201, n72202, n72203, n72204, n72205, n72206, n72207, n72208, n72209, n72210, n72211, n72212, n72213, n72214, n72215, n72216, n72217, n72218, n72219, n72220, n72221, n72222, n72223, n72224, n72225, n72226, n72227, n72228, n72229, n72230, n72231, n72232, n72233, n72234, n72235, n72236, n72237, n72238, n72239, n72240, n72241, n72242, n72243, n72244, n72245, n72246, n72247, n72248, n72249, n72250, n72251, n72252, n72253, n72254, n72255, n72256, n72257, n72258, n72259, n72260, n72261, n72262, n72263, n72264, n72265, n72266, n72267, n72268, n72269, n72270, n72271, n72272, n72273, n72274, n72275, n72276, n72277, n72278, n72279, n72280, n72281, n72282, n72283, n72284, n72285, n72286, n72287, n72288, n72289, n72290, n72291, n72292, n72293, n72294, n72295, n72296, n72297, n72298, n72299, n72300, n72301, n72302, n72303, n72304, n72305, n72306, n72307, n72308, n72309, n72310, n72311, n72312, n72313, n72314, n72315, n72316, n72317, n72318, n72319, n72320, n72321, n72322, n72323, n72324, n72325, n72326, n72327, n72328, n72329, n72330, n72331, n72332, n72333, n72334, n72335, n72336, n72337, n72338, n72339, n72340, n72341, n72342, n72343, n72344, n72345, n72346, n72347, n72348, n72349, n72350, n72351, n72352, n72353, n72354, n72355, n72356, n72357, n72358, n72359, n72360, n72361, n72362, n72363, n72364, n72365, n72366, n72367, n72368, n72369, n72370, n72371, n72372, n72373, n72374, n72375, n72376, n72377, n72378, n72379, n72380, n72381, n72382, n72383, n72384, n72385, n72386, n72387, n72388, n72389, n72390, n72391, n72392, n72393, n72394, n72395, n72396, n72397, n72398, n72399, n72400, n72401, n72402, n72403, n72404, n72405, n72406, n72407, n72408, n72409, n72410, n72411, n72412, n72413, n72414, n72415, n72416, n72417, n72418, n72419, n72420, n72421, n72422, n72423, n72424, n72425, n72426, n72427, n72428, n72429, n72430, n72431, n72432, n72433, n72434, n72435, n72436, n72437, n72438, n72439, n72440, n72441, n72442, n72443, n72444, n72445, n72446, n72447, n72448, n72449, n72450, n72451, n72452, n72453, n72454, n72455, n72456, n72457, n72458, n72459, n72460, n72461, n72462, n72463, n72464, n72465, n72466, n72467, n72468, n72469, n72470, n72471, n72472, n72473, n72474, n72475, n72476, n72477, n72478, n72479, n72480, n72481, n72482, n72483, n72484, n72485, n72486, n72487, n72488, n72489, n72490, n72491, n72492, n72493, n72494, n72495, n72496, n72497, n72498, n72499, n72500, n72501, n72502, n72503, n72504, n72505, n72506, n72507, n72508, n72509, n72510, n72511, n72512, n72513, n72514, n72515, n72516, n72517, n72518, n72519, n72520, n72521, n72522, n72523, n72524, n72525, n72526, n72527, n72528, n72529, n72530, n72531, n72532, n72533, n72534, n72535, n72536, n72537, n72538, n72539, n72540, n72541, n72542, n72543, n72544, n72545, n72546, n72547, n72548, n72549, n72550, n72551, n72552, n72553, n72554, n72555, n72556, n72557, n72558, n72559, n72560, n72561, n72562, n72563, n72564, n72565, n72566, n72567, n72568, n72569, n72570, n72571, n72572, n72573, n72574, n72575, n72576, n72577, n72578, n72579, n72580, n72581, n72582, n72583, n72584, n72585, n72586, n72587, n72588, n72589, n72590, n72591, n72592, n72593, n72594, n72595, n72596, n72597, n72598, n72599, n72600, n72601, n72602, n72603, n72604, n72605, n72606, n72607, n72608, n72609, n72610, n72611, n72612, n72613, n72614, n72615, n72616, n72617, n72618, n72619, n72620, n72621, n72622, n72623, n72624, n72625, n72626, n72627, n72628, n72629, n72630, n72631, n72632, n72633, n72634, n72635, n72636, n72637, n72638, n72639, n72640, n72641, n72642, n72643, n72644, n72645, n72646, n72647, n72648, n72649, n72650, n72651, n72652, n72653, n72654, n72655, n72656, n72657, n72658, n72659, n72660, n72661, n72662, n72663, n72664, n72665, n72666, n72667, n72668, n72669, n72670, n72671, n72672, n72673, n72674, n72675, n72676, n72677, n72678, n72679, n72680, n72681, n72682, n72683, n72684, n72685, n72686, n72687, n72688, n72689, n72690, n72691, n72692, n72693, n72694, n72695, n72696, n72697, n72698, n72699, n72700, n72701, n72702, n72703, n72704, n72705, n72706, n72707, n72708, n72709, n72710, n72711, n72712, n72713, n72714, n72715, n72716, n72717, n72718, n72719, n72720, n72721, n72722, n72723, n72724, n72725, n72726, n72727, n72728, n72729, n72730, n72731, n72732, n72733, n72734, n72735, n72736, n72737, n72738, n72739, n72740, n72741, n72742, n72743, n72744, n72745, n72746, n72747, n72748, n72749, n72750, n72751, n72752, n72753, n72754, n72755, n72756, n72757, n72758, n72759, n72760, n72761, n72762, n72763, n72764, n72765, n72766, n72767, n72768, n72769, n72770, n72771, n72772, n72773, n72774, n72775, n72776, n72777, n72778, n72779, n72780, n72781, n72782, n72783, n72784, n72785, n72786, n72787, n72788, n72789, n72790, n72791, n72792, n72793, n72794, n72795, n72796, n72797, n72798, n72799, n72800, n72801, n72802, n72803, n72804, n72805, n72806, n72807, n72808, n72809, n72810, n72811, n72812, n72813, n72814, n72815, n72816, n72817, n72818, n72819, n72820, n72821, n72822, n72823, n72824, n72825, n72826, n72827, n72828, n72829, n72830, n72831, n72832, n72833, n72834, n72835, n72836, n72837, n72838, n72839, n72840, n72841, n72842, n72843, n72844, n72845, n72846, n72847, n72848, n72849, n72850, n72851, n72852, n72853, n72854, n72855, n72856, n72857, n72858, n72859, n72860, n72861, n72862, n72863, n72864, n72865, n72866, n72867, n72868, n72869, n72870, n72871, n72872, n72873, n72874, n72875, n72876, n72877, n72878, n72879, n72880, n72881, n72882, n72883, n72884, n72885, n72886, n72887, n72888, n72889, n72890, n72891, n72892, n72893, n72894, n72895, n72896, n72897, n72898, n72899, n72900, n72901, n72902, n72903, n72904, n72905, n72906, n72907, n72908, n72909, n72910, n72911, n72912, n72913, n72914, n72915, n72916, n72917, n72918, n72919, n72920, n72921, n72922, n72923, n72924, n72925, n72926, n72927, n72928, n72929, n72930, n72931, n72932, n72933, n72934, n72935, n72936, n72937, n72938, n72939, n72940, n72941, n72942, n72943, n72944, n72945, n72946, n72947, n72948, n72949, n72950, n72951, n72952, n72953, n72954, n72955, n72956, n72957, n72958, n72959, n72960, n72961, n72962, n72963, n72964, n72965, n72966, n72967, n72968, n72969, n72970, n72971, n72972, n72973, n72974, n72975, n72976, n72977, n72978, n72979, n72980, n72981, n72982, n72983, n72984, n72985, n72986, n72987, n72988, n72989, n72990, n72991, n72992, n72993, n72994, n72995, n72996, n72997, n72998, n72999, n73000, n73001, n73002, n73003, n73004, n73005, n73006, n73007, n73008, n73009, n73010, n73011, n73012, n73013, n73014, n73015, n73016, n73017, n73018, n73019, n73020, n73021, n73022, n73023, n73024, n73025, n73026, n73027, n73028, n73029, n73030, n73031, n73032, n73033, n73034, n73035, n73036, n73037, n73038, n73039, n73040, n73041, n73042, n73043, n73044, n73045, n73046, n73047, n73048, n73049, n73050, n73051, n73052, n73053, n73054, n73055, n73056, n73057, n73058, n73059, n73060, n73061, n73062, n73063, n73064, n73065, n73066, n73067, n73068, n73069, n73070, n73071, n73072, n73073, n73074, n73075, n73076, n73077, n73078, n73079, n73080, n73081, n73082, n73083, n73084, n73085, n73086, n73087, n73088, n73089, n73090, n73091, n73092, n73093, n73094, n73095, n73096, n73097, n73098, n73099, n73100, n73101, n73102, n73103, n73104, n73105, n73106, n73107, n73108, n73109, n73110, n73111, n73112, n73113, n73114, n73115, n73116, n73117, n73118, n73119, n73120, n73121, n73122, n73123, n73124, n73125, n73126, n73127, n73128, n73129, n73130, n73131, n73132, n73133, n73134, n73135, n73136, n73137, n73138, n73139, n73140, n73141, n73142, n73143, n73144, n73145, n73146, n73147, n73148, n73149, n73150, n73151, n73152, n73153, n73154, n73155, n73156, n73157, n73158, n73159, n73160, n73161, n73162, n73163, n73164, n73165, n73166, n73167, n73168, n73169, n73170, n73171, n73172, n73173, n73174, n73175, n73176, n73177, n73178, n73179, n73180, n73181, n73182, n73183, n73184, n73185, n73186, n73187, n73188, n73189, n73190, n73191, n73192, n73193, n73194, n73195, n73196, n73197, n73198, n73199, n73200, n73201, n73202, n73203, n73204, n73205, n73206, n73207, n73208, n73209, n73210, n73211, n73212, n73213, n73214, n73215, n73216, n73217, n73218, n73219, n73220, n73221, n73222, n73223, n73224, n73225, n73226, n73227, n73228, n73229, n73230, n73231, n73232, n73233, n73234, n73235, n73236, n73237, n73238, n73239, n73240, n73241, n73242, n73243, n73244, n73245, n73246, n73247, n73248, n73249, n73250, n73251, n73252, n73253, n73254, n73255, n73256, n73257, n73258, n73259, n73260, n73261, n73262, n73263, n73264, n73265, n73266, n73267, n73268, n73269, n73270, n73271, n73272, n73273, n73274, n73275, n73276, n73277, n73278, n73279, n73280, n73281, n73282, n73283, n73284, n73285, n73286, n73287, n73288, n73289, n73290, n73291, n73292, n73293, n73294, n73295, n73296, n73297, n73298, n73299, n73300, n73301, n73302, n73303, n73304, n73305, n73306, n73307, n73308, n73309, n73310, n73311, n73312, n73313, n73314, n73315, n73316, n73317, n73318, n73319, n73320, n73321, n73322, n73323, n73324, n73325, n73326, n73327, n73328, n73329, n73330, n73331, n73332, n73333, n73334, n73335, n73336, n73337, n73338, n73339, n73340, n73341, n73342, n73343, n73344, n73345, n73346, n73347, n73348, n73349, n73350, n73351, n73352, n73353, n73354, n73355, n73356, n73357, n73358, n73359, n73360, n73361, n73362, n73363, n73364, n73365, n73366, n73367, n73368, n73369, n73370, n73371, n73372, n73373, n73374, n73375, n73376, n73377, n73378, n73379, n73380, n73381, n73382, n73383, n73384, n73385, n73386, n73387, n73388, n73389, n73390, n73391, n73392, n73393, n73394, n73395, n73396, n73397, n73398, n73399, n73400, n73401, n73402, n73403, n73404, n73405, n73406, n73407, n73408, n73409, n73410, n73411, n73412, n73413, n73414, n73415, n73416, n73417, n73418, n73419, n73420, n73421, n73422, n73423, n73424, n73425, n73426, n73427, n73428, n73429, n73430, n73431, n73432, n73433, n73434, n73435, n73436, n73437, n73438, n73439, n73440, n73441, n73442, n73443, n73444, n73445, n73446, n73447, n73448, n73449, n73450, n73451, n73452, n73453, n73454, n73455, n73456, n73457, n73458, n73459, n73460, n73461, n73462, n73463, n73464, n73465, n73466, n73467, n73468, n73469, n73470, n73471, n73472, n73473, n73474, n73475, n73476, n73477, n73478, n73479, n73480, n73481, n73482, n73483, n73484, n73485, n73486, n73487, n73488, n73489, n73490, n73491, n73492, n73493, n73494, n73495, n73496, n73497, n73498, n73499, n73500, n73501, n73502, n73503, n73504, n73505, n73506, n73507, n73508, n73509, n73510, n73511, n73512, n73513, n73514, n73515, n73516, n73517, n73518, n73519, n73520, n73521, n73522, n73523, n73524, n73525, n73526, n73527, n73528, n73529, n73530, n73531, n73532, n73533, n73534, n73535, n73536, n73537, n73538, n73539, n73540, n73541, n73542, n73543, n73544, n73545, n73546, n73547, n73548, n73549, n73550, n73551, n73552, n73553, n73554, n73555, n73556, n73557, n73558, n73559, n73560, n73561, n73562, n73563, n73564, n73565, n73566, n73567, n73568, n73569, n73570, n73571, n73572, n73573, n73574, n73575, n73576, n73577, n73578, n73579, n73580, n73581, n73582, n73583, n73584, n73585, n73586, n73587, n73588, n73589, n73590, n73591, n73592, n73593, n73594, n73595, n73596, n73597, n73598, n73599, n73600, n73601, n73602, n73603, n73604, n73605, n73606, n73607, n73608, n73609, n73610, n73611, n73612, n73613, n73614, n73615, n73616, n73617, n73618, n73619, n73620, n73621, n73622, n73623, n73624, n73625, n73626, n73627, n73628, n73629, n73630, n73631, n73632, n73633, n73634, n73635, n73636, n73637, n73638, n73639, n73640, n73641, n73642, n73643, n73644, n73645, n73646, n73647, n73648, n73649, n73650, n73651, n73652, n73653, n73654, n73655, n73656, n73657, n73658, n73659, n73660, n73661, n73662, n73663, n73664, n73665, n73666, n73667, n73668, n73669, n73670, n73671, n73672, n73673, n73674, n73675, n73676, n73677, n73678, n73679, n73680, n73681, n73682, n73683, n73684, n73685, n73686, n73687, n73688, n73689, n73690, n73691, n73692, n73693, n73694, n73695, n73696, n73697, n73698, n73699, n73700, n73701, n73702, n73703, n73704, n73705, n73706, n73707, n73708, n73709, n73710, n73711, n73712, n73713, n73714, n73715, n73716, n73717, n73718, n73719, n73720, n73721, n73722, n73723, n73724, n73725, n73726, n73727, n73728, n73729, n73730, n73731, n73732, n73733, n73734, n73735, n73736, n73737, n73738, n73739, n73740, n73741, n73742, n73743, n73744, n73745, n73746, n73747, n73748, n73749, n73750, n73751, n73752, n73753, n73754, n73755, n73756, n73757, n73758, n73759, n73760, n73761, n73762, n73763, n73764, n73765, n73766, n73767, n73768, n73769, n73770, n73771, n73772, n73773, n73774, n73775, n73776, n73777, n73778, n73779, n73780, n73781, n73782, n73783, n73784, n73785, n73786, n73787, n73788, n73789, n73790, n73791, n73792, n73793, n73794, n73795, n73796, n73797, n73798, n73799, n73800, n73801, n73802, n73803, n73804, n73805, n73806, n73807, n73808, n73809, n73810, n73811, n73812, n73813, n73814, n73815, n73816, n73817, n73818, n73819, n73820, n73821, n73822, n73823, n73824, n73825, n73826, n73827, n73828, n73829, n73830, n73831, n73832, n73833, n73834, n73835, n73836, n73837, n73838, n73839, n73840, n73841, n73842, n73843, n73844, n73845, n73846, n73847, n73848, n73849, n73850, n73851, n73852, n73853, n73854, n73855, n73856, n73857, n73858, n73859, n73860, n73861, n73862, n73863, n73864, n73865, n73866, n73867, n73868, n73869, n73870, n73871, n73872, n73873, n73874, n73875, n73876, n73877, n73878, n73879, n73880, n73881, n73882, n73883, n73884, n73885, n73886, n73887, n73888, n73889, n73890, n73891, n73892, n73893, n73894, n73895, n73896, n73897, n73898, n73899, n73900, n73901, n73902, n73903, n73904, n73905, n73906, n73907, n73908, n73909, n73910, n73911, n73912, n73913, n73914, n73915, n73916, n73917, n73918, n73919, n73920, n73921, n73922, n73923, n73924, n73925, n73926, n73927, n73928, n73929, n73930, n73931, n73932, n73933, n73934, n73935, n73936, n73937, n73938, n73939, n73940, n73941, n73942, n73943, n73944, n73945, n73946, n73947, n73948, n73949, n73950, n73951, n73952, n73953, n73954, n73955, n73956, n73957, n73958, n73959, n73960, n73961, n73962, n73963, n73964, n73965, n73966, n73967, n73968, n73969, n73970, n73971, n73972, n73973, n73974, n73975, n73976, n73977, n73978, n73979, n73980, n73981, n73982, n73983, n73984, n73985, n73986, n73987, n73988, n73989, n73990, n73991, n73992, n73993, n73994, n73995, n73996, n73997, n73998, n73999, n74000, n74001, n74002, n74003, n74004, n74005, n74006, n74007, n74008, n74009, n74010, n74011, n74012, n74013, n74014, n74015, n74016, n74017, n74018, n74019, n74020, n74021, n74022, n74023, n74024, n74025, n74026, n74027, n74028, n74029, n74030, n74031, n74032, n74033, n74034, n74035, n74036, n74037, n74038, n74039, n74040, n74041, n74042, n74043, n74044, n74045, n74046, n74047, n74048, n74049, n74050, n74051, n74052, n74053, n74054, n74055, n74056, n74057, n74058, n74059, n74060, n74061, n74062, n74063, n74064, n74065, n74066, n74067, n74068, n74069, n74070, n74071, n74072, n74073, n74074, n74075, n74076, n74077, n74078, n74079, n74080, n74081, n74082, n74083, n74084, n74085, n74086, n74087, n74088, n74089, n74090, n74091, n74092, n74093, n74094, n74095, n74096, n74097, n74098, n74099, n74100, n74101, n74102, n74103, n74104, n74105, n74106, n74107, n74108, n74109, n74110, n74111, n74112, n74113, n74114, n74115, n74116, n74117, n74118, n74119, n74120, n74121, n74122, n74123, n74124, n74125, n74126, n74127, n74128, n74129, n74130, n74131, n74132, n74133, n74134, n74135, n74136, n74137, n74138, n74139, n74140, n74141, n74142, n74143, n74144, n74145, n74146, n74147, n74148, n74149, n74150, n74151, n74152, n74153, n74154, n74155, n74156, n74157, n74158, n74159, n74160, n74161, n74162, n74163, n74164, n74165, n74166, n74167, n74168, n74169, n74170, n74171, n74172, n74173, n74174, n74175, n74176, n74177, n74178, n74179, n74180, n74181, n74182, n74183, n74184, n74185, n74186, n74187, n74188, n74189, n74190, n74191, n74192, n74193, n74194, n74195, n74196, n74197, n74198, n74199, n74200, n74201, n74202, n74203, n74204, n74205, n74206, n74207, n74208, n74209, n74210, n74211, n74212, n74213, n74214, n74215, n74216, n74217, n74218, n74219, n74220, n74221, n74222, n74223, n74224, n74225, n74226, n74227, n74228, n74229, n74230, n74231, n74232, n74233, n74234, n74235, n74236, n74237, n74238, n74239, n74240, n74241, n74242, n74243, n74244, n74245, n74246, n74247, n74248, n74249, n74250, n74251, n74252, n74253, n74254, n74255, n74256, n74257, n74258, n74259, n74260, n74261, n74262, n74263, n74264, n74265, n74266, n74267, n74268, n74269, n74270, n74271, n74272, n74273, n74274, n74275, n74276, n74277, n74278, n74279, n74280, n74281, n74282, n74283, n74284, n74285, n74286, n74287, n74288, n74289, n74290, n74291, n74292, n74293, n74294, n74295, n74296, n74297, n74298, n74299, n74300, n74301, n74302, n74303, n74304, n74305, n74306, n74307, n74308, n74309, n74310, n74311, n74312, n74313, n74314, n74315, n74316, n74317, n74318, n74319, n74320, n74321, n74322, n74323, n74324, n74325, n74326, n74327, n74328, n74329, n74330, n74331, n74332, n74333, n74334, n74335, n74336, n74337, n74338, n74339, n74340, n74341, n74342, n74343, n74344, n74345, n74346, n74347, n74348, n74349, n74350, n74351, n74352, n74353, n74354, n74355, n74356, n74357, n74358, n74359, n74360, n74361, n74362, n74363, n74364, n74365, n74366, n74367, n74368, n74369, n74370, n74371, n74372, n74373, n74374, n74375, n74376, n74377, n74378, n74379, n74380, n74381, n74382, n74383, n74384, n74385, n74386, n74387, n74388, n74389, n74390, n74391, n74392, n74393, n74394, n74395, n74396, n74397, n74398, n74399, n74400, n74401, n74402, n74403, n74404, n74405, n74406, n74407, n74408, n74409, n74410, n74411, n74412, n74413, n74414, n74415, n74416, n74417, n74418, n74419, n74420, n74421, n74422, n74423, n74424, n74425, n74426, n74427, n74428, n74429, n74430, n74431, n74432, n74433, n74434, n74435, n74436, n74437, n74438, n74439, n74440, n74441, n74442, n74443, n74444, n74445, n74446, n74447, n74448, n74449, n74450, n74451, n74452, n74453, n74454, n74455, n74456, n74457, n74458, n74459, n74460, n74461, n74462, n74463, n74464, n74465, n74466, n74467, n74468, n74469, n74470, n74471, n74472, n74473, n74474, n74475, n74476, n74477, n74478, n74479, n74480, n74481, n74482, n74483, n74484, n74485, n74486, n74487, n74488, n74489, n74490, n74491, n74492, n74493, n74494, n74495, n74496, n74497, n74498, n74499, n74500, n74501, n74502, n74503, n74504, n74505, n74506, n74507, n74508, n74509, n74510, n74511, n74512, n74513, n74514, n74515, n74516, n74517, n74518, n74519, n74520, n74521, n74522, n74523, n74524, n74525, n74526, n74527, n74528, n74529, n74530, n74531, n74532, n74533, n74534, n74535, n74536, n74537, n74538, n74539, n74540, n74541, n74542, n74543, n74544, n74545, n74546, n74547, n74548, n74549, n74550, n74551, n74552, n74553, n74554, n74555, n74556, n74557, n74558, n74559, n74560, n74561, n74562, n74563, n74564, n74565, n74566, n74567, n74568, n74569, n74570, n74571, n74572, n74573, n74574, n74575, n74576, n74577, n74578, n74579, n74580, n74581, n74582, n74583, n74584, n74585, n74586, n74587, n74588, n74589, n74590, n74591, n74592, n74593, n74594, n74595, n74596, n74597, n74598, n74599, n74600, n74601, n74602, n74603, n74604, n74605, n74606, n74607, n74608, n74609, n74610, n74611, n74612, n74613, n74614, n74615, n74616, n74617, n74618, n74619, n74620, n74621, n74622, n74623, n74624, n74625, n74626, n74627, n74628, n74629, n74630, n74631, n74632, n74633, n74634, n74635, n74636, n74637, n74638, n74639, n74640, n74641, n74642, n74643, n74644, n74645, n74646, n74647, n74648, n74649, n74650, n74651, n74652, n74653, n74654, n74655, n74656, n74657, n74658, n74659, n74660, n74661, n74662, n74663, n74664, n74665, n74666, n74667, n74668, n74669, n74670, n74671, n74672, n74673, n74674, n74675, n74676, n74677, n74678, n74679, n74680, n74681, n74682, n74683, n74684, n74685, n74686, n74687, n74688, n74689, n74690, n74691, n74692, n74693, n74694, n74695, n74696, n74697, n74698, n74699, n74700, n74701, n74702, n74703, n74704, n74705, n74706, n74707, n74708, n74709, n74710, n74711, n74712, n74713, n74714, n74715, n74716, n74717, n74718, n74719, n74720, n74721, n74722, n74723, n74724, n74725, n74726, n74727, n74728, n74729, n74730, n74731, n74732, n74733, n74734, n74735, n74736, n74737, n74738, n74739, n74740;
  assign n17 = x0 & x8;
  assign n18 = x1 & x8;
  assign n19 = x0 & x9;
  assign n20 = n18 & n19;
  assign n21 = n18 | n19;
  assign n22 = ~n20 & n21;
  assign n23 = x2 & x8;
  assign n24 = x1 & x9;
  assign n25 = n23 & n24;
  assign n26 = n23 | n24;
  assign n27 = ~n25 & n26;
  assign n28 = n20 & n27;
  assign n29 = n20 | n27;
  assign n30 = ~n28 & n29;
  assign n31 = x0 & x10;
  assign n32 = n30 & n31;
  assign n33 = n30 | n31;
  assign n34 = ~n32 & n33;
  assign n441 = n20 | n25;
  assign n442 = (n25 & n27) | (n25 & n441) | (n27 & n441);
  assign n36 = x3 & x8;
  assign n37 = x2 & x9;
  assign n38 = n36 & n37;
  assign n39 = n36 | n37;
  assign n40 = ~n38 & n39;
  assign n41 = n442 & n40;
  assign n42 = n442 | n40;
  assign n43 = ~n41 & n42;
  assign n44 = x1 & x10;
  assign n45 = n43 & n44;
  assign n46 = n43 | n44;
  assign n47 = ~n45 & n46;
  assign n48 = n32 & n47;
  assign n49 = n32 | n47;
  assign n50 = ~n48 & n49;
  assign n51 = x0 & x11;
  assign n52 = n50 & n51;
  assign n53 = n50 | n51;
  assign n54 = ~n52 & n53;
  assign n443 = n32 | n45;
  assign n444 = (n45 & n47) | (n45 & n443) | (n47 & n443);
  assign n445 = n38 | n40;
  assign n446 = (n38 & n442) | (n38 & n445) | (n442 & n445);
  assign n57 = x4 & x8;
  assign n58 = x3 & x9;
  assign n59 = n57 & n58;
  assign n60 = n57 | n58;
  assign n61 = ~n59 & n60;
  assign n62 = n446 & n61;
  assign n63 = n446 | n61;
  assign n64 = ~n62 & n63;
  assign n65 = x2 & x10;
  assign n66 = n64 & n65;
  assign n67 = n64 | n65;
  assign n68 = ~n66 & n67;
  assign n69 = n444 & n68;
  assign n70 = n444 | n68;
  assign n71 = ~n69 & n70;
  assign n72 = x1 & x11;
  assign n73 = n71 & n72;
  assign n74 = n71 | n72;
  assign n75 = ~n73 & n74;
  assign n76 = n52 & n75;
  assign n77 = n52 | n75;
  assign n78 = ~n76 & n77;
  assign n79 = x0 & x12;
  assign n80 = n78 & n79;
  assign n81 = n78 | n79;
  assign n82 = ~n80 & n81;
  assign n447 = n52 | n73;
  assign n448 = (n73 & n75) | (n73 & n447) | (n75 & n447);
  assign n86 = x5 & x8;
  assign n87 = x4 & x9;
  assign n88 = n86 & n87;
  assign n89 = n86 | n87;
  assign n90 = ~n88 & n89;
  assign n449 = n59 | n61;
  assign n451 = n90 & n449;
  assign n452 = n59 & n90;
  assign n453 = (n446 & n451) | (n446 & n452) | (n451 & n452);
  assign n454 = n90 | n449;
  assign n455 = n59 | n90;
  assign n456 = (n446 & n454) | (n446 & n455) | (n454 & n455);
  assign n93 = ~n453 & n456;
  assign n94 = x3 & x10;
  assign n95 = n93 & n94;
  assign n96 = n93 | n94;
  assign n97 = ~n95 & n96;
  assign n457 = n66 & n97;
  assign n458 = (n69 & n97) | (n69 & n457) | (n97 & n457);
  assign n459 = n66 | n97;
  assign n460 = n69 | n459;
  assign n100 = ~n458 & n460;
  assign n101 = x2 & x11;
  assign n102 = n100 & n101;
  assign n103 = n100 | n101;
  assign n104 = ~n102 & n103;
  assign n105 = n448 & n104;
  assign n106 = n448 | n104;
  assign n107 = ~n105 & n106;
  assign n108 = x1 & x12;
  assign n109 = n107 & n108;
  assign n110 = n107 | n108;
  assign n111 = ~n109 & n110;
  assign n112 = n80 & n111;
  assign n113 = n80 | n111;
  assign n114 = ~n112 & n113;
  assign n115 = x0 & x13;
  assign n116 = n114 & n115;
  assign n117 = n114 | n115;
  assign n118 = ~n116 & n117;
  assign n461 = n80 | n109;
  assign n462 = (n109 & n111) | (n109 & n461) | (n111 & n461);
  assign n120 = n102 | n105;
  assign n123 = x6 & x8;
  assign n124 = x5 & x9;
  assign n125 = n123 & n124;
  assign n126 = n123 | n124;
  assign n127 = ~n125 & n126;
  assign n463 = n88 & n127;
  assign n464 = (n127 & n453) | (n127 & n463) | (n453 & n463);
  assign n465 = n88 | n127;
  assign n466 = n453 | n465;
  assign n130 = ~n464 & n466;
  assign n131 = x4 & x10;
  assign n132 = n130 & n131;
  assign n133 = n130 | n131;
  assign n134 = ~n132 & n133;
  assign n467 = n95 & n134;
  assign n468 = (n134 & n458) | (n134 & n467) | (n458 & n467);
  assign n469 = n95 | n134;
  assign n470 = n458 | n469;
  assign n137 = ~n468 & n470;
  assign n138 = x3 & x11;
  assign n139 = n137 & n138;
  assign n140 = n137 | n138;
  assign n141 = ~n139 & n140;
  assign n142 = n120 & n141;
  assign n143 = n120 | n141;
  assign n144 = ~n142 & n143;
  assign n145 = x2 & x12;
  assign n146 = n144 & n145;
  assign n147 = n144 | n145;
  assign n148 = ~n146 & n147;
  assign n149 = n462 & n148;
  assign n150 = n462 | n148;
  assign n151 = ~n149 & n150;
  assign n152 = x1 & x13;
  assign n153 = n151 & n152;
  assign n154 = n151 | n152;
  assign n155 = ~n153 & n154;
  assign n156 = n116 & n155;
  assign n157 = n116 | n155;
  assign n158 = ~n156 & n157;
  assign n159 = x0 & x14;
  assign n160 = n158 & n159;
  assign n161 = n158 | n159;
  assign n162 = ~n160 & n161;
  assign n2628 = n115 | n152;
  assign n2629 = (n114 & n152) | (n114 & n2628) | (n152 & n2628);
  assign n598 = (n116 & n151) | (n116 & n2629) | (n151 & n2629);
  assign n472 = (n153 & n155) | (n153 & n598) | (n155 & n598);
  assign n473 = n146 | n462;
  assign n474 = (n146 & n148) | (n146 & n473) | (n148 & n473);
  assign n475 = n139 | n141;
  assign n476 = (n120 & n139) | (n120 & n475) | (n139 & n475);
  assign n168 = x7 & x8;
  assign n169 = x6 & x9;
  assign n170 = n168 & n169;
  assign n171 = n168 | n169;
  assign n172 = ~n170 & n171;
  assign n599 = n88 | n125;
  assign n600 = (n125 & n127) | (n125 & n599) | (n127 & n599);
  assign n480 = n172 & n600;
  assign n478 = n125 | n127;
  assign n481 = n172 & n478;
  assign n482 = (n453 & n480) | (n453 & n481) | (n480 & n481);
  assign n483 = n172 | n600;
  assign n484 = n172 | n478;
  assign n485 = (n453 & n483) | (n453 & n484) | (n483 & n484);
  assign n175 = ~n482 & n485;
  assign n176 = x5 & x10;
  assign n177 = n175 & n176;
  assign n178 = n175 | n176;
  assign n179 = ~n177 & n178;
  assign n486 = n132 & n179;
  assign n487 = (n179 & n468) | (n179 & n486) | (n468 & n486);
  assign n488 = n132 | n179;
  assign n489 = n468 | n488;
  assign n182 = ~n487 & n489;
  assign n183 = x4 & x11;
  assign n184 = n182 & n183;
  assign n185 = n182 | n183;
  assign n186 = ~n184 & n185;
  assign n187 = n476 & n186;
  assign n188 = n476 | n186;
  assign n189 = ~n187 & n188;
  assign n190 = x3 & x12;
  assign n191 = n189 & n190;
  assign n192 = n189 | n190;
  assign n193 = ~n191 & n192;
  assign n194 = n474 & n193;
  assign n195 = n474 | n193;
  assign n196 = ~n194 & n195;
  assign n197 = x2 & x13;
  assign n198 = n196 & n197;
  assign n199 = n196 | n197;
  assign n200 = ~n198 & n199;
  assign n201 = n472 & n200;
  assign n202 = n472 | n200;
  assign n203 = ~n201 & n202;
  assign n204 = x1 & x14;
  assign n205 = n203 & n204;
  assign n206 = n203 | n204;
  assign n207 = ~n205 & n206;
  assign n208 = n160 & n207;
  assign n209 = n160 | n207;
  assign n210 = ~n208 & n209;
  assign n211 = x0 & x15;
  assign n212 = n210 & n211;
  assign n213 = n210 | n211;
  assign n214 = ~n212 & n213;
  assign n490 = n160 | n205;
  assign n491 = (n205 & n207) | (n205 & n490) | (n207 & n490);
  assign n216 = n198 | n201;
  assign n217 = n191 | n194;
  assign n492 = n184 | n186;
  assign n493 = (n184 & n476) | (n184 & n492) | (n476 & n492);
  assign n221 = x7 & x9;
  assign n497 = n170 & n221;
  assign n2630 = (n172 & n221) | (n172 & n497) | (n221 & n497);
  assign n2632 = (n478 & n2630) | (n478 & n497) | (n2630 & n497);
  assign n2633 = (n600 & n2630) | (n600 & n497) | (n2630 & n497);
  assign n605 = (n453 & n2632) | (n453 & n2633) | (n2632 & n2633);
  assign n499 = n170 | n221;
  assign n2634 = n172 | n499;
  assign n2635 = (n478 & n499) | (n478 & n2634) | (n499 & n2634);
  assign n2636 = (n499 & n600) | (n499 & n2634) | (n600 & n2634);
  assign n608 = (n453 & n2635) | (n453 & n2636) | (n2635 & n2636);
  assign n224 = ~n605 & n608;
  assign n225 = x6 & x10;
  assign n226 = n224 & n225;
  assign n227 = n224 | n225;
  assign n228 = ~n226 & n227;
  assign n495 = n177 | n179;
  assign n609 = n228 & n495;
  assign n601 = n132 | n177;
  assign n602 = (n177 & n179) | (n177 & n601) | (n179 & n601);
  assign n610 = n228 & n602;
  assign n611 = (n468 & n609) | (n468 & n610) | (n609 & n610);
  assign n612 = n228 | n495;
  assign n613 = n228 | n602;
  assign n614 = (n468 & n612) | (n468 & n613) | (n612 & n613);
  assign n231 = ~n611 & n614;
  assign n232 = x5 & x11;
  assign n233 = n231 & n232;
  assign n234 = n231 | n232;
  assign n235 = ~n233 & n234;
  assign n236 = n493 & n235;
  assign n237 = n493 | n235;
  assign n238 = ~n236 & n237;
  assign n239 = x4 & x12;
  assign n240 = n238 & n239;
  assign n241 = n238 | n239;
  assign n242 = ~n240 & n241;
  assign n243 = n217 & n242;
  assign n244 = n217 | n242;
  assign n245 = ~n243 & n244;
  assign n246 = x3 & x13;
  assign n247 = n245 & n246;
  assign n248 = n245 | n246;
  assign n249 = ~n247 & n248;
  assign n250 = n216 & n249;
  assign n251 = n216 | n249;
  assign n252 = ~n250 & n251;
  assign n253 = x2 & x14;
  assign n254 = n252 & n253;
  assign n255 = n252 | n253;
  assign n256 = ~n254 & n255;
  assign n257 = n491 & n256;
  assign n258 = n491 | n256;
  assign n259 = ~n257 & n258;
  assign n260 = x1 & x15;
  assign n261 = n259 & n260;
  assign n262 = n259 | n260;
  assign n263 = ~n261 & n262;
  assign n264 = n212 & n263;
  assign n265 = n212 | n263;
  assign n266 = ~n264 & n265;
  assign n2637 = n211 | n260;
  assign n2638 = (n210 & n260) | (n210 & n2637) | (n260 & n2637);
  assign n616 = (n212 & n259) | (n212 & n2638) | (n259 & n2638);
  assign n502 = (n261 & n263) | (n261 & n616) | (n263 & n616);
  assign n503 = n254 | n491;
  assign n504 = (n254 & n256) | (n254 & n503) | (n256 & n503);
  assign n269 = n247 | n250;
  assign n505 = n240 | n242;
  assign n506 = (n217 & n240) | (n217 & n505) | (n240 & n505);
  assign n273 = x7 & x10;
  assign n512 = n221 & n273;
  assign n617 = n170 & n512;
  assign n2639 = (n172 & n512) | (n172 & n617) | (n512 & n617);
  assign n2640 = n512 & n617;
  assign n2641 = (n478 & n2639) | (n478 & n2640) | (n2639 & n2640);
  assign n2642 = (n600 & n2639) | (n600 & n2640) | (n2639 & n2640);
  assign n620 = (n453 & n2641) | (n453 & n2642) | (n2641 & n2642);
  assign n515 = n221 | n273;
  assign n621 = (n170 & n273) | (n170 & n515) | (n273 & n515);
  assign n2643 = (n172 & n515) | (n172 & n621) | (n515 & n621);
  assign n2644 = n515 & n621;
  assign n2645 = (n478 & n2643) | (n478 & n2644) | (n2643 & n2644);
  assign n2646 = (n600 & n2643) | (n600 & n2644) | (n2643 & n2644);
  assign n624 = (n453 & n2645) | (n453 & n2646) | (n2645 & n2646);
  assign n276 = ~n620 & n624;
  assign n518 = n226 & n276;
  assign n625 = (n228 & n276) | (n228 & n518) | (n276 & n518);
  assign n626 = (n495 & n518) | (n495 & n625) | (n518 & n625);
  assign n627 = (n518 & n602) | (n518 & n625) | (n602 & n625);
  assign n628 = (n468 & n626) | (n468 & n627) | (n626 & n627);
  assign n521 = n226 | n276;
  assign n629 = n228 | n521;
  assign n630 = (n495 & n521) | (n495 & n629) | (n521 & n629);
  assign n631 = (n521 & n602) | (n521 & n629) | (n602 & n629);
  assign n632 = (n468 & n630) | (n468 & n631) | (n630 & n631);
  assign n279 = ~n628 & n632;
  assign n280 = x6 & x11;
  assign n281 = n279 & n280;
  assign n282 = n279 | n280;
  assign n283 = ~n281 & n282;
  assign n507 = n233 | n235;
  assign n633 = n283 & n507;
  assign n634 = n233 & n283;
  assign n635 = (n493 & n633) | (n493 & n634) | (n633 & n634);
  assign n636 = n283 | n507;
  assign n637 = n233 | n283;
  assign n638 = (n493 & n636) | (n493 & n637) | (n636 & n637);
  assign n286 = ~n635 & n638;
  assign n287 = x5 & x12;
  assign n288 = n286 & n287;
  assign n289 = n286 | n287;
  assign n290 = ~n288 & n289;
  assign n291 = n506 & n290;
  assign n292 = n506 | n290;
  assign n293 = ~n291 & n292;
  assign n294 = x4 & x13;
  assign n295 = n293 & n294;
  assign n296 = n293 | n294;
  assign n297 = ~n295 & n296;
  assign n298 = n269 & n297;
  assign n299 = n269 | n297;
  assign n300 = ~n298 & n299;
  assign n301 = x3 & x14;
  assign n302 = n300 & n301;
  assign n303 = n300 | n301;
  assign n304 = ~n302 & n303;
  assign n305 = n504 & n304;
  assign n306 = n504 | n304;
  assign n307 = ~n305 & n306;
  assign n308 = x2 & x15;
  assign n309 = n307 & n308;
  assign n310 = n307 | n308;
  assign n311 = ~n309 & n310;
  assign n312 = n502 & n311;
  assign n313 = n502 | n311;
  assign n314 = ~n312 & n313;
  assign n523 = n309 | n502;
  assign n524 = (n309 & n311) | (n309 & n523) | (n311 & n523);
  assign n525 = n302 | n504;
  assign n526 = (n302 & n304) | (n302 & n525) | (n304 & n525);
  assign n527 = n295 | n297;
  assign n528 = (n269 & n295) | (n269 & n527) | (n295 & n527);
  assign n321 = x7 & x11;
  assign n2647 = n321 & n2642;
  assign n2648 = n321 & n2641;
  assign n2649 = (n453 & n2647) | (n453 & n2648) | (n2647 & n2648);
  assign n534 = (n321 & n628) | (n321 & n2649) | (n628 & n2649);
  assign n2650 = n321 | n2642;
  assign n2651 = n321 | n2641;
  assign n2652 = (n453 & n2650) | (n453 & n2651) | (n2650 & n2651);
  assign n536 = n628 | n2652;
  assign n324 = ~n534 & n536;
  assign n538 = n281 & n324;
  assign n639 = (n283 & n324) | (n283 & n538) | (n324 & n538);
  assign n640 = (n507 & n538) | (n507 & n639) | (n538 & n639);
  assign n641 = (n233 & n538) | (n233 & n639) | (n538 & n639);
  assign n642 = (n493 & n640) | (n493 & n641) | (n640 & n641);
  assign n541 = n281 | n324;
  assign n643 = n283 | n541;
  assign n644 = (n507 & n541) | (n507 & n643) | (n541 & n643);
  assign n645 = (n233 & n541) | (n233 & n643) | (n541 & n643);
  assign n646 = (n493 & n644) | (n493 & n645) | (n644 & n645);
  assign n327 = ~n642 & n646;
  assign n328 = x6 & x12;
  assign n329 = n327 & n328;
  assign n330 = n327 | n328;
  assign n331 = ~n329 & n330;
  assign n529 = n288 | n290;
  assign n647 = n331 & n529;
  assign n648 = n288 & n331;
  assign n649 = (n506 & n647) | (n506 & n648) | (n647 & n648);
  assign n650 = n331 | n529;
  assign n651 = n288 | n331;
  assign n652 = (n506 & n650) | (n506 & n651) | (n650 & n651);
  assign n334 = ~n649 & n652;
  assign n335 = x5 & x13;
  assign n336 = n334 & n335;
  assign n337 = n334 | n335;
  assign n338 = ~n336 & n337;
  assign n339 = n528 & n338;
  assign n340 = n528 | n338;
  assign n341 = ~n339 & n340;
  assign n342 = x4 & x14;
  assign n343 = n341 & n342;
  assign n344 = n341 | n342;
  assign n345 = ~n343 & n344;
  assign n346 = n526 & n345;
  assign n347 = n526 | n345;
  assign n348 = ~n346 & n347;
  assign n349 = x3 & x15;
  assign n350 = n348 & n349;
  assign n351 = n348 | n349;
  assign n352 = ~n350 & n351;
  assign n353 = n524 & n352;
  assign n354 = n524 | n352;
  assign n355 = ~n353 & n354;
  assign n356 = n350 | n353;
  assign n361 = x7 & x12;
  assign n653 = n361 & n2649;
  assign n654 = n321 & n361;
  assign n655 = (n628 & n653) | (n628 & n654) | (n653 & n654);
  assign n548 = (n361 & n642) | (n361 & n655) | (n642 & n655);
  assign n656 = n361 | n2649;
  assign n657 = n321 | n361;
  assign n658 = (n628 & n656) | (n628 & n657) | (n656 & n657);
  assign n550 = n642 | n658;
  assign n364 = ~n548 & n550;
  assign n552 = n329 & n364;
  assign n659 = (n331 & n364) | (n331 & n552) | (n364 & n552);
  assign n660 = (n529 & n552) | (n529 & n659) | (n552 & n659);
  assign n661 = (n288 & n552) | (n288 & n659) | (n552 & n659);
  assign n662 = (n506 & n660) | (n506 & n661) | (n660 & n661);
  assign n555 = n329 | n364;
  assign n663 = n331 | n555;
  assign n664 = (n529 & n555) | (n529 & n663) | (n555 & n663);
  assign n665 = (n288 & n555) | (n288 & n663) | (n555 & n663);
  assign n666 = (n506 & n664) | (n506 & n665) | (n664 & n665);
  assign n367 = ~n662 & n666;
  assign n368 = x6 & x13;
  assign n369 = n367 & n368;
  assign n370 = n367 | n368;
  assign n371 = ~n369 & n370;
  assign n543 = n336 | n338;
  assign n667 = n371 & n543;
  assign n668 = n336 & n371;
  assign n669 = (n528 & n667) | (n528 & n668) | (n667 & n668);
  assign n670 = n371 | n543;
  assign n671 = n336 | n371;
  assign n672 = (n528 & n670) | (n528 & n671) | (n670 & n671);
  assign n374 = ~n669 & n672;
  assign n375 = x5 & x14;
  assign n376 = n374 & n375;
  assign n377 = n374 | n375;
  assign n378 = ~n376 & n377;
  assign n673 = n343 & n378;
  assign n674 = (n346 & n378) | (n346 & n673) | (n378 & n673);
  assign n675 = n343 | n378;
  assign n676 = n346 | n675;
  assign n381 = ~n674 & n676;
  assign n382 = x4 & x15;
  assign n383 = n381 & n382;
  assign n384 = n381 | n382;
  assign n385 = ~n383 & n384;
  assign n386 = n356 & n385;
  assign n387 = n356 | n385;
  assign n388 = ~n386 & n387;
  assign n677 = n383 | n385;
  assign n678 = (n356 & n383) | (n356 & n677) | (n383 & n677);
  assign n357 = n343 | n346;
  assign n393 = x7 & x13;
  assign n680 = n361 & n393;
  assign n3415 = n680 & n2649;
  assign n2654 = n393 & n654;
  assign n2655 = (n628 & n3415) | (n628 & n2654) | (n3415 & n2654);
  assign n681 = (n642 & n2655) | (n642 & n680) | (n2655 & n680);
  assign n562 = (n393 & n662) | (n393 & n681) | (n662 & n681);
  assign n683 = n361 | n393;
  assign n3416 = (n393 & n683) | (n393 & n2649) | (n683 & n2649);
  assign n2657 = n393 | n654;
  assign n2658 = (n628 & n3416) | (n628 & n2657) | (n3416 & n2657);
  assign n684 = (n642 & n2658) | (n642 & n683) | (n2658 & n683);
  assign n564 = n662 | n684;
  assign n396 = ~n562 & n564;
  assign n566 = n369 & n396;
  assign n685 = (n371 & n396) | (n371 & n566) | (n396 & n566);
  assign n686 = (n543 & n566) | (n543 & n685) | (n566 & n685);
  assign n687 = (n336 & n566) | (n336 & n685) | (n566 & n685);
  assign n688 = (n528 & n686) | (n528 & n687) | (n686 & n687);
  assign n569 = n369 | n396;
  assign n689 = n371 | n569;
  assign n690 = (n543 & n569) | (n543 & n689) | (n569 & n689);
  assign n691 = (n336 & n569) | (n336 & n689) | (n569 & n689);
  assign n692 = (n528 & n690) | (n528 & n691) | (n690 & n691);
  assign n399 = ~n688 & n692;
  assign n400 = x6 & x14;
  assign n401 = n399 & n400;
  assign n402 = n399 | n400;
  assign n403 = ~n401 & n402;
  assign n557 = n376 | n378;
  assign n693 = n403 & n557;
  assign n694 = n376 & n403;
  assign n695 = (n357 & n693) | (n357 & n694) | (n693 & n694);
  assign n696 = n403 | n557;
  assign n697 = n376 | n403;
  assign n698 = (n357 & n696) | (n357 & n697) | (n696 & n697);
  assign n406 = ~n695 & n698;
  assign n407 = x5 & x15;
  assign n408 = n406 & n407;
  assign n409 = n406 | n407;
  assign n410 = ~n408 & n409;
  assign n411 = n678 & n410;
  assign n412 = n678 | n410;
  assign n413 = ~n411 & n412;
  assign n571 = n408 | n410;
  assign n572 = (n678 & n408) | (n678 & n571) | (n408 & n571);
  assign n417 = x7 & x14;
  assign n2660 = n417 & n680;
  assign n11787 = n2649 & n2660;
  assign n700 = n393 & n417;
  assign n11788 = n654 & n700;
  assign n3419 = (n628 & n11787) | (n628 & n11788) | (n11787 & n11788);
  assign n2661 = (n642 & n3419) | (n642 & n2660) | (n3419 & n2660);
  assign n701 = (n662 & n2661) | (n662 & n700) | (n2661 & n700);
  assign n576 = (n417 & n688) | (n417 & n701) | (n688 & n701);
  assign n2663 = n417 | n680;
  assign n11789 = (n417 & n2649) | (n417 & n2663) | (n2649 & n2663);
  assign n703 = n393 | n417;
  assign n11790 = (n417 & n654) | (n417 & n703) | (n654 & n703);
  assign n3422 = (n628 & n11789) | (n628 & n11790) | (n11789 & n11790);
  assign n2664 = (n642 & n3422) | (n642 & n2663) | (n3422 & n2663);
  assign n704 = (n662 & n2664) | (n662 & n703) | (n2664 & n703);
  assign n578 = n688 | n704;
  assign n420 = ~n576 & n578;
  assign n580 = n401 & n420;
  assign n705 = (n403 & n420) | (n403 & n580) | (n420 & n580);
  assign n706 = (n557 & n580) | (n557 & n705) | (n580 & n705);
  assign n707 = (n376 & n580) | (n376 & n705) | (n580 & n705);
  assign n708 = (n357 & n706) | (n357 & n707) | (n706 & n707);
  assign n583 = n401 | n420;
  assign n709 = n403 | n583;
  assign n710 = (n557 & n583) | (n557 & n709) | (n583 & n709);
  assign n711 = (n376 & n583) | (n376 & n709) | (n583 & n709);
  assign n712 = (n357 & n710) | (n357 & n711) | (n710 & n711);
  assign n423 = ~n708 & n712;
  assign n424 = x6 & x15;
  assign n425 = n423 & n424;
  assign n426 = n423 | n424;
  assign n427 = ~n425 & n426;
  assign n428 = n572 & n427;
  assign n429 = n572 | n427;
  assign n430 = ~n428 & n429;
  assign n433 = x7 & x15;
  assign n714 = n417 & n433;
  assign n11794 = n680 & n714;
  assign n15521 = n2649 & n11794;
  assign n11792 = n433 & n11788;
  assign n11793 = (n628 & n15521) | (n628 & n11792) | (n15521 & n11792);
  assign n3425 = (n642 & n11793) | (n642 & n11794) | (n11793 & n11794);
  assign n2666 = n433 & n700;
  assign n2667 = (n662 & n3425) | (n662 & n2666) | (n3425 & n2666);
  assign n715 = (n688 & n2667) | (n688 & n714) | (n2667 & n714);
  assign n588 = (n433 & n708) | (n433 & n715) | (n708 & n715);
  assign n717 = n417 | n433;
  assign n11798 = (n433 & n680) | (n433 & n717) | (n680 & n717);
  assign n15522 = (n433 & n2649) | (n433 & n11798) | (n2649 & n11798);
  assign n11796 = n433 | n11788;
  assign n11797 = (n628 & n15522) | (n628 & n11796) | (n15522 & n11796);
  assign n3428 = (n642 & n11797) | (n642 & n11798) | (n11797 & n11798);
  assign n2669 = n433 | n700;
  assign n2670 = (n662 & n3428) | (n662 & n2669) | (n3428 & n2669);
  assign n718 = (n688 & n2670) | (n688 & n717) | (n2670 & n717);
  assign n590 = n708 | n718;
  assign n436 = ~n588 & n590;
  assign n592 = n425 & n436;
  assign n719 = (n427 & n436) | (n427 & n592) | (n436 & n592);
  assign n593 = (n572 & n719) | (n572 & n592) | (n719 & n592);
  assign n595 = n425 | n436;
  assign n720 = n427 | n595;
  assign n596 = (n572 & n720) | (n572 & n595) | (n720 & n595);
  assign n439 = ~n593 & n596;
  assign n721 = n588 | n719;
  assign n722 = n588 | n592;
  assign n723 = (n572 & n721) | (n572 & n722) | (n721 & n722);
  assign n756 = x16 & x32;
  assign n757 = x17 & x32;
  assign n758 = x16 & x33;
  assign n759 = n757 & n758;
  assign n760 = n757 | n758;
  assign n761 = ~n759 & n760;
  assign n762 = x18 & x32;
  assign n763 = x17 & x33;
  assign n764 = n762 & n763;
  assign n765 = n762 | n763;
  assign n766 = ~n764 & n765;
  assign n767 = n759 & n766;
  assign n768 = n759 | n766;
  assign n769 = ~n767 & n768;
  assign n770 = x16 & x34;
  assign n771 = n769 & n770;
  assign n772 = n769 | n770;
  assign n773 = ~n771 & n772;
  assign n2671 = n759 | n764;
  assign n2672 = (n764 & n766) | (n764 & n2671) | (n766 & n2671);
  assign n775 = x19 & x32;
  assign n776 = x18 & x33;
  assign n777 = n775 & n776;
  assign n778 = n775 | n776;
  assign n779 = ~n777 & n778;
  assign n780 = n2672 & n779;
  assign n781 = n2672 | n779;
  assign n782 = ~n780 & n781;
  assign n783 = x17 & x34;
  assign n784 = n782 & n783;
  assign n785 = n782 | n783;
  assign n786 = ~n784 & n785;
  assign n787 = n771 & n786;
  assign n788 = n771 | n786;
  assign n789 = ~n787 & n788;
  assign n790 = x16 & x35;
  assign n791 = n789 & n790;
  assign n792 = n789 | n790;
  assign n793 = ~n791 & n792;
  assign n2673 = n771 | n784;
  assign n2674 = (n784 & n786) | (n784 & n2673) | (n786 & n2673);
  assign n2675 = n777 | n779;
  assign n2676 = (n777 & n2672) | (n777 & n2675) | (n2672 & n2675);
  assign n796 = x20 & x32;
  assign n797 = x19 & x33;
  assign n798 = n796 & n797;
  assign n799 = n796 | n797;
  assign n800 = ~n798 & n799;
  assign n801 = n2676 & n800;
  assign n802 = n2676 | n800;
  assign n803 = ~n801 & n802;
  assign n804 = x18 & x34;
  assign n805 = n803 & n804;
  assign n806 = n803 | n804;
  assign n807 = ~n805 & n806;
  assign n808 = n2674 & n807;
  assign n809 = n2674 | n807;
  assign n810 = ~n808 & n809;
  assign n811 = x17 & x35;
  assign n812 = n810 & n811;
  assign n813 = n810 | n811;
  assign n814 = ~n812 & n813;
  assign n815 = n791 & n814;
  assign n816 = n791 | n814;
  assign n817 = ~n815 & n816;
  assign n818 = x16 & x36;
  assign n819 = n817 & n818;
  assign n820 = n817 | n818;
  assign n821 = ~n819 & n820;
  assign n2677 = n791 | n812;
  assign n2678 = (n812 & n814) | (n812 & n2677) | (n814 & n2677);
  assign n825 = x21 & x32;
  assign n826 = x20 & x33;
  assign n827 = n825 & n826;
  assign n828 = n825 | n826;
  assign n829 = ~n827 & n828;
  assign n2679 = n798 | n800;
  assign n2681 = n829 & n2679;
  assign n2682 = n798 & n829;
  assign n2683 = (n2676 & n2681) | (n2676 & n2682) | (n2681 & n2682);
  assign n2684 = n829 | n2679;
  assign n2685 = n798 | n829;
  assign n2686 = (n2676 & n2684) | (n2676 & n2685) | (n2684 & n2685);
  assign n832 = ~n2683 & n2686;
  assign n833 = x19 & x34;
  assign n834 = n832 & n833;
  assign n835 = n832 | n833;
  assign n836 = ~n834 & n835;
  assign n2687 = n805 & n836;
  assign n2688 = (n808 & n836) | (n808 & n2687) | (n836 & n2687);
  assign n2689 = n805 | n836;
  assign n2690 = n808 | n2689;
  assign n839 = ~n2688 & n2690;
  assign n840 = x18 & x35;
  assign n841 = n839 & n840;
  assign n842 = n839 | n840;
  assign n843 = ~n841 & n842;
  assign n844 = n2678 & n843;
  assign n845 = n2678 | n843;
  assign n846 = ~n844 & n845;
  assign n847 = x17 & x36;
  assign n848 = n846 & n847;
  assign n849 = n846 | n847;
  assign n850 = ~n848 & n849;
  assign n851 = n819 & n850;
  assign n852 = n819 | n850;
  assign n853 = ~n851 & n852;
  assign n854 = x16 & x37;
  assign n855 = n853 & n854;
  assign n856 = n853 | n854;
  assign n857 = ~n855 & n856;
  assign n2691 = n819 | n848;
  assign n2692 = (n848 & n850) | (n848 & n2691) | (n850 & n2691);
  assign n859 = n841 | n844;
  assign n862 = x22 & x32;
  assign n863 = x21 & x33;
  assign n864 = n862 & n863;
  assign n865 = n862 | n863;
  assign n866 = ~n864 & n865;
  assign n2693 = n827 & n866;
  assign n2694 = (n866 & n2683) | (n866 & n2693) | (n2683 & n2693);
  assign n2695 = n827 | n866;
  assign n2696 = n2683 | n2695;
  assign n869 = ~n2694 & n2696;
  assign n870 = x20 & x34;
  assign n871 = n869 & n870;
  assign n872 = n869 | n870;
  assign n873 = ~n871 & n872;
  assign n2697 = n834 & n873;
  assign n2698 = (n873 & n2688) | (n873 & n2697) | (n2688 & n2697);
  assign n2699 = n834 | n873;
  assign n2700 = n2688 | n2699;
  assign n876 = ~n2698 & n2700;
  assign n877 = x19 & x35;
  assign n878 = n876 & n877;
  assign n879 = n876 | n877;
  assign n880 = ~n878 & n879;
  assign n881 = n859 & n880;
  assign n882 = n859 | n880;
  assign n883 = ~n881 & n882;
  assign n884 = x18 & x36;
  assign n885 = n883 & n884;
  assign n886 = n883 | n884;
  assign n887 = ~n885 & n886;
  assign n888 = n2692 & n887;
  assign n889 = n2692 | n887;
  assign n890 = ~n888 & n889;
  assign n891 = x17 & x37;
  assign n892 = n890 & n891;
  assign n893 = n890 | n891;
  assign n894 = ~n892 & n893;
  assign n895 = n855 & n894;
  assign n896 = n855 | n894;
  assign n897 = ~n895 & n896;
  assign n898 = x16 & x38;
  assign n899 = n897 & n898;
  assign n900 = n897 | n898;
  assign n901 = ~n899 & n900;
  assign n11799 = n854 | n891;
  assign n11800 = (n853 & n891) | (n853 & n11799) | (n891 & n11799);
  assign n3430 = (n855 & n890) | (n855 & n11800) | (n890 & n11800);
  assign n2702 = (n892 & n894) | (n892 & n3430) | (n894 & n3430);
  assign n2703 = n885 | n2692;
  assign n2704 = (n885 & n887) | (n885 & n2703) | (n887 & n2703);
  assign n2705 = n878 | n880;
  assign n2706 = (n859 & n878) | (n859 & n2705) | (n878 & n2705);
  assign n907 = x23 & x32;
  assign n908 = x22 & x33;
  assign n909 = n907 & n908;
  assign n910 = n907 | n908;
  assign n911 = ~n909 & n910;
  assign n3431 = n827 | n864;
  assign n3432 = (n864 & n866) | (n864 & n3431) | (n866 & n3431);
  assign n2710 = n911 & n3432;
  assign n2708 = n864 | n866;
  assign n2711 = n911 & n2708;
  assign n2712 = (n2683 & n2710) | (n2683 & n2711) | (n2710 & n2711);
  assign n2713 = n911 | n3432;
  assign n2714 = n911 | n2708;
  assign n2715 = (n2683 & n2713) | (n2683 & n2714) | (n2713 & n2714);
  assign n914 = ~n2712 & n2715;
  assign n915 = x21 & x34;
  assign n916 = n914 & n915;
  assign n917 = n914 | n915;
  assign n918 = ~n916 & n917;
  assign n2716 = n871 & n918;
  assign n2717 = (n918 & n2698) | (n918 & n2716) | (n2698 & n2716);
  assign n2718 = n871 | n918;
  assign n2719 = n2698 | n2718;
  assign n921 = ~n2717 & n2719;
  assign n922 = x20 & x35;
  assign n923 = n921 & n922;
  assign n924 = n921 | n922;
  assign n925 = ~n923 & n924;
  assign n926 = n2706 & n925;
  assign n927 = n2706 | n925;
  assign n928 = ~n926 & n927;
  assign n929 = x19 & x36;
  assign n930 = n928 & n929;
  assign n931 = n928 | n929;
  assign n932 = ~n930 & n931;
  assign n933 = n2704 & n932;
  assign n934 = n2704 | n932;
  assign n935 = ~n933 & n934;
  assign n936 = x18 & x37;
  assign n937 = n935 & n936;
  assign n938 = n935 | n936;
  assign n939 = ~n937 & n938;
  assign n940 = n2702 & n939;
  assign n941 = n2702 | n939;
  assign n942 = ~n940 & n941;
  assign n943 = x17 & x38;
  assign n944 = n942 & n943;
  assign n945 = n942 | n943;
  assign n946 = ~n944 & n945;
  assign n947 = n899 & n946;
  assign n948 = n899 | n946;
  assign n949 = ~n947 & n948;
  assign n950 = x16 & x39;
  assign n951 = n949 & n950;
  assign n952 = n949 | n950;
  assign n953 = ~n951 & n952;
  assign n2720 = n899 | n944;
  assign n2721 = (n944 & n946) | (n944 & n2720) | (n946 & n2720);
  assign n955 = n937 | n940;
  assign n956 = n930 | n933;
  assign n2722 = n923 | n925;
  assign n2723 = (n923 & n2706) | (n923 & n2722) | (n2706 & n2722);
  assign n960 = x24 & x32;
  assign n961 = x23 & x33;
  assign n962 = n960 & n961;
  assign n963 = n960 | n961;
  assign n964 = ~n962 & n963;
  assign n2727 = n909 & n964;
  assign n3435 = (n964 & n2711) | (n964 & n2727) | (n2711 & n2727);
  assign n3436 = (n964 & n2710) | (n964 & n2727) | (n2710 & n2727);
  assign n3437 = (n2683 & n3435) | (n2683 & n3436) | (n3435 & n3436);
  assign n2729 = n909 | n964;
  assign n3438 = n2711 | n2729;
  assign n3439 = n2710 | n2729;
  assign n3440 = (n2683 & n3438) | (n2683 & n3439) | (n3438 & n3439);
  assign n967 = ~n3437 & n3440;
  assign n968 = x22 & x34;
  assign n969 = n967 & n968;
  assign n970 = n967 | n968;
  assign n971 = ~n969 & n970;
  assign n2725 = n916 | n918;
  assign n3441 = n971 & n2725;
  assign n3433 = n871 | n916;
  assign n3434 = (n916 & n918) | (n916 & n3433) | (n918 & n3433);
  assign n3442 = n971 & n3434;
  assign n3443 = (n2698 & n3441) | (n2698 & n3442) | (n3441 & n3442);
  assign n3444 = n971 | n2725;
  assign n3445 = n971 | n3434;
  assign n3446 = (n2698 & n3444) | (n2698 & n3445) | (n3444 & n3445);
  assign n974 = ~n3443 & n3446;
  assign n975 = x21 & x35;
  assign n976 = n974 & n975;
  assign n977 = n974 | n975;
  assign n978 = ~n976 & n977;
  assign n979 = n2723 & n978;
  assign n980 = n2723 | n978;
  assign n981 = ~n979 & n980;
  assign n982 = x20 & x36;
  assign n983 = n981 & n982;
  assign n984 = n981 | n982;
  assign n985 = ~n983 & n984;
  assign n986 = n956 & n985;
  assign n987 = n956 | n985;
  assign n988 = ~n986 & n987;
  assign n989 = x19 & x37;
  assign n990 = n988 & n989;
  assign n991 = n988 | n989;
  assign n992 = ~n990 & n991;
  assign n993 = n955 & n992;
  assign n994 = n955 | n992;
  assign n995 = ~n993 & n994;
  assign n996 = x18 & x38;
  assign n997 = n995 & n996;
  assign n998 = n995 | n996;
  assign n999 = ~n997 & n998;
  assign n1000 = n2721 & n999;
  assign n1001 = n2721 | n999;
  assign n1002 = ~n1000 & n1001;
  assign n1003 = x17 & x39;
  assign n1004 = n1002 & n1003;
  assign n1005 = n1002 | n1003;
  assign n1006 = ~n1004 & n1005;
  assign n1007 = n951 & n1006;
  assign n1008 = n951 | n1006;
  assign n1009 = ~n1007 & n1008;
  assign n1010 = x16 & x40;
  assign n1011 = n1009 & n1010;
  assign n1012 = n1009 | n1010;
  assign n1013 = ~n1011 & n1012;
  assign n11801 = n950 | n1003;
  assign n11802 = (n949 & n1003) | (n949 & n11801) | (n1003 & n11801);
  assign n3448 = (n951 & n1002) | (n951 & n11802) | (n1002 & n11802);
  assign n2732 = (n1004 & n1006) | (n1004 & n3448) | (n1006 & n3448);
  assign n2733 = n997 | n2721;
  assign n2734 = (n997 & n999) | (n997 & n2733) | (n999 & n2733);
  assign n1016 = n990 | n993;
  assign n2735 = n983 | n985;
  assign n2736 = (n956 & n983) | (n956 & n2735) | (n983 & n2735);
  assign n2726 = (n2698 & n3434) | (n2698 & n2725) | (n3434 & n2725);
  assign n1021 = x25 & x32;
  assign n1022 = x24 & x33;
  assign n1023 = n1021 & n1022;
  assign n1024 = n1021 | n1022;
  assign n1025 = ~n1023 & n1024;
  assign n3449 = n909 | n962;
  assign n3450 = (n962 & n964) | (n962 & n3449) | (n964 & n3449);
  assign n2744 = n1025 & n3450;
  assign n2742 = n962 | n964;
  assign n2745 = n1025 & n2742;
  assign n3451 = (n2711 & n2744) | (n2711 & n2745) | (n2744 & n2745);
  assign n3452 = (n2710 & n2744) | (n2710 & n2745) | (n2744 & n2745);
  assign n3453 = (n2683 & n3451) | (n2683 & n3452) | (n3451 & n3452);
  assign n2747 = n1025 | n3450;
  assign n2748 = n1025 | n2742;
  assign n3454 = (n2711 & n2747) | (n2711 & n2748) | (n2747 & n2748);
  assign n3455 = (n2710 & n2747) | (n2710 & n2748) | (n2747 & n2748);
  assign n3456 = (n2683 & n3454) | (n2683 & n3455) | (n3454 & n3455);
  assign n1028 = ~n3453 & n3456;
  assign n1029 = x23 & x34;
  assign n1030 = n1028 & n1029;
  assign n1031 = n1028 | n1029;
  assign n1032 = ~n1030 & n1031;
  assign n2739 = n969 | n971;
  assign n2750 = n1032 & n2739;
  assign n2751 = n969 & n1032;
  assign n2752 = (n2726 & n2750) | (n2726 & n2751) | (n2750 & n2751);
  assign n2753 = n1032 | n2739;
  assign n2754 = n969 | n1032;
  assign n2755 = (n2726 & n2753) | (n2726 & n2754) | (n2753 & n2754);
  assign n1035 = ~n2752 & n2755;
  assign n1036 = x22 & x35;
  assign n1037 = n1035 & n1036;
  assign n1038 = n1035 | n1036;
  assign n1039 = ~n1037 & n1038;
  assign n2737 = n976 | n978;
  assign n3457 = n1039 & n2737;
  assign n3458 = n976 & n1039;
  assign n3459 = (n2723 & n3457) | (n2723 & n3458) | (n3457 & n3458);
  assign n3460 = n1039 | n2737;
  assign n3461 = n976 | n1039;
  assign n3462 = (n2723 & n3460) | (n2723 & n3461) | (n3460 & n3461);
  assign n1042 = ~n3459 & n3462;
  assign n1043 = x21 & x36;
  assign n1044 = n1042 & n1043;
  assign n1045 = n1042 | n1043;
  assign n1046 = ~n1044 & n1045;
  assign n1047 = n2736 & n1046;
  assign n1048 = n2736 | n1046;
  assign n1049 = ~n1047 & n1048;
  assign n1050 = x20 & x37;
  assign n1051 = n1049 & n1050;
  assign n1052 = n1049 | n1050;
  assign n1053 = ~n1051 & n1052;
  assign n1054 = n1016 & n1053;
  assign n1055 = n1016 | n1053;
  assign n1056 = ~n1054 & n1055;
  assign n1057 = x19 & x38;
  assign n1058 = n1056 & n1057;
  assign n1059 = n1056 | n1057;
  assign n1060 = ~n1058 & n1059;
  assign n1061 = n2734 & n1060;
  assign n1062 = n2734 | n1060;
  assign n1063 = ~n1061 & n1062;
  assign n1064 = x18 & x39;
  assign n1065 = n1063 & n1064;
  assign n1066 = n1063 | n1064;
  assign n1067 = ~n1065 & n1066;
  assign n1068 = n2732 & n1067;
  assign n1069 = n2732 | n1067;
  assign n1070 = ~n1068 & n1069;
  assign n1071 = x17 & x40;
  assign n1072 = n1070 & n1071;
  assign n1073 = n1070 | n1071;
  assign n1074 = ~n1072 & n1073;
  assign n1075 = n1011 & n1074;
  assign n1076 = n1011 | n1074;
  assign n1077 = ~n1075 & n1076;
  assign n1078 = x16 & x41;
  assign n1079 = n1077 & n1078;
  assign n1080 = n1077 | n1078;
  assign n1081 = ~n1079 & n1080;
  assign n11803 = n1010 | n1071;
  assign n11804 = (n1009 & n1071) | (n1009 & n11803) | (n1071 & n11803);
  assign n3464 = (n1011 & n1070) | (n1011 & n11804) | (n1070 & n11804);
  assign n2757 = (n1072 & n1074) | (n1072 & n3464) | (n1074 & n3464);
  assign n2758 = n1065 | n2732;
  assign n2759 = (n1065 & n1067) | (n1065 & n2758) | (n1067 & n2758);
  assign n2760 = n1058 | n2734;
  assign n2761 = (n1058 & n1060) | (n1058 & n2760) | (n1060 & n2760);
  assign n2762 = n1051 | n1053;
  assign n2763 = (n1016 & n1051) | (n1016 & n2762) | (n1051 & n2762);
  assign n2738 = (n976 & n2723) | (n976 & n2737) | (n2723 & n2737);
  assign n3465 = n1023 | n1025;
  assign n3466 = (n1023 & n3450) | (n1023 & n3465) | (n3450 & n3465);
  assign n3467 = (n1023 & n2742) | (n1023 & n3465) | (n2742 & n3465);
  assign n3468 = (n2711 & n3466) | (n2711 & n3467) | (n3466 & n3467);
  assign n3469 = (n2710 & n3466) | (n2710 & n3467) | (n3466 & n3467);
  assign n3470 = (n2683 & n3468) | (n2683 & n3469) | (n3468 & n3469);
  assign n1090 = x26 & x32;
  assign n1091 = x25 & x33;
  assign n1092 = n1090 & n1091;
  assign n1093 = n1090 | n1091;
  assign n1094 = ~n1092 & n1093;
  assign n1095 = n3470 & n1094;
  assign n1096 = n3470 | n1094;
  assign n1097 = ~n1095 & n1096;
  assign n1098 = x24 & x34;
  assign n1099 = n1097 & n1098;
  assign n1100 = n1097 | n1098;
  assign n1101 = ~n1099 & n1100;
  assign n2771 = n1030 & n1101;
  assign n3471 = (n1101 & n2750) | (n1101 & n2771) | (n2750 & n2771);
  assign n3472 = (n1101 & n2751) | (n1101 & n2771) | (n2751 & n2771);
  assign n3473 = (n2726 & n3471) | (n2726 & n3472) | (n3471 & n3472);
  assign n2773 = n1030 | n1101;
  assign n3474 = n2750 | n2773;
  assign n3475 = n2751 | n2773;
  assign n3476 = (n2726 & n3474) | (n2726 & n3475) | (n3474 & n3475);
  assign n1104 = ~n3473 & n3476;
  assign n1105 = x23 & x35;
  assign n1106 = n1104 & n1105;
  assign n1107 = n1104 | n1105;
  assign n1108 = ~n1106 & n1107;
  assign n2766 = n1037 | n1039;
  assign n2775 = n1108 & n2766;
  assign n2776 = n1037 & n1108;
  assign n2777 = (n2738 & n2775) | (n2738 & n2776) | (n2775 & n2776);
  assign n2778 = n1108 | n2766;
  assign n2779 = n1037 | n1108;
  assign n2780 = (n2738 & n2778) | (n2738 & n2779) | (n2778 & n2779);
  assign n1111 = ~n2777 & n2780;
  assign n1112 = x22 & x36;
  assign n1113 = n1111 & n1112;
  assign n1114 = n1111 | n1112;
  assign n1115 = ~n1113 & n1114;
  assign n2764 = n1044 | n1046;
  assign n3477 = n1115 & n2764;
  assign n3478 = n1044 & n1115;
  assign n3479 = (n2736 & n3477) | (n2736 & n3478) | (n3477 & n3478);
  assign n3480 = n1115 | n2764;
  assign n3481 = n1044 | n1115;
  assign n3482 = (n2736 & n3480) | (n2736 & n3481) | (n3480 & n3481);
  assign n1118 = ~n3479 & n3482;
  assign n1119 = x21 & x37;
  assign n1120 = n1118 & n1119;
  assign n1121 = n1118 | n1119;
  assign n1122 = ~n1120 & n1121;
  assign n1123 = n2763 & n1122;
  assign n1124 = n2763 | n1122;
  assign n1125 = ~n1123 & n1124;
  assign n1126 = x20 & x38;
  assign n1127 = n1125 & n1126;
  assign n1128 = n1125 | n1126;
  assign n1129 = ~n1127 & n1128;
  assign n1130 = n2761 & n1129;
  assign n1131 = n2761 | n1129;
  assign n1132 = ~n1130 & n1131;
  assign n1133 = x19 & x39;
  assign n1134 = n1132 & n1133;
  assign n1135 = n1132 | n1133;
  assign n1136 = ~n1134 & n1135;
  assign n1137 = n2759 & n1136;
  assign n1138 = n2759 | n1136;
  assign n1139 = ~n1137 & n1138;
  assign n1140 = x18 & x40;
  assign n1141 = n1139 & n1140;
  assign n1142 = n1139 | n1140;
  assign n1143 = ~n1141 & n1142;
  assign n1144 = n2757 & n1143;
  assign n1145 = n2757 | n1143;
  assign n1146 = ~n1144 & n1145;
  assign n1147 = x17 & x41;
  assign n1148 = n1146 & n1147;
  assign n1149 = n1146 | n1147;
  assign n1150 = ~n1148 & n1149;
  assign n1151 = n1079 & n1150;
  assign n1152 = n1079 | n1150;
  assign n1153 = ~n1151 & n1152;
  assign n1154 = x16 & x42;
  assign n1155 = n1153 & n1154;
  assign n1156 = n1153 | n1154;
  assign n1157 = ~n1155 & n1156;
  assign n2781 = n1079 | n1148;
  assign n2782 = (n1148 & n1150) | (n1148 & n2781) | (n1150 & n2781);
  assign n1159 = n1141 | n1144;
  assign n1160 = n1134 | n1137;
  assign n2765 = (n1044 & n2736) | (n1044 & n2764) | (n2736 & n2764);
  assign n2788 = n1099 | n1101;
  assign n3483 = n1030 | n1099;
  assign n3484 = (n1099 & n1101) | (n1099 & n3483) | (n1101 & n3483);
  assign n3485 = (n2750 & n2788) | (n2750 & n3484) | (n2788 & n3484);
  assign n3486 = (n2751 & n2788) | (n2751 & n3484) | (n2788 & n3484);
  assign n3487 = (n2726 & n3485) | (n2726 & n3486) | (n3485 & n3486);
  assign n1167 = x27 & x32;
  assign n1168 = x26 & x33;
  assign n1169 = n1167 & n1168;
  assign n1170 = n1167 | n1168;
  assign n1171 = ~n1169 & n1170;
  assign n2790 = n1092 | n1094;
  assign n2792 = n1171 & n2790;
  assign n2793 = n1092 & n1171;
  assign n2794 = (n3470 & n2792) | (n3470 & n2793) | (n2792 & n2793);
  assign n2795 = n1171 | n2790;
  assign n2796 = n1092 | n1171;
  assign n2797 = (n3470 & n2795) | (n3470 & n2796) | (n2795 & n2796);
  assign n1174 = ~n2794 & n2797;
  assign n1175 = x25 & x34;
  assign n1176 = n1174 & n1175;
  assign n1177 = n1174 | n1175;
  assign n1178 = ~n1176 & n1177;
  assign n1179 = n3487 & n1178;
  assign n1180 = n3487 | n1178;
  assign n1181 = ~n1179 & n1180;
  assign n1182 = x24 & x35;
  assign n1183 = n1181 & n1182;
  assign n1184 = n1181 | n1182;
  assign n1185 = ~n1183 & n1184;
  assign n2798 = n1106 & n1185;
  assign n2799 = (n1185 & n2777) | (n1185 & n2798) | (n2777 & n2798);
  assign n2800 = n1106 | n1185;
  assign n2801 = n2777 | n2800;
  assign n1188 = ~n2799 & n2801;
  assign n1189 = x23 & x36;
  assign n1190 = n1188 & n1189;
  assign n1191 = n1188 | n1189;
  assign n1192 = ~n1190 & n1191;
  assign n2785 = n1113 | n1115;
  assign n2802 = n1192 & n2785;
  assign n2803 = n1113 & n1192;
  assign n2804 = (n2765 & n2802) | (n2765 & n2803) | (n2802 & n2803);
  assign n2805 = n1192 | n2785;
  assign n2806 = n1113 | n1192;
  assign n2807 = (n2765 & n2805) | (n2765 & n2806) | (n2805 & n2806);
  assign n1195 = ~n2804 & n2807;
  assign n1196 = x22 & x37;
  assign n1197 = n1195 & n1196;
  assign n1198 = n1195 | n1196;
  assign n1199 = ~n1197 & n1198;
  assign n2783 = n1120 | n1122;
  assign n3488 = n1199 & n2783;
  assign n3489 = n1120 & n1199;
  assign n3490 = (n2763 & n3488) | (n2763 & n3489) | (n3488 & n3489);
  assign n3491 = n1199 | n2783;
  assign n3492 = n1120 | n1199;
  assign n3493 = (n2763 & n3491) | (n2763 & n3492) | (n3491 & n3492);
  assign n1202 = ~n3490 & n3493;
  assign n1203 = x21 & x38;
  assign n1204 = n1202 & n1203;
  assign n1205 = n1202 | n1203;
  assign n1206 = ~n1204 & n1205;
  assign n3494 = n1127 & n1206;
  assign n3495 = (n1130 & n1206) | (n1130 & n3494) | (n1206 & n3494);
  assign n3496 = n1127 | n1206;
  assign n3497 = n1130 | n3496;
  assign n1209 = ~n3495 & n3497;
  assign n1210 = x20 & x39;
  assign n1211 = n1209 & n1210;
  assign n1212 = n1209 | n1210;
  assign n1213 = ~n1211 & n1212;
  assign n1214 = n1160 & n1213;
  assign n1215 = n1160 | n1213;
  assign n1216 = ~n1214 & n1215;
  assign n1217 = x19 & x40;
  assign n1218 = n1216 & n1217;
  assign n1219 = n1216 | n1217;
  assign n1220 = ~n1218 & n1219;
  assign n1221 = n1159 & n1220;
  assign n1222 = n1159 | n1220;
  assign n1223 = ~n1221 & n1222;
  assign n1224 = x18 & x41;
  assign n1225 = n1223 & n1224;
  assign n1226 = n1223 | n1224;
  assign n1227 = ~n1225 & n1226;
  assign n1228 = n2782 & n1227;
  assign n1229 = n2782 | n1227;
  assign n1230 = ~n1228 & n1229;
  assign n1231 = x17 & x42;
  assign n1232 = n1230 & n1231;
  assign n1233 = n1230 | n1231;
  assign n1234 = ~n1232 & n1233;
  assign n1235 = n1155 & n1234;
  assign n1236 = n1155 | n1234;
  assign n1237 = ~n1235 & n1236;
  assign n1238 = x16 & x43;
  assign n1239 = n1237 & n1238;
  assign n1240 = n1237 | n1238;
  assign n1241 = ~n1239 & n1240;
  assign n11805 = n1154 | n1231;
  assign n11806 = (n1153 & n1231) | (n1153 & n11805) | (n1231 & n11805);
  assign n3499 = (n1155 & n1230) | (n1155 & n11806) | (n1230 & n11806);
  assign n2809 = (n1232 & n1234) | (n1232 & n3499) | (n1234 & n3499);
  assign n2810 = n1225 | n2782;
  assign n2811 = (n1225 & n1227) | (n1225 & n2810) | (n1227 & n2810);
  assign n1244 = n1218 | n1221;
  assign n3500 = n1211 | n1213;
  assign n3501 = (n1160 & n1211) | (n1160 & n3500) | (n1211 & n3500);
  assign n1161 = n1127 | n1130;
  assign n2784 = (n1120 & n2763) | (n1120 & n2783) | (n2763 & n2783);
  assign n1252 = x28 & x32;
  assign n1253 = x27 & x33;
  assign n1254 = n1252 & n1253;
  assign n1255 = n1252 | n1253;
  assign n1256 = ~n1254 & n1255;
  assign n3502 = n1169 | n1171;
  assign n3503 = (n1169 & n2790) | (n1169 & n3502) | (n2790 & n3502);
  assign n2821 = n1256 & n3503;
  assign n3504 = n1092 | n1169;
  assign n3505 = (n1169 & n1171) | (n1169 & n3504) | (n1171 & n3504);
  assign n2822 = n1256 & n3505;
  assign n2823 = (n3470 & n2821) | (n3470 & n2822) | (n2821 & n2822);
  assign n2824 = n1256 | n3503;
  assign n2825 = n1256 | n3505;
  assign n2826 = (n3470 & n2824) | (n3470 & n2825) | (n2824 & n2825);
  assign n1259 = ~n2823 & n2826;
  assign n1260 = x26 & x34;
  assign n1261 = n1259 & n1260;
  assign n1262 = n1259 | n1260;
  assign n1263 = ~n1261 & n1262;
  assign n2816 = n1176 | n1178;
  assign n2827 = n1263 & n2816;
  assign n2828 = n1176 & n1263;
  assign n2829 = (n3487 & n2827) | (n3487 & n2828) | (n2827 & n2828);
  assign n2830 = n1263 | n2816;
  assign n2831 = n1176 | n1263;
  assign n2832 = (n3487 & n2830) | (n3487 & n2831) | (n2830 & n2831);
  assign n1266 = ~n2829 & n2832;
  assign n1267 = x25 & x35;
  assign n1268 = n1266 & n1267;
  assign n1269 = n1266 | n1267;
  assign n1270 = ~n1268 & n1269;
  assign n2833 = n1183 & n1270;
  assign n3506 = (n1270 & n2798) | (n1270 & n2833) | (n2798 & n2833);
  assign n3507 = (n1185 & n1270) | (n1185 & n2833) | (n1270 & n2833);
  assign n3508 = (n2777 & n3506) | (n2777 & n3507) | (n3506 & n3507);
  assign n2835 = n1183 | n1270;
  assign n3509 = n2798 | n2835;
  assign n3510 = n1185 | n2835;
  assign n3511 = (n2777 & n3509) | (n2777 & n3510) | (n3509 & n3510);
  assign n1273 = ~n3508 & n3511;
  assign n1274 = x24 & x36;
  assign n1275 = n1273 & n1274;
  assign n1276 = n1273 | n1274;
  assign n1277 = ~n1275 & n1276;
  assign n2837 = n1190 & n1277;
  assign n2838 = (n1277 & n2804) | (n1277 & n2837) | (n2804 & n2837);
  assign n2839 = n1190 | n1277;
  assign n2840 = n2804 | n2839;
  assign n1280 = ~n2838 & n2840;
  assign n1281 = x23 & x37;
  assign n1282 = n1280 & n1281;
  assign n1283 = n1280 | n1281;
  assign n1284 = ~n1282 & n1283;
  assign n2814 = n1197 | n1199;
  assign n2841 = n1284 & n2814;
  assign n2842 = n1197 & n1284;
  assign n2843 = (n2784 & n2841) | (n2784 & n2842) | (n2841 & n2842);
  assign n2844 = n1284 | n2814;
  assign n2845 = n1197 | n1284;
  assign n2846 = (n2784 & n2844) | (n2784 & n2845) | (n2844 & n2845);
  assign n1287 = ~n2843 & n2846;
  assign n1288 = x22 & x38;
  assign n1289 = n1287 & n1288;
  assign n1290 = n1287 | n1288;
  assign n1291 = ~n1289 & n1290;
  assign n2812 = n1204 | n1206;
  assign n3512 = n1291 & n2812;
  assign n3513 = n1204 & n1291;
  assign n3514 = (n1161 & n3512) | (n1161 & n3513) | (n3512 & n3513);
  assign n3515 = n1291 | n2812;
  assign n3516 = n1204 | n1291;
  assign n3517 = (n1161 & n3515) | (n1161 & n3516) | (n3515 & n3516);
  assign n1294 = ~n3514 & n3517;
  assign n1295 = x21 & x39;
  assign n1296 = n1294 & n1295;
  assign n1297 = n1294 | n1295;
  assign n1298 = ~n1296 & n1297;
  assign n1299 = n3501 & n1298;
  assign n1300 = n3501 | n1298;
  assign n1301 = ~n1299 & n1300;
  assign n1302 = x20 & x40;
  assign n1303 = n1301 & n1302;
  assign n1304 = n1301 | n1302;
  assign n1305 = ~n1303 & n1304;
  assign n1306 = n1244 & n1305;
  assign n1307 = n1244 | n1305;
  assign n1308 = ~n1306 & n1307;
  assign n1309 = x19 & x41;
  assign n1310 = n1308 & n1309;
  assign n1311 = n1308 | n1309;
  assign n1312 = ~n1310 & n1311;
  assign n1313 = n2811 & n1312;
  assign n1314 = n2811 | n1312;
  assign n1315 = ~n1313 & n1314;
  assign n1316 = x18 & x42;
  assign n1317 = n1315 & n1316;
  assign n1318 = n1315 | n1316;
  assign n1319 = ~n1317 & n1318;
  assign n1320 = n2809 & n1319;
  assign n1321 = n2809 | n1319;
  assign n1322 = ~n1320 & n1321;
  assign n1323 = x17 & x43;
  assign n1324 = n1322 & n1323;
  assign n1325 = n1322 | n1323;
  assign n1326 = ~n1324 & n1325;
  assign n1327 = n1239 & n1326;
  assign n1328 = n1239 | n1326;
  assign n1329 = ~n1327 & n1328;
  assign n1330 = x16 & x44;
  assign n1331 = n1329 & n1330;
  assign n1332 = n1329 | n1330;
  assign n1333 = ~n1331 & n1332;
  assign n11807 = n1238 | n1323;
  assign n11808 = (n1237 & n1323) | (n1237 & n11807) | (n1323 & n11807);
  assign n3519 = (n1239 & n1322) | (n1239 & n11808) | (n1322 & n11808);
  assign n2848 = (n1324 & n1326) | (n1324 & n3519) | (n1326 & n3519);
  assign n2849 = n1317 | n2809;
  assign n2850 = (n1317 & n1319) | (n1317 & n2849) | (n1319 & n2849);
  assign n2851 = n1310 | n2811;
  assign n2852 = (n1310 & n1312) | (n1310 & n2851) | (n1312 & n2851);
  assign n3520 = n1303 | n1305;
  assign n3521 = (n1244 & n1303) | (n1244 & n3520) | (n1303 & n3520);
  assign n2853 = n1296 | n1298;
  assign n2854 = (n3501 & n1296) | (n3501 & n2853) | (n1296 & n2853);
  assign n2813 = (n1161 & n1204) | (n1161 & n2812) | (n1204 & n2812);
  assign n2858 = n1268 | n1270;
  assign n3522 = n1183 | n1268;
  assign n3523 = (n1268 & n1270) | (n1268 & n3522) | (n1270 & n3522);
  assign n3524 = (n2798 & n2858) | (n2798 & n3523) | (n2858 & n3523);
  assign n3525 = (n1185 & n2858) | (n1185 & n3523) | (n2858 & n3523);
  assign n3526 = (n2777 & n3524) | (n2777 & n3525) | (n3524 & n3525);
  assign n1345 = x29 & x32;
  assign n1346 = x28 & x33;
  assign n1347 = n1345 & n1346;
  assign n1348 = n1345 | n1346;
  assign n1349 = ~n1347 & n1348;
  assign n3531 = n1254 | n1256;
  assign n11809 = n1349 & n3531;
  assign n11810 = n1254 & n1349;
  assign n11811 = (n3503 & n11809) | (n3503 & n11810) | (n11809 & n11810);
  assign n3533 = (n1254 & n3505) | (n1254 & n3531) | (n3505 & n3531);
  assign n3535 = n1349 & n3533;
  assign n3536 = (n3470 & n11811) | (n3470 & n3535) | (n11811 & n3535);
  assign n11812 = n1349 | n3531;
  assign n11813 = n1254 | n1349;
  assign n11814 = (n3503 & n11812) | (n3503 & n11813) | (n11812 & n11813);
  assign n3538 = n1349 | n3533;
  assign n3539 = (n3470 & n11814) | (n3470 & n3538) | (n11814 & n3538);
  assign n1352 = ~n3536 & n3539;
  assign n1353 = x27 & x34;
  assign n1354 = n1352 & n1353;
  assign n1355 = n1352 | n1353;
  assign n1356 = ~n1354 & n1355;
  assign n3527 = n1261 | n1263;
  assign n3528 = (n1261 & n2816) | (n1261 & n3527) | (n2816 & n3527);
  assign n3540 = n1356 & n3528;
  assign n3529 = n1176 | n1261;
  assign n3530 = (n1261 & n1263) | (n1261 & n3529) | (n1263 & n3529);
  assign n3541 = n1356 & n3530;
  assign n3542 = (n3487 & n3540) | (n3487 & n3541) | (n3540 & n3541);
  assign n3543 = n1356 | n3528;
  assign n3544 = n1356 | n3530;
  assign n3545 = (n3487 & n3543) | (n3487 & n3544) | (n3543 & n3544);
  assign n1359 = ~n3542 & n3545;
  assign n1360 = x26 & x35;
  assign n1361 = n1359 & n1360;
  assign n1362 = n1359 | n1360;
  assign n1363 = ~n1361 & n1362;
  assign n1364 = n3526 & n1363;
  assign n1365 = n3526 | n1363;
  assign n1366 = ~n1364 & n1365;
  assign n1367 = x25 & x36;
  assign n1368 = n1366 & n1367;
  assign n1369 = n1366 | n1367;
  assign n1370 = ~n1368 & n1369;
  assign n2866 = n1275 & n1370;
  assign n2867 = (n1370 & n2838) | (n1370 & n2866) | (n2838 & n2866);
  assign n2868 = n1275 | n1370;
  assign n2869 = n2838 | n2868;
  assign n1373 = ~n2867 & n2869;
  assign n1374 = x24 & x37;
  assign n1375 = n1373 & n1374;
  assign n1376 = n1373 | n1374;
  assign n1377 = ~n1375 & n1376;
  assign n2870 = n1282 & n1377;
  assign n2871 = (n1377 & n2843) | (n1377 & n2870) | (n2843 & n2870);
  assign n2872 = n1282 | n1377;
  assign n2873 = n2843 | n2872;
  assign n1380 = ~n2871 & n2873;
  assign n1381 = x23 & x38;
  assign n1382 = n1380 & n1381;
  assign n1383 = n1380 | n1381;
  assign n1384 = ~n1382 & n1383;
  assign n2855 = n1289 | n1291;
  assign n2874 = n1384 & n2855;
  assign n2875 = n1289 & n1384;
  assign n2876 = (n2813 & n2874) | (n2813 & n2875) | (n2874 & n2875);
  assign n2877 = n1384 | n2855;
  assign n2878 = n1289 | n1384;
  assign n2879 = (n2813 & n2877) | (n2813 & n2878) | (n2877 & n2878);
  assign n1387 = ~n2876 & n2879;
  assign n1388 = x22 & x39;
  assign n1389 = n1387 & n1388;
  assign n1390 = n1387 | n1388;
  assign n1391 = ~n1389 & n1390;
  assign n1392 = n2854 & n1391;
  assign n1393 = n2854 | n1391;
  assign n1394 = ~n1392 & n1393;
  assign n1395 = x21 & x40;
  assign n1396 = n1394 & n1395;
  assign n1397 = n1394 | n1395;
  assign n1398 = ~n1396 & n1397;
  assign n1399 = n3521 & n1398;
  assign n1400 = n3521 | n1398;
  assign n1401 = ~n1399 & n1400;
  assign n1402 = x20 & x41;
  assign n1403 = n1401 & n1402;
  assign n1404 = n1401 | n1402;
  assign n1405 = ~n1403 & n1404;
  assign n1406 = n2852 & n1405;
  assign n1407 = n2852 | n1405;
  assign n1408 = ~n1406 & n1407;
  assign n1409 = x19 & x42;
  assign n1410 = n1408 & n1409;
  assign n1411 = n1408 | n1409;
  assign n1412 = ~n1410 & n1411;
  assign n1413 = n2850 & n1412;
  assign n1414 = n2850 | n1412;
  assign n1415 = ~n1413 & n1414;
  assign n1416 = x18 & x43;
  assign n1417 = n1415 & n1416;
  assign n1418 = n1415 | n1416;
  assign n1419 = ~n1417 & n1418;
  assign n1420 = n2848 & n1419;
  assign n1421 = n2848 | n1419;
  assign n1422 = ~n1420 & n1421;
  assign n1423 = x17 & x44;
  assign n1424 = n1422 & n1423;
  assign n1425 = n1422 | n1423;
  assign n1426 = ~n1424 & n1425;
  assign n1427 = n1331 & n1426;
  assign n1428 = n1331 | n1426;
  assign n1429 = ~n1427 & n1428;
  assign n1430 = x16 & x45;
  assign n1431 = n1429 & n1430;
  assign n1432 = n1429 | n1430;
  assign n1433 = ~n1431 & n1432;
  assign n2880 = n1331 | n1424;
  assign n2881 = (n1424 & n1426) | (n1424 & n2880) | (n1426 & n2880);
  assign n2882 = n1417 | n2848;
  assign n2883 = (n1417 & n1419) | (n1417 & n2882) | (n1419 & n2882);
  assign n2884 = n1410 | n2850;
  assign n2885 = (n1410 & n1412) | (n1410 & n2884) | (n1412 & n2884);
  assign n2886 = n1403 | n2852;
  assign n2887 = (n1403 & n1405) | (n1403 & n2886) | (n1405 & n2886);
  assign n2888 = n1396 | n1398;
  assign n2889 = (n3521 & n1396) | (n3521 & n2888) | (n1396 & n2888);
  assign n1446 = x30 & x32;
  assign n1447 = x29 & x33;
  assign n1448 = n1446 & n1447;
  assign n1449 = n1446 | n1447;
  assign n1450 = ~n1448 & n1449;
  assign n2896 = n1347 | n1349;
  assign n2898 = n1450 & n2896;
  assign n2899 = n1347 & n1450;
  assign n3532 = (n1254 & n3503) | (n1254 & n3531) | (n3503 & n3531);
  assign n3546 = (n2898 & n2899) | (n2898 & n3532) | (n2899 & n3532);
  assign n3547 = (n2898 & n2899) | (n2898 & n3533) | (n2899 & n3533);
  assign n3548 = (n3470 & n3546) | (n3470 & n3547) | (n3546 & n3547);
  assign n2901 = n1450 | n2896;
  assign n2902 = n1347 | n1450;
  assign n3549 = (n2901 & n2902) | (n2901 & n3532) | (n2902 & n3532);
  assign n3550 = (n2901 & n2902) | (n2901 & n3533) | (n2902 & n3533);
  assign n3551 = (n3470 & n3549) | (n3470 & n3550) | (n3549 & n3550);
  assign n1453 = ~n3548 & n3551;
  assign n1454 = x28 & x34;
  assign n1455 = n1453 & n1454;
  assign n1456 = n1453 | n1454;
  assign n1457 = ~n1455 & n1456;
  assign n2894 = n1354 | n1356;
  assign n2904 = n1457 & n2894;
  assign n2905 = n1354 & n1457;
  assign n3552 = (n2904 & n2905) | (n2904 & n3528) | (n2905 & n3528);
  assign n3553 = (n2904 & n2905) | (n2904 & n3530) | (n2905 & n3530);
  assign n3554 = (n3487 & n3552) | (n3487 & n3553) | (n3552 & n3553);
  assign n2907 = n1457 | n2894;
  assign n2908 = n1354 | n1457;
  assign n3555 = (n2907 & n2908) | (n2907 & n3528) | (n2908 & n3528);
  assign n3556 = (n2907 & n2908) | (n2907 & n3530) | (n2908 & n3530);
  assign n3557 = (n3487 & n3555) | (n3487 & n3556) | (n3555 & n3556);
  assign n1460 = ~n3554 & n3557;
  assign n1461 = x27 & x35;
  assign n1462 = n1460 & n1461;
  assign n1463 = n1460 | n1461;
  assign n1464 = ~n1462 & n1463;
  assign n2892 = n1361 | n1363;
  assign n2910 = n1464 & n2892;
  assign n2911 = n1361 & n1464;
  assign n2912 = (n3526 & n2910) | (n3526 & n2911) | (n2910 & n2911);
  assign n2913 = n1464 | n2892;
  assign n2914 = n1361 | n1464;
  assign n2915 = (n3526 & n2913) | (n3526 & n2914) | (n2913 & n2914);
  assign n1467 = ~n2912 & n2915;
  assign n1468 = x26 & x36;
  assign n1469 = n1467 & n1468;
  assign n1470 = n1467 | n1468;
  assign n1471 = ~n1469 & n1470;
  assign n2916 = n1368 & n1471;
  assign n3558 = (n1471 & n2866) | (n1471 & n2916) | (n2866 & n2916);
  assign n3559 = (n1370 & n1471) | (n1370 & n2916) | (n1471 & n2916);
  assign n3560 = (n2838 & n3558) | (n2838 & n3559) | (n3558 & n3559);
  assign n2918 = n1368 | n1471;
  assign n3561 = n2866 | n2918;
  assign n3562 = n1370 | n2918;
  assign n3563 = (n2838 & n3561) | (n2838 & n3562) | (n3561 & n3562);
  assign n1474 = ~n3560 & n3563;
  assign n1475 = x25 & x37;
  assign n1476 = n1474 & n1475;
  assign n1477 = n1474 | n1475;
  assign n1478 = ~n1476 & n1477;
  assign n2920 = n1375 & n1478;
  assign n2921 = (n1478 & n2871) | (n1478 & n2920) | (n2871 & n2920);
  assign n2922 = n1375 | n1478;
  assign n2923 = n2871 | n2922;
  assign n1481 = ~n2921 & n2923;
  assign n1482 = x24 & x38;
  assign n1483 = n1481 & n1482;
  assign n1484 = n1481 | n1482;
  assign n1485 = ~n1483 & n1484;
  assign n2924 = n1382 & n1485;
  assign n2925 = (n1485 & n2876) | (n1485 & n2924) | (n2876 & n2924);
  assign n2926 = n1382 | n1485;
  assign n2927 = n2876 | n2926;
  assign n1488 = ~n2925 & n2927;
  assign n1489 = x23 & x39;
  assign n1490 = n1488 & n1489;
  assign n1491 = n1488 | n1489;
  assign n1492 = ~n1490 & n1491;
  assign n2890 = n1389 | n1391;
  assign n2928 = n1492 & n2890;
  assign n2929 = n1389 & n1492;
  assign n2930 = (n2854 & n2928) | (n2854 & n2929) | (n2928 & n2929);
  assign n2931 = n1492 | n2890;
  assign n2932 = n1389 | n1492;
  assign n2933 = (n2854 & n2931) | (n2854 & n2932) | (n2931 & n2932);
  assign n1495 = ~n2930 & n2933;
  assign n1496 = x22 & x40;
  assign n1497 = n1495 & n1496;
  assign n1498 = n1495 | n1496;
  assign n1499 = ~n1497 & n1498;
  assign n1500 = n2889 & n1499;
  assign n1501 = n2889 | n1499;
  assign n1502 = ~n1500 & n1501;
  assign n1503 = x21 & x41;
  assign n1504 = n1502 & n1503;
  assign n1505 = n1502 | n1503;
  assign n1506 = ~n1504 & n1505;
  assign n1507 = n2887 & n1506;
  assign n1508 = n2887 | n1506;
  assign n1509 = ~n1507 & n1508;
  assign n1510 = x20 & x42;
  assign n1511 = n1509 & n1510;
  assign n1512 = n1509 | n1510;
  assign n1513 = ~n1511 & n1512;
  assign n1514 = n2885 & n1513;
  assign n1515 = n2885 | n1513;
  assign n1516 = ~n1514 & n1515;
  assign n1517 = x19 & x43;
  assign n1518 = n1516 & n1517;
  assign n1519 = n1516 | n1517;
  assign n1520 = ~n1518 & n1519;
  assign n1521 = n2883 & n1520;
  assign n1522 = n2883 | n1520;
  assign n1523 = ~n1521 & n1522;
  assign n1524 = x18 & x44;
  assign n1525 = n1523 & n1524;
  assign n1526 = n1523 | n1524;
  assign n1527 = ~n1525 & n1526;
  assign n1528 = n2881 & n1527;
  assign n1529 = n2881 | n1527;
  assign n1530 = ~n1528 & n1529;
  assign n1531 = x17 & x45;
  assign n1532 = n1530 & n1531;
  assign n1533 = n1530 | n1531;
  assign n1534 = ~n1532 & n1533;
  assign n1535 = n1431 & n1534;
  assign n1536 = n1431 | n1534;
  assign n1537 = ~n1535 & n1536;
  assign n1538 = x16 & x46;
  assign n1539 = n1537 & n1538;
  assign n1540 = n1537 | n1538;
  assign n1541 = ~n1539 & n1540;
  assign n11815 = n1430 | n1531;
  assign n11816 = (n1429 & n1531) | (n1429 & n11815) | (n1531 & n11815);
  assign n3565 = (n1431 & n1530) | (n1431 & n11816) | (n1530 & n11816);
  assign n2935 = (n1532 & n1534) | (n1532 & n3565) | (n1534 & n3565);
  assign n3566 = n1525 | n2881;
  assign n3567 = (n1525 & n1527) | (n1525 & n3566) | (n1527 & n3566);
  assign n1544 = n1518 | n1521;
  assign n1545 = n1511 | n1514;
  assign n2939 = n1469 | n1471;
  assign n3568 = n1368 | n1469;
  assign n3569 = (n1469 & n1471) | (n1469 & n3568) | (n1471 & n3568);
  assign n3570 = (n2866 & n2939) | (n2866 & n3569) | (n2939 & n3569);
  assign n3571 = (n1370 & n2939) | (n1370 & n3569) | (n2939 & n3569);
  assign n3572 = (n2838 & n3570) | (n2838 & n3571) | (n3570 & n3571);
  assign n3573 = n1455 | n1457;
  assign n3574 = (n1455 & n2894) | (n1455 & n3573) | (n2894 & n3573);
  assign n3575 = n1354 | n1455;
  assign n3576 = (n1455 & n1457) | (n1455 & n3575) | (n1457 & n3575);
  assign n3577 = (n3528 & n3574) | (n3528 & n3576) | (n3574 & n3576);
  assign n3578 = (n3530 & n3574) | (n3530 & n3576) | (n3574 & n3576);
  assign n3579 = (n3487 & n3577) | (n3487 & n3578) | (n3577 & n3578);
  assign n1555 = x31 & x32;
  assign n1556 = x30 & x33;
  assign n1557 = n1555 & n1556;
  assign n1558 = n1555 | n1556;
  assign n1559 = ~n1557 & n1558;
  assign n3580 = n1448 | n1450;
  assign n3581 = (n1448 & n2896) | (n1448 & n3580) | (n2896 & n3580);
  assign n2947 = n1559 & n3581;
  assign n3582 = n1347 | n1448;
  assign n3583 = (n1448 & n1450) | (n1448 & n3582) | (n1450 & n3582);
  assign n2948 = n1559 & n3583;
  assign n3584 = (n2947 & n2948) | (n2947 & n3532) | (n2948 & n3532);
  assign n3585 = (n2947 & n2948) | (n2947 & n3533) | (n2948 & n3533);
  assign n3586 = (n3470 & n3584) | (n3470 & n3585) | (n3584 & n3585);
  assign n2950 = n1559 | n3581;
  assign n2951 = n1559 | n3583;
  assign n3587 = (n2950 & n2951) | (n2950 & n3532) | (n2951 & n3532);
  assign n3588 = (n2950 & n2951) | (n2950 & n3533) | (n2951 & n3533);
  assign n3589 = (n3470 & n3587) | (n3470 & n3588) | (n3587 & n3588);
  assign n1562 = ~n3586 & n3589;
  assign n1563 = x29 & x34;
  assign n1564 = n1562 & n1563;
  assign n1565 = n1562 | n1563;
  assign n1566 = ~n1564 & n1565;
  assign n1567 = n3579 & n1566;
  assign n1568 = n3579 | n1566;
  assign n1569 = ~n1567 & n1568;
  assign n1570 = x28 & x35;
  assign n1571 = n1569 & n1570;
  assign n1572 = n1569 | n1570;
  assign n1573 = ~n1571 & n1572;
  assign n2953 = n1462 & n1573;
  assign n3590 = (n1573 & n2910) | (n1573 & n2953) | (n2910 & n2953);
  assign n3591 = (n1573 & n2911) | (n1573 & n2953) | (n2911 & n2953);
  assign n3592 = (n3526 & n3590) | (n3526 & n3591) | (n3590 & n3591);
  assign n2955 = n1462 | n1573;
  assign n3593 = n2910 | n2955;
  assign n3594 = n2911 | n2955;
  assign n3595 = (n3526 & n3593) | (n3526 & n3594) | (n3593 & n3594);
  assign n1576 = ~n3592 & n3595;
  assign n1577 = x27 & x36;
  assign n1578 = n1576 & n1577;
  assign n1579 = n1576 | n1577;
  assign n1580 = ~n1578 & n1579;
  assign n1581 = n3572 & n1580;
  assign n1582 = n3572 | n1580;
  assign n1583 = ~n1581 & n1582;
  assign n1584 = x26 & x37;
  assign n1585 = n1583 & n1584;
  assign n1586 = n1583 | n1584;
  assign n1587 = ~n1585 & n1586;
  assign n2957 = n1476 & n1587;
  assign n2958 = (n1587 & n2921) | (n1587 & n2957) | (n2921 & n2957);
  assign n2959 = n1476 | n1587;
  assign n2960 = n2921 | n2959;
  assign n1590 = ~n2958 & n2960;
  assign n1591 = x25 & x38;
  assign n1592 = n1590 & n1591;
  assign n1593 = n1590 | n1591;
  assign n1594 = ~n1592 & n1593;
  assign n2961 = n1483 & n1594;
  assign n2962 = (n1594 & n2925) | (n1594 & n2961) | (n2925 & n2961);
  assign n2963 = n1483 | n1594;
  assign n2964 = n2925 | n2963;
  assign n1597 = ~n2962 & n2964;
  assign n1598 = x24 & x39;
  assign n1599 = n1597 & n1598;
  assign n1600 = n1597 | n1598;
  assign n1601 = ~n1599 & n1600;
  assign n2965 = n1490 & n1601;
  assign n2966 = (n1601 & n2930) | (n1601 & n2965) | (n2930 & n2965);
  assign n2967 = n1490 | n1601;
  assign n2968 = n2930 | n2967;
  assign n1604 = ~n2966 & n2968;
  assign n1605 = x23 & x40;
  assign n1606 = n1604 & n1605;
  assign n1607 = n1604 | n1605;
  assign n1608 = ~n1606 & n1607;
  assign n2936 = n1497 | n1499;
  assign n2969 = n1608 & n2936;
  assign n2970 = n1497 & n1608;
  assign n2971 = (n2889 & n2969) | (n2889 & n2970) | (n2969 & n2970);
  assign n2972 = n1608 | n2936;
  assign n2973 = n1497 | n1608;
  assign n2974 = (n2889 & n2972) | (n2889 & n2973) | (n2972 & n2973);
  assign n1611 = ~n2971 & n2974;
  assign n1612 = x22 & x41;
  assign n1613 = n1611 & n1612;
  assign n1614 = n1611 | n1612;
  assign n1615 = ~n1613 & n1614;
  assign n2975 = n1504 & n1615;
  assign n2976 = (n1507 & n1615) | (n1507 & n2975) | (n1615 & n2975);
  assign n2977 = n1504 | n1615;
  assign n2978 = n1507 | n2977;
  assign n1618 = ~n2976 & n2978;
  assign n1619 = x21 & x42;
  assign n1620 = n1618 & n1619;
  assign n1621 = n1618 | n1619;
  assign n1622 = ~n1620 & n1621;
  assign n1623 = n1545 & n1622;
  assign n1624 = n1545 | n1622;
  assign n1625 = ~n1623 & n1624;
  assign n1626 = x20 & x43;
  assign n1627 = n1625 & n1626;
  assign n1628 = n1625 | n1626;
  assign n1629 = ~n1627 & n1628;
  assign n1630 = n1544 & n1629;
  assign n1631 = n1544 | n1629;
  assign n1632 = ~n1630 & n1631;
  assign n1633 = x19 & x44;
  assign n1634 = n1632 & n1633;
  assign n1635 = n1632 | n1633;
  assign n1636 = ~n1634 & n1635;
  assign n1637 = n3567 & n1636;
  assign n1638 = n3567 | n1636;
  assign n1639 = ~n1637 & n1638;
  assign n1640 = x18 & x45;
  assign n1641 = n1639 & n1640;
  assign n1642 = n1639 | n1640;
  assign n1643 = ~n1641 & n1642;
  assign n1644 = n2935 & n1643;
  assign n1645 = n2935 | n1643;
  assign n1646 = ~n1644 & n1645;
  assign n1647 = x17 & x46;
  assign n1648 = n1646 & n1647;
  assign n1649 = n1646 | n1647;
  assign n1650 = ~n1648 & n1649;
  assign n1651 = n1539 & n1650;
  assign n1652 = n1539 | n1650;
  assign n1653 = ~n1651 & n1652;
  assign n1654 = x16 & x47;
  assign n1655 = n1653 & n1654;
  assign n1656 = n1653 | n1654;
  assign n1657 = ~n1655 & n1656;
  assign n11817 = n1538 | n1647;
  assign n11818 = (n1537 & n1647) | (n1537 & n11817) | (n1647 & n11817);
  assign n3597 = (n1539 & n1646) | (n1539 & n11818) | (n1646 & n11818);
  assign n2980 = (n1648 & n1650) | (n1648 & n3597) | (n1650 & n3597);
  assign n2981 = n1641 | n2935;
  assign n2982 = (n1641 & n1643) | (n1641 & n2981) | (n1643 & n2981);
  assign n3598 = n1634 | n3567;
  assign n3599 = (n1634 & n1636) | (n1634 & n3598) | (n1636 & n3598);
  assign n1661 = n1627 | n1630;
  assign n2983 = n1620 | n1622;
  assign n2984 = (n1545 & n1620) | (n1545 & n2983) | (n1620 & n2983);
  assign n2988 = n1571 | n1573;
  assign n3600 = n1462 | n1571;
  assign n3601 = (n1571 & n1573) | (n1571 & n3600) | (n1573 & n3600);
  assign n3602 = (n2910 & n2988) | (n2910 & n3601) | (n2988 & n3601);
  assign n3603 = (n2911 & n2988) | (n2911 & n3601) | (n2988 & n3601);
  assign n3604 = (n3526 & n3602) | (n3526 & n3603) | (n3602 & n3603);
  assign n1672 = x31 & x33;
  assign n3605 = n1557 | n1559;
  assign n3610 = (n1557 & n3583) | (n1557 & n3605) | (n3583 & n3605);
  assign n2996 = n1672 & n3610;
  assign n3608 = n1557 & n1672;
  assign n11819 = (n1559 & n1672) | (n1559 & n3608) | (n1672 & n3608);
  assign n3609 = (n3581 & n11819) | (n3581 & n3608) | (n11819 & n3608);
  assign n3611 = (n2996 & n3532) | (n2996 & n3609) | (n3532 & n3609);
  assign n3612 = (n2996 & n3533) | (n2996 & n3609) | (n3533 & n3609);
  assign n3613 = (n3470 & n3611) | (n3470 & n3612) | (n3611 & n3612);
  assign n2999 = n1672 | n3610;
  assign n3615 = n1557 | n1672;
  assign n11820 = n1559 | n3615;
  assign n3616 = (n3581 & n11820) | (n3581 & n3615) | (n11820 & n3615);
  assign n3617 = (n2999 & n3532) | (n2999 & n3616) | (n3532 & n3616);
  assign n3618 = (n2999 & n3533) | (n2999 & n3616) | (n3533 & n3616);
  assign n3619 = (n3470 & n3617) | (n3470 & n3618) | (n3617 & n3618);
  assign n1675 = ~n3613 & n3619;
  assign n1676 = x30 & x34;
  assign n1677 = n1675 & n1676;
  assign n1678 = n1675 | n1676;
  assign n1679 = ~n1677 & n1678;
  assign n2990 = n1564 | n1566;
  assign n3001 = n1679 & n2990;
  assign n3002 = n1564 & n1679;
  assign n3003 = (n3579 & n3001) | (n3579 & n3002) | (n3001 & n3002);
  assign n3004 = n1679 | n2990;
  assign n3005 = n1564 | n1679;
  assign n3006 = (n3579 & n3004) | (n3579 & n3005) | (n3004 & n3005);
  assign n1682 = ~n3003 & n3006;
  assign n1683 = x29 & x35;
  assign n1684 = n1682 & n1683;
  assign n1685 = n1682 | n1683;
  assign n1686 = ~n1684 & n1685;
  assign n1687 = n3604 & n1686;
  assign n1688 = n3604 | n1686;
  assign n1689 = ~n1687 & n1688;
  assign n1690 = x28 & x36;
  assign n1691 = n1689 & n1690;
  assign n1692 = n1689 | n1690;
  assign n1693 = ~n1691 & n1692;
  assign n2985 = n1578 | n1580;
  assign n3007 = n1693 & n2985;
  assign n3008 = n1578 & n1693;
  assign n3009 = (n3572 & n3007) | (n3572 & n3008) | (n3007 & n3008);
  assign n3010 = n1693 | n2985;
  assign n3011 = n1578 | n1693;
  assign n3012 = (n3572 & n3010) | (n3572 & n3011) | (n3010 & n3011);
  assign n1696 = ~n3009 & n3012;
  assign n1697 = x27 & x37;
  assign n1698 = n1696 & n1697;
  assign n1699 = n1696 | n1697;
  assign n1700 = ~n1698 & n1699;
  assign n3013 = n1585 & n1700;
  assign n3620 = (n1700 & n2957) | (n1700 & n3013) | (n2957 & n3013);
  assign n3621 = (n1587 & n1700) | (n1587 & n3013) | (n1700 & n3013);
  assign n3622 = (n2921 & n3620) | (n2921 & n3621) | (n3620 & n3621);
  assign n3015 = n1585 | n1700;
  assign n3623 = n2957 | n3015;
  assign n3624 = n1587 | n3015;
  assign n3625 = (n2921 & n3623) | (n2921 & n3624) | (n3623 & n3624);
  assign n1703 = ~n3622 & n3625;
  assign n1704 = x26 & x38;
  assign n1705 = n1703 & n1704;
  assign n1706 = n1703 | n1704;
  assign n1707 = ~n1705 & n1706;
  assign n3017 = n1592 & n1707;
  assign n3018 = (n1707 & n2962) | (n1707 & n3017) | (n2962 & n3017);
  assign n3019 = n1592 | n1707;
  assign n3020 = n2962 | n3019;
  assign n1710 = ~n3018 & n3020;
  assign n1711 = x25 & x39;
  assign n1712 = n1710 & n1711;
  assign n1713 = n1710 | n1711;
  assign n1714 = ~n1712 & n1713;
  assign n3021 = n1599 & n1714;
  assign n3022 = (n1714 & n2966) | (n1714 & n3021) | (n2966 & n3021);
  assign n3023 = n1599 | n1714;
  assign n3024 = n2966 | n3023;
  assign n1717 = ~n3022 & n3024;
  assign n1718 = x24 & x40;
  assign n1719 = n1717 & n1718;
  assign n1720 = n1717 | n1718;
  assign n1721 = ~n1719 & n1720;
  assign n3025 = n1606 & n1721;
  assign n3026 = (n1721 & n2971) | (n1721 & n3025) | (n2971 & n3025);
  assign n3027 = n1606 | n1721;
  assign n3028 = n2971 | n3027;
  assign n1724 = ~n3026 & n3028;
  assign n1725 = x23 & x41;
  assign n1726 = n1724 & n1725;
  assign n1727 = n1724 | n1725;
  assign n1728 = ~n1726 & n1727;
  assign n3029 = n1613 & n1728;
  assign n3030 = (n1728 & n2976) | (n1728 & n3029) | (n2976 & n3029);
  assign n3031 = n1613 | n1728;
  assign n3032 = n2976 | n3031;
  assign n1731 = ~n3030 & n3032;
  assign n1732 = x22 & x42;
  assign n1733 = n1731 & n1732;
  assign n1734 = n1731 | n1732;
  assign n1735 = ~n1733 & n1734;
  assign n1736 = n2984 & n1735;
  assign n1737 = n2984 | n1735;
  assign n1738 = ~n1736 & n1737;
  assign n1739 = x21 & x43;
  assign n1740 = n1738 & n1739;
  assign n1741 = n1738 | n1739;
  assign n1742 = ~n1740 & n1741;
  assign n1743 = n1661 & n1742;
  assign n1744 = n1661 | n1742;
  assign n1745 = ~n1743 & n1744;
  assign n1746 = x20 & x44;
  assign n1747 = n1745 & n1746;
  assign n1748 = n1745 | n1746;
  assign n1749 = ~n1747 & n1748;
  assign n1750 = n3599 & n1749;
  assign n1751 = n3599 | n1749;
  assign n1752 = ~n1750 & n1751;
  assign n1753 = x19 & x45;
  assign n1754 = n1752 & n1753;
  assign n1755 = n1752 | n1753;
  assign n1756 = ~n1754 & n1755;
  assign n1757 = n2982 & n1756;
  assign n1758 = n2982 | n1756;
  assign n1759 = ~n1757 & n1758;
  assign n1760 = x18 & x46;
  assign n1761 = n1759 & n1760;
  assign n1762 = n1759 | n1760;
  assign n1763 = ~n1761 & n1762;
  assign n1764 = n2980 & n1763;
  assign n1765 = n2980 | n1763;
  assign n1766 = ~n1764 & n1765;
  assign n1767 = x17 & x47;
  assign n1768 = n1766 & n1767;
  assign n1769 = n1766 | n1767;
  assign n1770 = ~n1768 & n1769;
  assign n1771 = n1655 & n1770;
  assign n1772 = n1655 | n1770;
  assign n1773 = ~n1771 & n1772;
  assign n11821 = n1654 | n1767;
  assign n11822 = (n1653 & n1767) | (n1653 & n11821) | (n1767 & n11821);
  assign n3627 = (n1655 & n1766) | (n1655 & n11822) | (n1766 & n11822);
  assign n3034 = (n1768 & n1770) | (n1768 & n3627) | (n1770 & n3627);
  assign n3035 = n1761 | n2980;
  assign n3036 = (n1761 & n1763) | (n1761 & n3035) | (n1763 & n3035);
  assign n3037 = n1754 | n2982;
  assign n3038 = (n1754 & n1756) | (n1754 & n3037) | (n1756 & n3037);
  assign n3628 = n1747 | n3599;
  assign n3629 = (n1747 & n1749) | (n1747 & n3628) | (n1749 & n3628);
  assign n3039 = n1740 | n1742;
  assign n3040 = (n1661 & n1740) | (n1661 & n3039) | (n1740 & n3039);
  assign n3041 = n1733 | n1735;
  assign n3042 = (n1733 & n2984) | (n1733 & n3041) | (n2984 & n3041);
  assign n3044 = n1698 | n1700;
  assign n3630 = n1585 | n1698;
  assign n3631 = (n1698 & n1700) | (n1698 & n3630) | (n1700 & n3630);
  assign n3632 = (n2957 & n3044) | (n2957 & n3631) | (n3044 & n3631);
  assign n3633 = (n1587 & n3044) | (n1587 & n3631) | (n3044 & n3631);
  assign n3634 = (n2921 & n3632) | (n2921 & n3633) | (n3632 & n3633);
  assign n1788 = x31 & x34;
  assign n1789 = n3613 & n1788;
  assign n1790 = n3613 | n1788;
  assign n1791 = ~n1789 & n1790;
  assign n3635 = n1677 | n1679;
  assign n3636 = (n1677 & n2990) | (n1677 & n3635) | (n2990 & n3635);
  assign n3051 = n1791 & n3636;
  assign n3637 = n1564 | n1677;
  assign n3638 = (n1677 & n1679) | (n1677 & n3637) | (n1679 & n3637);
  assign n3052 = n1791 & n3638;
  assign n3053 = (n3579 & n3051) | (n3579 & n3052) | (n3051 & n3052);
  assign n3054 = n1791 | n3636;
  assign n3055 = n1791 | n3638;
  assign n3056 = (n3579 & n3054) | (n3579 & n3055) | (n3054 & n3055);
  assign n1794 = ~n3053 & n3056;
  assign n1795 = x30 & x35;
  assign n1796 = n1794 & n1795;
  assign n1797 = n1794 | n1795;
  assign n1798 = ~n1796 & n1797;
  assign n3046 = n1684 | n1686;
  assign n3057 = n1798 & n3046;
  assign n3058 = n1684 & n1798;
  assign n3059 = (n3604 & n3057) | (n3604 & n3058) | (n3057 & n3058);
  assign n3060 = n1798 | n3046;
  assign n3061 = n1684 | n1798;
  assign n3062 = (n3604 & n3060) | (n3604 & n3061) | (n3060 & n3061);
  assign n1801 = ~n3059 & n3062;
  assign n1802 = x29 & x36;
  assign n1803 = n1801 & n1802;
  assign n1804 = n1801 | n1802;
  assign n1805 = ~n1803 & n1804;
  assign n3063 = n1691 & n1805;
  assign n3639 = (n1805 & n3008) | (n1805 & n3063) | (n3008 & n3063);
  assign n3640 = (n1805 & n3007) | (n1805 & n3063) | (n3007 & n3063);
  assign n3641 = (n3572 & n3639) | (n3572 & n3640) | (n3639 & n3640);
  assign n3065 = n1691 | n1805;
  assign n3642 = n3008 | n3065;
  assign n3643 = n3007 | n3065;
  assign n3644 = (n3572 & n3642) | (n3572 & n3643) | (n3642 & n3643);
  assign n1808 = ~n3641 & n3644;
  assign n1809 = x28 & x37;
  assign n1810 = n1808 & n1809;
  assign n1811 = n1808 | n1809;
  assign n1812 = ~n1810 & n1811;
  assign n1813 = n3634 & n1812;
  assign n1814 = n3634 | n1812;
  assign n1815 = ~n1813 & n1814;
  assign n1816 = x27 & x38;
  assign n1817 = n1815 & n1816;
  assign n1818 = n1815 | n1816;
  assign n1819 = ~n1817 & n1818;
  assign n3067 = n1705 & n1819;
  assign n3068 = (n1819 & n3018) | (n1819 & n3067) | (n3018 & n3067);
  assign n3069 = n1705 | n1819;
  assign n3070 = n3018 | n3069;
  assign n1822 = ~n3068 & n3070;
  assign n1823 = x26 & x39;
  assign n1824 = n1822 & n1823;
  assign n1825 = n1822 | n1823;
  assign n1826 = ~n1824 & n1825;
  assign n3071 = n1712 & n1826;
  assign n3072 = (n1826 & n3022) | (n1826 & n3071) | (n3022 & n3071);
  assign n3073 = n1712 | n1826;
  assign n3074 = n3022 | n3073;
  assign n1829 = ~n3072 & n3074;
  assign n1830 = x25 & x40;
  assign n1831 = n1829 & n1830;
  assign n1832 = n1829 | n1830;
  assign n1833 = ~n1831 & n1832;
  assign n3075 = n1719 & n1833;
  assign n3076 = (n1833 & n3026) | (n1833 & n3075) | (n3026 & n3075);
  assign n3077 = n1719 | n1833;
  assign n3078 = n3026 | n3077;
  assign n1836 = ~n3076 & n3078;
  assign n1837 = x24 & x41;
  assign n1838 = n1836 & n1837;
  assign n1839 = n1836 | n1837;
  assign n1840 = ~n1838 & n1839;
  assign n3079 = n1726 & n1840;
  assign n3080 = (n1840 & n3030) | (n1840 & n3079) | (n3030 & n3079);
  assign n3081 = n1726 | n1840;
  assign n3082 = n3030 | n3081;
  assign n1843 = ~n3080 & n3082;
  assign n1844 = x23 & x42;
  assign n1845 = n1843 & n1844;
  assign n1846 = n1843 | n1844;
  assign n1847 = ~n1845 & n1846;
  assign n1848 = n3042 & n1847;
  assign n1849 = n3042 | n1847;
  assign n1850 = ~n1848 & n1849;
  assign n1851 = x22 & x43;
  assign n1852 = n1850 & n1851;
  assign n1853 = n1850 | n1851;
  assign n1854 = ~n1852 & n1853;
  assign n1855 = n3040 & n1854;
  assign n1856 = n3040 | n1854;
  assign n1857 = ~n1855 & n1856;
  assign n1858 = x21 & x44;
  assign n1859 = n1857 & n1858;
  assign n1860 = n1857 | n1858;
  assign n1861 = ~n1859 & n1860;
  assign n1862 = n3629 & n1861;
  assign n1863 = n3629 | n1861;
  assign n1864 = ~n1862 & n1863;
  assign n1865 = x20 & x45;
  assign n1866 = n1864 & n1865;
  assign n1867 = n1864 | n1865;
  assign n1868 = ~n1866 & n1867;
  assign n1869 = n3038 & n1868;
  assign n1870 = n3038 | n1868;
  assign n1871 = ~n1869 & n1870;
  assign n1872 = x19 & x46;
  assign n1873 = n1871 & n1872;
  assign n1874 = n1871 | n1872;
  assign n1875 = ~n1873 & n1874;
  assign n1876 = n3036 & n1875;
  assign n1877 = n3036 | n1875;
  assign n1878 = ~n1876 & n1877;
  assign n1879 = x18 & x47;
  assign n1880 = n1878 & n1879;
  assign n1881 = n1878 | n1879;
  assign n1882 = ~n1880 & n1881;
  assign n1883 = n3034 & n1882;
  assign n1884 = n3034 | n1882;
  assign n1885 = ~n1883 & n1884;
  assign n3083 = n1880 | n3034;
  assign n3084 = (n1880 & n1882) | (n1880 & n3083) | (n1882 & n3083);
  assign n3085 = n1873 | n3036;
  assign n3086 = (n1873 & n1875) | (n1873 & n3085) | (n1875 & n3085);
  assign n3087 = n1866 | n3038;
  assign n3088 = (n1866 & n1868) | (n1866 & n3087) | (n1868 & n3087);
  assign n3089 = n1859 | n1861;
  assign n3090 = (n3629 & n1859) | (n3629 & n3089) | (n1859 & n3089);
  assign n3091 = n1852 | n1854;
  assign n3092 = (n1852 & n3040) | (n1852 & n3091) | (n3040 & n3091);
  assign n3093 = n1845 | n1847;
  assign n3094 = (n1845 & n3042) | (n1845 & n3093) | (n3042 & n3093);
  assign n3098 = n1803 | n1805;
  assign n3645 = n1691 | n1803;
  assign n3646 = (n1803 & n1805) | (n1803 & n3645) | (n1805 & n3645);
  assign n3647 = (n3008 & n3098) | (n3008 & n3646) | (n3098 & n3646);
  assign n3648 = (n3007 & n3098) | (n3007 & n3646) | (n3098 & n3646);
  assign n3649 = (n3572 & n3647) | (n3572 & n3648) | (n3647 & n3648);
  assign n1900 = x31 & x35;
  assign n3654 = n1788 & n1900;
  assign n3655 = n3613 & n3654;
  assign n11823 = (n1791 & n1900) | (n1791 & n3655) | (n1900 & n3655);
  assign n15523 = n1900 & n3654;
  assign n15524 = n3613 & n15523;
  assign n11825 = (n3636 & n11823) | (n3636 & n15524) | (n11823 & n15524);
  assign n11826 = (n3638 & n11823) | (n3638 & n15524) | (n11823 & n15524);
  assign n3658 = (n3579 & n11825) | (n3579 & n11826) | (n11825 & n11826);
  assign n3659 = n1788 | n1900;
  assign n3660 = (n1900 & n3613) | (n1900 & n3659) | (n3613 & n3659);
  assign n11827 = n1791 | n3660;
  assign n11828 = (n3636 & n3660) | (n3636 & n11827) | (n3660 & n11827);
  assign n11829 = (n3638 & n3660) | (n3638 & n11827) | (n3660 & n11827);
  assign n3663 = (n3579 & n11828) | (n3579 & n11829) | (n11828 & n11829);
  assign n1903 = ~n3658 & n3663;
  assign n3650 = n1796 | n1798;
  assign n3651 = (n1796 & n3046) | (n1796 & n3650) | (n3046 & n3650);
  assign n3664 = n1903 & n3651;
  assign n3652 = n1684 | n1796;
  assign n3653 = (n1796 & n1798) | (n1796 & n3652) | (n1798 & n3652);
  assign n3665 = n1903 & n3653;
  assign n3666 = (n3604 & n3664) | (n3604 & n3665) | (n3664 & n3665);
  assign n3667 = n1903 | n3651;
  assign n3668 = n1903 | n3653;
  assign n3669 = (n3604 & n3667) | (n3604 & n3668) | (n3667 & n3668);
  assign n1906 = ~n3666 & n3669;
  assign n1907 = x30 & x36;
  assign n1908 = n1906 & n1907;
  assign n1909 = n1906 | n1907;
  assign n1910 = ~n1908 & n1909;
  assign n1911 = n3649 & n1910;
  assign n1912 = n3649 | n1910;
  assign n1913 = ~n1911 & n1912;
  assign n1914 = x29 & x37;
  assign n1915 = n1913 & n1914;
  assign n1916 = n1913 | n1914;
  assign n1917 = ~n1915 & n1916;
  assign n3095 = n1810 | n1812;
  assign n3107 = n1917 & n3095;
  assign n3108 = n1810 & n1917;
  assign n3109 = (n3634 & n3107) | (n3634 & n3108) | (n3107 & n3108);
  assign n3110 = n1917 | n3095;
  assign n3111 = n1810 | n1917;
  assign n3112 = (n3634 & n3110) | (n3634 & n3111) | (n3110 & n3111);
  assign n1920 = ~n3109 & n3112;
  assign n1921 = x28 & x38;
  assign n1922 = n1920 & n1921;
  assign n1923 = n1920 | n1921;
  assign n1924 = ~n1922 & n1923;
  assign n3113 = n1817 & n1924;
  assign n3670 = (n1924 & n3067) | (n1924 & n3113) | (n3067 & n3113);
  assign n3671 = (n1819 & n1924) | (n1819 & n3113) | (n1924 & n3113);
  assign n3672 = (n3018 & n3670) | (n3018 & n3671) | (n3670 & n3671);
  assign n3115 = n1817 | n1924;
  assign n3673 = n3067 | n3115;
  assign n3674 = n1819 | n3115;
  assign n3675 = (n3018 & n3673) | (n3018 & n3674) | (n3673 & n3674);
  assign n1927 = ~n3672 & n3675;
  assign n1928 = x27 & x39;
  assign n1929 = n1927 & n1928;
  assign n1930 = n1927 | n1928;
  assign n1931 = ~n1929 & n1930;
  assign n3117 = n1824 & n1931;
  assign n3118 = (n1931 & n3072) | (n1931 & n3117) | (n3072 & n3117);
  assign n3119 = n1824 | n1931;
  assign n3120 = n3072 | n3119;
  assign n1934 = ~n3118 & n3120;
  assign n1935 = x26 & x40;
  assign n1936 = n1934 & n1935;
  assign n1937 = n1934 | n1935;
  assign n1938 = ~n1936 & n1937;
  assign n3121 = n1831 & n1938;
  assign n3122 = (n1938 & n3076) | (n1938 & n3121) | (n3076 & n3121);
  assign n3123 = n1831 | n1938;
  assign n3124 = n3076 | n3123;
  assign n1941 = ~n3122 & n3124;
  assign n1942 = x25 & x41;
  assign n1943 = n1941 & n1942;
  assign n1944 = n1941 | n1942;
  assign n1945 = ~n1943 & n1944;
  assign n3125 = n1838 & n1945;
  assign n3126 = (n1945 & n3080) | (n1945 & n3125) | (n3080 & n3125);
  assign n3127 = n1838 | n1945;
  assign n3128 = n3080 | n3127;
  assign n1948 = ~n3126 & n3128;
  assign n1949 = x24 & x42;
  assign n1950 = n1948 & n1949;
  assign n1951 = n1948 | n1949;
  assign n1952 = ~n1950 & n1951;
  assign n1953 = n3094 & n1952;
  assign n1954 = n3094 | n1952;
  assign n1955 = ~n1953 & n1954;
  assign n1956 = x23 & x43;
  assign n1957 = n1955 & n1956;
  assign n1958 = n1955 | n1956;
  assign n1959 = ~n1957 & n1958;
  assign n1960 = n3092 & n1959;
  assign n1961 = n3092 | n1959;
  assign n1962 = ~n1960 & n1961;
  assign n1963 = x22 & x44;
  assign n1964 = n1962 & n1963;
  assign n1965 = n1962 | n1963;
  assign n1966 = ~n1964 & n1965;
  assign n1967 = n3090 & n1966;
  assign n1968 = n3090 | n1966;
  assign n1969 = ~n1967 & n1968;
  assign n1970 = x21 & x45;
  assign n1971 = n1969 & n1970;
  assign n1972 = n1969 | n1970;
  assign n1973 = ~n1971 & n1972;
  assign n1974 = n3088 & n1973;
  assign n1975 = n3088 | n1973;
  assign n1976 = ~n1974 & n1975;
  assign n1977 = x20 & x46;
  assign n1978 = n1976 & n1977;
  assign n1979 = n1976 | n1977;
  assign n1980 = ~n1978 & n1979;
  assign n1981 = n3086 & n1980;
  assign n1982 = n3086 | n1980;
  assign n1983 = ~n1981 & n1982;
  assign n1984 = x19 & x47;
  assign n1985 = n1983 & n1984;
  assign n1986 = n1983 | n1984;
  assign n1987 = ~n1985 & n1986;
  assign n1988 = n3084 & n1987;
  assign n1989 = n3084 | n1987;
  assign n1990 = ~n1988 & n1989;
  assign n1991 = n1985 | n1988;
  assign n1992 = n1978 | n1981;
  assign n1993 = n1971 | n1974;
  assign n3129 = n1964 | n1966;
  assign n3130 = (n1964 & n3090) | (n1964 & n3129) | (n3090 & n3129);
  assign n3131 = n1957 | n1959;
  assign n3132 = (n1957 & n3092) | (n1957 & n3131) | (n3092 & n3131);
  assign n3133 = n1950 | n1952;
  assign n3134 = (n1950 & n3094) | (n1950 & n3133) | (n3094 & n3133);
  assign n3136 = n1922 | n1924;
  assign n3676 = n1817 | n1922;
  assign n3677 = (n1922 & n1924) | (n1922 & n3676) | (n1924 & n3676);
  assign n3678 = (n3067 & n3136) | (n3067 & n3677) | (n3136 & n3677);
  assign n3679 = (n1819 & n3136) | (n1819 & n3677) | (n3136 & n3677);
  assign n3680 = (n3018 & n3678) | (n3018 & n3679) | (n3678 & n3679);
  assign n2004 = x31 & x36;
  assign n66353 = n2004 & n3654;
  assign n66354 = n3613 & n66353;
  assign n49823 = n1900 & n2004;
  assign n49824 = (n1791 & n66354) | (n1791 & n49823) | (n66354 & n49823);
  assign n66355 = n3654 & n49823;
  assign n49826 = n3613 & n66355;
  assign n15527 = (n3636 & n49824) | (n3636 & n49826) | (n49824 & n49826);
  assign n15528 = (n3638 & n49824) | (n3638 & n49826) | (n49824 & n49826);
  assign n11832 = (n3579 & n15527) | (n3579 & n15528) | (n15527 & n15528);
  assign n3682 = (n1903 & n2004) | (n1903 & n11832) | (n2004 & n11832);
  assign n3683 = (n11832 & n3651) | (n11832 & n3682) | (n3651 & n3682);
  assign n3684 = (n11832 & n3653) | (n11832 & n3682) | (n3653 & n3682);
  assign n3685 = (n3604 & n3683) | (n3604 & n3684) | (n3683 & n3684);
  assign n66356 = n2004 | n3654;
  assign n66357 = (n2004 & n3613) | (n2004 & n66356) | (n3613 & n66356);
  assign n49828 = n1900 | n2004;
  assign n49829 = (n1791 & n66357) | (n1791 & n49828) | (n66357 & n49828);
  assign n66358 = (n2004 & n3654) | (n2004 & n49828) | (n3654 & n49828);
  assign n49831 = (n2004 & n3613) | (n2004 & n66358) | (n3613 & n66358);
  assign n15531 = (n3636 & n49829) | (n3636 & n49831) | (n49829 & n49831);
  assign n15532 = (n3638 & n49829) | (n3638 & n49831) | (n49829 & n49831);
  assign n11835 = (n3579 & n15531) | (n3579 & n15532) | (n15531 & n15532);
  assign n3687 = n1903 | n11835;
  assign n3688 = (n11835 & n3651) | (n11835 & n3687) | (n3651 & n3687);
  assign n3689 = (n11835 & n3653) | (n11835 & n3687) | (n3653 & n3687);
  assign n3690 = (n3604 & n3688) | (n3604 & n3689) | (n3688 & n3689);
  assign n2007 = ~n3685 & n3690;
  assign n3149 = n1908 & n2007;
  assign n3691 = (n1910 & n2007) | (n1910 & n3149) | (n2007 & n3149);
  assign n3150 = (n3649 & n3691) | (n3649 & n3149) | (n3691 & n3149);
  assign n3152 = n1908 | n2007;
  assign n3692 = n1910 | n3152;
  assign n3153 = (n3649 & n3692) | (n3649 & n3152) | (n3692 & n3152);
  assign n2010 = ~n3150 & n3153;
  assign n2011 = x30 & x37;
  assign n2012 = n2010 & n2011;
  assign n2013 = n2010 | n2011;
  assign n2014 = ~n2012 & n2013;
  assign n3154 = n1915 & n2014;
  assign n3693 = (n2014 & n3108) | (n2014 & n3154) | (n3108 & n3154);
  assign n3694 = (n2014 & n3107) | (n2014 & n3154) | (n3107 & n3154);
  assign n3695 = (n3634 & n3693) | (n3634 & n3694) | (n3693 & n3694);
  assign n3156 = n1915 | n2014;
  assign n3696 = n3108 | n3156;
  assign n3697 = n3107 | n3156;
  assign n3698 = (n3634 & n3696) | (n3634 & n3697) | (n3696 & n3697);
  assign n2017 = ~n3695 & n3698;
  assign n2018 = x29 & x38;
  assign n2019 = n2017 & n2018;
  assign n2020 = n2017 | n2018;
  assign n2021 = ~n2019 & n2020;
  assign n2022 = n3680 & n2021;
  assign n2023 = n3680 | n2021;
  assign n2024 = ~n2022 & n2023;
  assign n2025 = x28 & x39;
  assign n2026 = n2024 & n2025;
  assign n2027 = n2024 | n2025;
  assign n2028 = ~n2026 & n2027;
  assign n3158 = n1929 & n2028;
  assign n3159 = (n2028 & n3118) | (n2028 & n3158) | (n3118 & n3158);
  assign n3160 = n1929 | n2028;
  assign n3161 = n3118 | n3160;
  assign n2031 = ~n3159 & n3161;
  assign n2032 = x27 & x40;
  assign n2033 = n2031 & n2032;
  assign n2034 = n2031 | n2032;
  assign n2035 = ~n2033 & n2034;
  assign n3162 = n1936 & n2035;
  assign n3163 = (n2035 & n3122) | (n2035 & n3162) | (n3122 & n3162);
  assign n3164 = n1936 | n2035;
  assign n3165 = n3122 | n3164;
  assign n2038 = ~n3163 & n3165;
  assign n2039 = x26 & x41;
  assign n2040 = n2038 & n2039;
  assign n2041 = n2038 | n2039;
  assign n2042 = ~n2040 & n2041;
  assign n3166 = n1943 & n2042;
  assign n3167 = (n2042 & n3126) | (n2042 & n3166) | (n3126 & n3166);
  assign n3168 = n1943 | n2042;
  assign n3169 = n3126 | n3168;
  assign n2045 = ~n3167 & n3169;
  assign n2046 = x25 & x42;
  assign n2047 = n2045 & n2046;
  assign n2048 = n2045 | n2046;
  assign n2049 = ~n2047 & n2048;
  assign n2050 = n3134 & n2049;
  assign n2051 = n3134 | n2049;
  assign n2052 = ~n2050 & n2051;
  assign n2053 = x24 & x43;
  assign n2054 = n2052 & n2053;
  assign n2055 = n2052 | n2053;
  assign n2056 = ~n2054 & n2055;
  assign n2057 = n3132 & n2056;
  assign n2058 = n3132 | n2056;
  assign n2059 = ~n2057 & n2058;
  assign n2060 = x23 & x44;
  assign n2061 = n2059 & n2060;
  assign n2062 = n2059 | n2060;
  assign n2063 = ~n2061 & n2062;
  assign n2064 = n3130 & n2063;
  assign n2065 = n3130 | n2063;
  assign n2066 = ~n2064 & n2065;
  assign n2067 = x22 & x45;
  assign n2068 = n2066 & n2067;
  assign n2069 = n2066 | n2067;
  assign n2070 = ~n2068 & n2069;
  assign n2071 = n1993 & n2070;
  assign n2072 = n1993 | n2070;
  assign n2073 = ~n2071 & n2072;
  assign n2074 = x21 & x46;
  assign n2075 = n2073 & n2074;
  assign n2076 = n2073 | n2074;
  assign n2077 = ~n2075 & n2076;
  assign n2078 = n1992 & n2077;
  assign n2079 = n1992 | n2077;
  assign n2080 = ~n2078 & n2079;
  assign n2081 = x20 & x47;
  assign n2082 = n2080 & n2081;
  assign n2083 = n2080 | n2081;
  assign n2084 = ~n2082 & n2083;
  assign n2085 = n1991 & n2084;
  assign n2086 = n1991 | n2084;
  assign n2087 = ~n2085 & n2086;
  assign n2088 = n2082 | n2085;
  assign n2089 = n2075 | n2078;
  assign n3170 = n2068 | n2070;
  assign n3171 = (n1993 & n2068) | (n1993 & n3170) | (n2068 & n3170);
  assign n3172 = n2061 | n2063;
  assign n3173 = (n2061 & n3130) | (n2061 & n3172) | (n3130 & n3172);
  assign n3174 = n2054 | n2056;
  assign n3175 = (n2054 & n3132) | (n2054 & n3174) | (n3132 & n3174);
  assign n3176 = n2047 | n2049;
  assign n3177 = (n2047 & n3134) | (n2047 & n3176) | (n3134 & n3176);
  assign n3181 = n2012 | n2014;
  assign n3699 = n1915 | n2012;
  assign n3700 = (n2012 & n2014) | (n2012 & n3699) | (n2014 & n3699);
  assign n3701 = (n3108 & n3181) | (n3108 & n3700) | (n3181 & n3700);
  assign n3702 = (n3107 & n3181) | (n3107 & n3700) | (n3181 & n3700);
  assign n3703 = (n3634 & n3701) | (n3634 & n3702) | (n3701 & n3702);
  assign n2100 = x31 & x37;
  assign n3183 = n2100 & n3685;
  assign n3704 = (n2100 & n3183) | (n2100 & n3691) | (n3183 & n3691);
  assign n11836 = (n2007 & n2100) | (n2007 & n3183) | (n2100 & n3183);
  assign n15533 = n2100 & n3685;
  assign n11838 = (n1908 & n11836) | (n1908 & n15533) | (n11836 & n15533);
  assign n3706 = (n3649 & n3704) | (n3649 & n11838) | (n3704 & n11838);
  assign n3185 = n2100 | n3685;
  assign n3707 = n3185 | n3691;
  assign n11839 = n2007 | n3185;
  assign n11840 = (n1908 & n3185) | (n1908 & n11839) | (n3185 & n11839);
  assign n3709 = (n3649 & n3707) | (n3649 & n11840) | (n3707 & n11840);
  assign n2103 = ~n3706 & n3709;
  assign n2104 = n3703 & n2103;
  assign n2105 = n3703 | n2103;
  assign n2106 = ~n2104 & n2105;
  assign n2107 = x30 & x38;
  assign n2108 = n2106 & n2107;
  assign n2109 = n2106 | n2107;
  assign n2110 = ~n2108 & n2109;
  assign n3178 = n2019 | n2021;
  assign n3187 = n2110 & n3178;
  assign n3188 = n2019 & n2110;
  assign n3189 = (n3680 & n3187) | (n3680 & n3188) | (n3187 & n3188);
  assign n3190 = n2110 | n3178;
  assign n3191 = n2019 | n2110;
  assign n3192 = (n3680 & n3190) | (n3680 & n3191) | (n3190 & n3191);
  assign n2113 = ~n3189 & n3192;
  assign n2114 = x29 & x39;
  assign n2115 = n2113 & n2114;
  assign n2116 = n2113 | n2114;
  assign n2117 = ~n2115 & n2116;
  assign n3193 = n2026 & n2117;
  assign n3710 = (n2117 & n3158) | (n2117 & n3193) | (n3158 & n3193);
  assign n3711 = (n2028 & n2117) | (n2028 & n3193) | (n2117 & n3193);
  assign n3712 = (n3118 & n3710) | (n3118 & n3711) | (n3710 & n3711);
  assign n3195 = n2026 | n2117;
  assign n3713 = n3158 | n3195;
  assign n3714 = n2028 | n3195;
  assign n3715 = (n3118 & n3713) | (n3118 & n3714) | (n3713 & n3714);
  assign n2120 = ~n3712 & n3715;
  assign n2121 = x28 & x40;
  assign n2122 = n2120 & n2121;
  assign n2123 = n2120 | n2121;
  assign n2124 = ~n2122 & n2123;
  assign n3197 = n2033 & n2124;
  assign n3198 = (n2124 & n3163) | (n2124 & n3197) | (n3163 & n3197);
  assign n3199 = n2033 | n2124;
  assign n3200 = n3163 | n3199;
  assign n2127 = ~n3198 & n3200;
  assign n2128 = x27 & x41;
  assign n2129 = n2127 & n2128;
  assign n2130 = n2127 | n2128;
  assign n2131 = ~n2129 & n2130;
  assign n3201 = n2040 & n2131;
  assign n3202 = (n2131 & n3167) | (n2131 & n3201) | (n3167 & n3201);
  assign n3203 = n2040 | n2131;
  assign n3204 = n3167 | n3203;
  assign n2134 = ~n3202 & n3204;
  assign n2135 = x26 & x42;
  assign n2136 = n2134 & n2135;
  assign n2137 = n2134 | n2135;
  assign n2138 = ~n2136 & n2137;
  assign n2139 = n3177 & n2138;
  assign n2140 = n3177 | n2138;
  assign n2141 = ~n2139 & n2140;
  assign n2142 = x25 & x43;
  assign n2143 = n2141 & n2142;
  assign n2144 = n2141 | n2142;
  assign n2145 = ~n2143 & n2144;
  assign n2146 = n3175 & n2145;
  assign n2147 = n3175 | n2145;
  assign n2148 = ~n2146 & n2147;
  assign n2149 = x24 & x44;
  assign n2150 = n2148 & n2149;
  assign n2151 = n2148 | n2149;
  assign n2152 = ~n2150 & n2151;
  assign n2153 = n3173 & n2152;
  assign n2154 = n3173 | n2152;
  assign n2155 = ~n2153 & n2154;
  assign n2156 = x23 & x45;
  assign n2157 = n2155 & n2156;
  assign n2158 = n2155 | n2156;
  assign n2159 = ~n2157 & n2158;
  assign n2160 = n3171 & n2159;
  assign n2161 = n3171 | n2159;
  assign n2162 = ~n2160 & n2161;
  assign n2163 = x22 & x46;
  assign n2164 = n2162 & n2163;
  assign n2165 = n2162 | n2163;
  assign n2166 = ~n2164 & n2165;
  assign n2167 = n2089 & n2166;
  assign n2168 = n2089 | n2166;
  assign n2169 = ~n2167 & n2168;
  assign n2170 = x21 & x47;
  assign n2171 = n2169 & n2170;
  assign n2172 = n2169 | n2170;
  assign n2173 = ~n2171 & n2172;
  assign n2174 = n2088 & n2173;
  assign n2175 = n2088 | n2173;
  assign n2176 = ~n2174 & n2175;
  assign n2177 = n2171 | n2174;
  assign n3205 = n2164 | n2166;
  assign n3206 = (n2089 & n2164) | (n2089 & n3205) | (n2164 & n3205);
  assign n3207 = n2157 | n2159;
  assign n3208 = (n2157 & n3171) | (n2157 & n3207) | (n3171 & n3207);
  assign n3209 = n2150 | n2152;
  assign n3210 = (n2150 & n3173) | (n2150 & n3209) | (n3173 & n3209);
  assign n3211 = n2143 | n2145;
  assign n3212 = (n2143 & n3175) | (n2143 & n3211) | (n3175 & n3211);
  assign n3213 = n2136 | n2138;
  assign n3214 = (n2136 & n3177) | (n2136 & n3213) | (n3177 & n3213);
  assign n3216 = n2115 | n2117;
  assign n3716 = n2026 | n2115;
  assign n3717 = (n2115 & n2117) | (n2115 & n3716) | (n2117 & n3716);
  assign n3718 = (n3158 & n3216) | (n3158 & n3717) | (n3216 & n3717);
  assign n3719 = (n2028 & n3216) | (n2028 & n3717) | (n3216 & n3717);
  assign n3720 = (n3118 & n3718) | (n3118 & n3719) | (n3718 & n3719);
  assign n2188 = x31 & x38;
  assign n11844 = n2100 & n2188;
  assign n15534 = n3685 & n11844;
  assign n11845 = (n3691 & n15534) | (n3691 & n11844) | (n15534 & n11844);
  assign n11841 = n2188 & n11838;
  assign n11842 = (n3649 & n11845) | (n3649 & n11841) | (n11845 & n11841);
  assign n3722 = (n2103 & n2188) | (n2103 & n11842) | (n2188 & n11842);
  assign n3724 = n2188 & n11838;
  assign n3725 = (n3649 & n11845) | (n3649 & n3724) | (n11845 & n3724);
  assign n3222 = (n3703 & n3722) | (n3703 & n3725) | (n3722 & n3725);
  assign n11849 = n2100 | n2188;
  assign n15535 = (n2188 & n3685) | (n2188 & n11849) | (n3685 & n11849);
  assign n11850 = (n3691 & n15535) | (n3691 & n11849) | (n15535 & n11849);
  assign n11846 = n2188 | n11838;
  assign n11847 = (n3649 & n11850) | (n3649 & n11846) | (n11850 & n11846);
  assign n3727 = n2103 | n11847;
  assign n3729 = n2188 | n11838;
  assign n3730 = (n3649 & n11850) | (n3649 & n3729) | (n11850 & n3729);
  assign n3225 = (n3703 & n3727) | (n3703 & n3730) | (n3727 & n3730);
  assign n2191 = ~n3222 & n3225;
  assign n3226 = n2108 & n2191;
  assign n3731 = (n2191 & n3188) | (n2191 & n3226) | (n3188 & n3226);
  assign n3732 = (n2191 & n3187) | (n2191 & n3226) | (n3187 & n3226);
  assign n3733 = (n3680 & n3731) | (n3680 & n3732) | (n3731 & n3732);
  assign n3228 = n2108 | n2191;
  assign n3734 = n3188 | n3228;
  assign n3735 = n3187 | n3228;
  assign n3736 = (n3680 & n3734) | (n3680 & n3735) | (n3734 & n3735);
  assign n2194 = ~n3733 & n3736;
  assign n2195 = x30 & x39;
  assign n2196 = n2194 & n2195;
  assign n2197 = n2194 | n2195;
  assign n2198 = ~n2196 & n2197;
  assign n2199 = n3720 & n2198;
  assign n2200 = n3720 | n2198;
  assign n2201 = ~n2199 & n2200;
  assign n2202 = x29 & x40;
  assign n2203 = n2201 & n2202;
  assign n2204 = n2201 | n2202;
  assign n2205 = ~n2203 & n2204;
  assign n3230 = n2122 & n2205;
  assign n3231 = (n2205 & n3198) | (n2205 & n3230) | (n3198 & n3230);
  assign n3232 = n2122 | n2205;
  assign n3233 = n3198 | n3232;
  assign n2208 = ~n3231 & n3233;
  assign n2209 = x28 & x41;
  assign n2210 = n2208 & n2209;
  assign n2211 = n2208 | n2209;
  assign n2212 = ~n2210 & n2211;
  assign n3234 = n2129 & n2212;
  assign n3235 = (n2212 & n3202) | (n2212 & n3234) | (n3202 & n3234);
  assign n3236 = n2129 | n2212;
  assign n3237 = n3202 | n3236;
  assign n2215 = ~n3235 & n3237;
  assign n2216 = x27 & x42;
  assign n2217 = n2215 & n2216;
  assign n2218 = n2215 | n2216;
  assign n2219 = ~n2217 & n2218;
  assign n2220 = n3214 & n2219;
  assign n2221 = n3214 | n2219;
  assign n2222 = ~n2220 & n2221;
  assign n2223 = x26 & x43;
  assign n2224 = n2222 & n2223;
  assign n2225 = n2222 | n2223;
  assign n2226 = ~n2224 & n2225;
  assign n2227 = n3212 & n2226;
  assign n2228 = n3212 | n2226;
  assign n2229 = ~n2227 & n2228;
  assign n2230 = x25 & x44;
  assign n2231 = n2229 & n2230;
  assign n2232 = n2229 | n2230;
  assign n2233 = ~n2231 & n2232;
  assign n2234 = n3210 & n2233;
  assign n2235 = n3210 | n2233;
  assign n2236 = ~n2234 & n2235;
  assign n2237 = x24 & x45;
  assign n2238 = n2236 & n2237;
  assign n2239 = n2236 | n2237;
  assign n2240 = ~n2238 & n2239;
  assign n2241 = n3208 & n2240;
  assign n2242 = n3208 | n2240;
  assign n2243 = ~n2241 & n2242;
  assign n2244 = x23 & x46;
  assign n2245 = n2243 & n2244;
  assign n2246 = n2243 | n2244;
  assign n2247 = ~n2245 & n2246;
  assign n2248 = n3206 & n2247;
  assign n2249 = n3206 | n2247;
  assign n2250 = ~n2248 & n2249;
  assign n2251 = x22 & x47;
  assign n2252 = n2250 & n2251;
  assign n2253 = n2250 | n2251;
  assign n2254 = ~n2252 & n2253;
  assign n2255 = n2177 & n2254;
  assign n2256 = n2177 | n2254;
  assign n2257 = ~n2255 & n2256;
  assign n3238 = n2252 | n2254;
  assign n3239 = (n2177 & n2252) | (n2177 & n3238) | (n2252 & n3238);
  assign n3240 = n2245 | n2247;
  assign n3241 = (n2245 & n3206) | (n2245 & n3240) | (n3206 & n3240);
  assign n3242 = n2238 | n2240;
  assign n3243 = (n2238 & n3208) | (n2238 & n3242) | (n3208 & n3242);
  assign n3244 = n2231 | n2233;
  assign n3245 = (n2231 & n3210) | (n2231 & n3244) | (n3210 & n3244);
  assign n3246 = n2224 | n2226;
  assign n3247 = (n2224 & n3212) | (n2224 & n3246) | (n3212 & n3246);
  assign n3248 = n2217 | n2219;
  assign n3249 = (n2217 & n3214) | (n2217 & n3248) | (n3214 & n3248);
  assign n2268 = x31 & x39;
  assign n3253 = n2191 | n3222;
  assign n3737 = (n2108 & n3222) | (n2108 & n3253) | (n3222 & n3253);
  assign n3255 = n2268 & n3737;
  assign n49835 = n2268 & n11844;
  assign n66359 = n3685 & n49835;
  assign n49836 = (n3691 & n66359) | (n3691 & n49835) | (n66359 & n49835);
  assign n15537 = n2188 & n2268;
  assign n49837 = n11838 & n15537;
  assign n49833 = (n3649 & n49836) | (n3649 & n49837) | (n49836 & n49837);
  assign n15538 = (n2103 & n49833) | (n2103 & n15537) | (n49833 & n15537);
  assign n15541 = (n3649 & n49836) | (n3649 & n49837) | (n49836 & n49837);
  assign n11853 = (n3703 & n15538) | (n3703 & n15541) | (n15538 & n15541);
  assign n3739 = (n2191 & n2268) | (n2191 & n11853) | (n2268 & n11853);
  assign n3740 = (n3188 & n3255) | (n3188 & n3739) | (n3255 & n3739);
  assign n3741 = (n3187 & n3255) | (n3187 & n3739) | (n3255 & n3739);
  assign n3742 = (n3680 & n3740) | (n3680 & n3741) | (n3740 & n3741);
  assign n3258 = n2268 | n3737;
  assign n49841 = n2268 | n11844;
  assign n66360 = (n2268 & n3685) | (n2268 & n49841) | (n3685 & n49841);
  assign n49842 = (n3691 & n66360) | (n3691 & n49841) | (n66360 & n49841);
  assign n15543 = n2188 | n2268;
  assign n49843 = (n2268 & n11838) | (n2268 & n15543) | (n11838 & n15543);
  assign n49839 = (n3649 & n49842) | (n3649 & n49843) | (n49842 & n49843);
  assign n15544 = (n2103 & n49839) | (n2103 & n15543) | (n49839 & n15543);
  assign n15547 = (n3649 & n49842) | (n3649 & n49843) | (n49842 & n49843);
  assign n11856 = (n3703 & n15544) | (n3703 & n15547) | (n15544 & n15547);
  assign n3744 = n2191 | n11856;
  assign n3745 = (n3188 & n3258) | (n3188 & n3744) | (n3258 & n3744);
  assign n3746 = (n3187 & n3258) | (n3187 & n3744) | (n3258 & n3744);
  assign n3747 = (n3680 & n3745) | (n3680 & n3746) | (n3745 & n3746);
  assign n2271 = ~n3742 & n3747;
  assign n3262 = n2196 & n2271;
  assign n3748 = (n2198 & n2271) | (n2198 & n3262) | (n2271 & n3262);
  assign n3263 = (n3720 & n3748) | (n3720 & n3262) | (n3748 & n3262);
  assign n3265 = n2196 | n2271;
  assign n3749 = n2198 | n3265;
  assign n3266 = (n3720 & n3749) | (n3720 & n3265) | (n3749 & n3265);
  assign n2274 = ~n3263 & n3266;
  assign n2275 = x30 & x40;
  assign n2276 = n2274 & n2275;
  assign n2277 = n2274 | n2275;
  assign n2278 = ~n2276 & n2277;
  assign n3267 = n2203 & n2278;
  assign n3750 = (n2278 & n3230) | (n2278 & n3267) | (n3230 & n3267);
  assign n3751 = (n2205 & n2278) | (n2205 & n3267) | (n2278 & n3267);
  assign n3752 = (n3198 & n3750) | (n3198 & n3751) | (n3750 & n3751);
  assign n3269 = n2203 | n2278;
  assign n3753 = n3230 | n3269;
  assign n3754 = n2205 | n3269;
  assign n3755 = (n3198 & n3753) | (n3198 & n3754) | (n3753 & n3754);
  assign n2281 = ~n3752 & n3755;
  assign n2282 = x29 & x41;
  assign n2283 = n2281 & n2282;
  assign n2284 = n2281 | n2282;
  assign n2285 = ~n2283 & n2284;
  assign n3271 = n2210 & n2285;
  assign n3272 = (n2285 & n3235) | (n2285 & n3271) | (n3235 & n3271);
  assign n3273 = n2210 | n2285;
  assign n3274 = n3235 | n3273;
  assign n2288 = ~n3272 & n3274;
  assign n2289 = x28 & x42;
  assign n2290 = n2288 & n2289;
  assign n2291 = n2288 | n2289;
  assign n2292 = ~n2290 & n2291;
  assign n2293 = n3249 & n2292;
  assign n2294 = n3249 | n2292;
  assign n2295 = ~n2293 & n2294;
  assign n2296 = x27 & x43;
  assign n2297 = n2295 & n2296;
  assign n2298 = n2295 | n2296;
  assign n2299 = ~n2297 & n2298;
  assign n2300 = n3247 & n2299;
  assign n2301 = n3247 | n2299;
  assign n2302 = ~n2300 & n2301;
  assign n2303 = x26 & x44;
  assign n2304 = n2302 & n2303;
  assign n2305 = n2302 | n2303;
  assign n2306 = ~n2304 & n2305;
  assign n2307 = n3245 & n2306;
  assign n2308 = n3245 | n2306;
  assign n2309 = ~n2307 & n2308;
  assign n2310 = x25 & x45;
  assign n2311 = n2309 & n2310;
  assign n2312 = n2309 | n2310;
  assign n2313 = ~n2311 & n2312;
  assign n2314 = n3243 & n2313;
  assign n2315 = n3243 | n2313;
  assign n2316 = ~n2314 & n2315;
  assign n2317 = x24 & x46;
  assign n2318 = n2316 & n2317;
  assign n2319 = n2316 | n2317;
  assign n2320 = ~n2318 & n2319;
  assign n2321 = n3241 & n2320;
  assign n2322 = n3241 | n2320;
  assign n2323 = ~n2321 & n2322;
  assign n2324 = x23 & x47;
  assign n2325 = n2323 & n2324;
  assign n2326 = n2323 | n2324;
  assign n2327 = ~n2325 & n2326;
  assign n2328 = n3239 & n2327;
  assign n2329 = n3239 | n2327;
  assign n2330 = ~n2328 & n2329;
  assign n3275 = n2325 | n2327;
  assign n3276 = (n2325 & n3239) | (n2325 & n3275) | (n3239 & n3275);
  assign n3277 = n2318 | n2320;
  assign n3278 = (n2318 & n3241) | (n2318 & n3277) | (n3241 & n3277);
  assign n3279 = n2311 | n2313;
  assign n3280 = (n2311 & n3243) | (n2311 & n3279) | (n3243 & n3279);
  assign n3281 = n2304 | n2306;
  assign n3282 = (n2304 & n3245) | (n2304 & n3281) | (n3245 & n3281);
  assign n3283 = n2297 | n2299;
  assign n3284 = (n2297 & n3247) | (n2297 & n3283) | (n3247 & n3283);
  assign n3285 = n2290 | n2292;
  assign n3286 = (n2290 & n3249) | (n2290 & n3285) | (n3249 & n3285);
  assign n3288 = n2276 | n2278;
  assign n3756 = n2203 | n2276;
  assign n3757 = (n2276 & n2278) | (n2276 & n3756) | (n2278 & n3756);
  assign n3758 = (n3230 & n3288) | (n3230 & n3757) | (n3288 & n3757);
  assign n3759 = (n2205 & n3288) | (n2205 & n3757) | (n3288 & n3757);
  assign n3760 = (n3198 & n3758) | (n3198 & n3759) | (n3758 & n3759);
  assign n2340 = x31 & x40;
  assign n3290 = n2340 & n3742;
  assign n3761 = (n2340 & n3290) | (n2340 & n3748) | (n3290 & n3748);
  assign n11857 = (n2271 & n2340) | (n2271 & n3290) | (n2340 & n3290);
  assign n15548 = n2340 & n3742;
  assign n11859 = (n2196 & n11857) | (n2196 & n15548) | (n11857 & n15548);
  assign n3763 = (n3720 & n3761) | (n3720 & n11859) | (n3761 & n11859);
  assign n3292 = n2340 | n3742;
  assign n3764 = n3292 | n3748;
  assign n11860 = n2271 | n3292;
  assign n11861 = (n2196 & n3292) | (n2196 & n11860) | (n3292 & n11860);
  assign n3766 = (n3720 & n3764) | (n3720 & n11861) | (n3764 & n11861);
  assign n2343 = ~n3763 & n3766;
  assign n2344 = n3760 & n2343;
  assign n2345 = n3760 | n2343;
  assign n2346 = ~n2344 & n2345;
  assign n2347 = x30 & x41;
  assign n2348 = n2346 & n2347;
  assign n2349 = n2346 | n2347;
  assign n2350 = ~n2348 & n2349;
  assign n3294 = n2283 & n2350;
  assign n3295 = (n2350 & n3272) | (n2350 & n3294) | (n3272 & n3294);
  assign n3296 = n2283 | n2350;
  assign n3297 = n3272 | n3296;
  assign n2353 = ~n3295 & n3297;
  assign n2354 = x29 & x42;
  assign n2355 = n2353 & n2354;
  assign n2356 = n2353 | n2354;
  assign n2357 = ~n2355 & n2356;
  assign n2358 = n3286 & n2357;
  assign n2359 = n3286 | n2357;
  assign n2360 = ~n2358 & n2359;
  assign n2361 = x28 & x43;
  assign n2362 = n2360 & n2361;
  assign n2363 = n2360 | n2361;
  assign n2364 = ~n2362 & n2363;
  assign n2365 = n3284 & n2364;
  assign n2366 = n3284 | n2364;
  assign n2367 = ~n2365 & n2366;
  assign n2368 = x27 & x44;
  assign n2369 = n2367 & n2368;
  assign n2370 = n2367 | n2368;
  assign n2371 = ~n2369 & n2370;
  assign n2372 = n3282 & n2371;
  assign n2373 = n3282 | n2371;
  assign n2374 = ~n2372 & n2373;
  assign n2375 = x26 & x45;
  assign n2376 = n2374 & n2375;
  assign n2377 = n2374 | n2375;
  assign n2378 = ~n2376 & n2377;
  assign n2379 = n3280 & n2378;
  assign n2380 = n3280 | n2378;
  assign n2381 = ~n2379 & n2380;
  assign n2382 = x25 & x46;
  assign n2383 = n2381 & n2382;
  assign n2384 = n2381 | n2382;
  assign n2385 = ~n2383 & n2384;
  assign n2386 = n3278 & n2385;
  assign n2387 = n3278 | n2385;
  assign n2388 = ~n2386 & n2387;
  assign n2389 = x24 & x47;
  assign n2390 = n2388 & n2389;
  assign n2391 = n2388 | n2389;
  assign n2392 = ~n2390 & n2391;
  assign n2393 = n3276 & n2392;
  assign n2394 = n3276 | n2392;
  assign n2395 = ~n2393 & n2394;
  assign n3298 = n2390 | n2392;
  assign n3299 = (n2390 & n3276) | (n2390 & n3298) | (n3276 & n3298);
  assign n3300 = n2383 | n2385;
  assign n3301 = (n2383 & n3278) | (n2383 & n3300) | (n3278 & n3300);
  assign n3302 = n2376 | n2378;
  assign n3303 = (n2376 & n3280) | (n2376 & n3302) | (n3280 & n3302);
  assign n3304 = n2369 | n2371;
  assign n3305 = (n2369 & n3282) | (n2369 & n3304) | (n3282 & n3304);
  assign n3306 = n2362 | n2364;
  assign n3307 = (n2362 & n3284) | (n2362 & n3306) | (n3284 & n3306);
  assign n3308 = n2355 | n2357;
  assign n3309 = (n2355 & n3286) | (n2355 & n3308) | (n3286 & n3308);
  assign n2404 = x31 & x41;
  assign n11865 = n2340 & n2404;
  assign n15549 = n3742 & n11865;
  assign n11866 = (n3748 & n15549) | (n3748 & n11865) | (n15549 & n11865);
  assign n11862 = n2404 & n11859;
  assign n11863 = (n3720 & n11866) | (n3720 & n11862) | (n11866 & n11862);
  assign n3768 = (n2343 & n2404) | (n2343 & n11863) | (n2404 & n11863);
  assign n3770 = n2404 & n11859;
  assign n3771 = (n3720 & n11866) | (n3720 & n3770) | (n11866 & n3770);
  assign n3314 = (n3760 & n3768) | (n3760 & n3771) | (n3768 & n3771);
  assign n11870 = n2340 | n2404;
  assign n15550 = (n2404 & n3742) | (n2404 & n11870) | (n3742 & n11870);
  assign n11871 = (n3748 & n15550) | (n3748 & n11870) | (n15550 & n11870);
  assign n11867 = n2404 | n11859;
  assign n11868 = (n3720 & n11871) | (n3720 & n11867) | (n11871 & n11867);
  assign n3773 = n2343 | n11868;
  assign n3775 = n2404 | n11859;
  assign n3776 = (n3720 & n11871) | (n3720 & n3775) | (n11871 & n3775);
  assign n3317 = (n3760 & n3773) | (n3760 & n3776) | (n3773 & n3776);
  assign n2407 = ~n3314 & n3317;
  assign n3318 = n2348 & n2407;
  assign n3777 = (n2407 & n3294) | (n2407 & n3318) | (n3294 & n3318);
  assign n3778 = (n2350 & n2407) | (n2350 & n3318) | (n2407 & n3318);
  assign n3779 = (n3272 & n3777) | (n3272 & n3778) | (n3777 & n3778);
  assign n3320 = n2348 | n2407;
  assign n3780 = n3294 | n3320;
  assign n3781 = n2350 | n3320;
  assign n3782 = (n3272 & n3780) | (n3272 & n3781) | (n3780 & n3781);
  assign n2410 = ~n3779 & n3782;
  assign n2411 = x30 & x42;
  assign n2412 = n2410 & n2411;
  assign n2413 = n2410 | n2411;
  assign n2414 = ~n2412 & n2413;
  assign n2415 = n3309 & n2414;
  assign n2416 = n3309 | n2414;
  assign n2417 = ~n2415 & n2416;
  assign n2418 = x29 & x43;
  assign n2419 = n2417 & n2418;
  assign n2420 = n2417 | n2418;
  assign n2421 = ~n2419 & n2420;
  assign n2422 = n3307 & n2421;
  assign n2423 = n3307 | n2421;
  assign n2424 = ~n2422 & n2423;
  assign n2425 = x28 & x44;
  assign n2426 = n2424 & n2425;
  assign n2427 = n2424 | n2425;
  assign n2428 = ~n2426 & n2427;
  assign n2429 = n3305 & n2428;
  assign n2430 = n3305 | n2428;
  assign n2431 = ~n2429 & n2430;
  assign n2432 = x27 & x45;
  assign n2433 = n2431 & n2432;
  assign n2434 = n2431 | n2432;
  assign n2435 = ~n2433 & n2434;
  assign n2436 = n3303 & n2435;
  assign n2437 = n3303 | n2435;
  assign n2438 = ~n2436 & n2437;
  assign n2439 = x26 & x46;
  assign n2440 = n2438 & n2439;
  assign n2441 = n2438 | n2439;
  assign n2442 = ~n2440 & n2441;
  assign n2443 = n3301 & n2442;
  assign n2444 = n3301 | n2442;
  assign n2445 = ~n2443 & n2444;
  assign n2446 = x25 & x47;
  assign n2447 = n2445 & n2446;
  assign n2448 = n2445 | n2446;
  assign n2449 = ~n2447 & n2448;
  assign n2450 = n3299 & n2449;
  assign n2451 = n3299 | n2449;
  assign n2452 = ~n2450 & n2451;
  assign n3322 = n2447 | n2449;
  assign n3323 = (n2447 & n3299) | (n2447 & n3322) | (n3299 & n3322);
  assign n3324 = n2440 | n2442;
  assign n3325 = (n2440 & n3301) | (n2440 & n3324) | (n3301 & n3324);
  assign n3326 = n2433 | n2435;
  assign n3327 = (n2433 & n3303) | (n2433 & n3326) | (n3303 & n3326);
  assign n3328 = n2426 | n2428;
  assign n3329 = (n2426 & n3305) | (n2426 & n3328) | (n3305 & n3328);
  assign n3330 = n2419 | n2421;
  assign n3331 = (n2419 & n3307) | (n2419 & n3330) | (n3307 & n3330);
  assign n2460 = x31 & x42;
  assign n3335 = n2407 | n3314;
  assign n3783 = (n2348 & n3314) | (n2348 & n3335) | (n3314 & n3335);
  assign n3337 = n2460 & n3783;
  assign n49847 = n2460 & n11865;
  assign n66361 = n3742 & n49847;
  assign n49848 = (n3748 & n66361) | (n3748 & n49847) | (n66361 & n49847);
  assign n15552 = n2404 & n2460;
  assign n49849 = n11859 & n15552;
  assign n49845 = (n3720 & n49848) | (n3720 & n49849) | (n49848 & n49849);
  assign n15553 = (n2343 & n49845) | (n2343 & n15552) | (n49845 & n15552);
  assign n15556 = (n3720 & n49848) | (n3720 & n49849) | (n49848 & n49849);
  assign n11874 = (n3760 & n15553) | (n3760 & n15556) | (n15553 & n15556);
  assign n3785 = (n2407 & n2460) | (n2407 & n11874) | (n2460 & n11874);
  assign n3786 = (n3294 & n3337) | (n3294 & n3785) | (n3337 & n3785);
  assign n3787 = (n2350 & n3337) | (n2350 & n3785) | (n3337 & n3785);
  assign n3788 = (n3272 & n3786) | (n3272 & n3787) | (n3786 & n3787);
  assign n3340 = n2460 | n3783;
  assign n49853 = n2460 | n11865;
  assign n66362 = (n2460 & n3742) | (n2460 & n49853) | (n3742 & n49853);
  assign n49854 = (n3748 & n66362) | (n3748 & n49853) | (n66362 & n49853);
  assign n15558 = n2404 | n2460;
  assign n49855 = (n2460 & n11859) | (n2460 & n15558) | (n11859 & n15558);
  assign n49851 = (n3720 & n49854) | (n3720 & n49855) | (n49854 & n49855);
  assign n15559 = (n2343 & n49851) | (n2343 & n15558) | (n49851 & n15558);
  assign n15562 = (n3720 & n49854) | (n3720 & n49855) | (n49854 & n49855);
  assign n11877 = (n3760 & n15559) | (n3760 & n15562) | (n15559 & n15562);
  assign n3790 = n2407 | n11877;
  assign n3791 = (n3294 & n3340) | (n3294 & n3790) | (n3340 & n3790);
  assign n3792 = (n2350 & n3340) | (n2350 & n3790) | (n3340 & n3790);
  assign n3793 = (n3272 & n3791) | (n3272 & n3792) | (n3791 & n3792);
  assign n2463 = ~n3788 & n3793;
  assign n3795 = n2412 & n2463;
  assign n11878 = (n2414 & n2463) | (n2414 & n3795) | (n2463 & n3795);
  assign n3796 = (n3309 & n11878) | (n3309 & n3795) | (n11878 & n3795);
  assign n3798 = n2412 | n2463;
  assign n11879 = n2414 | n3798;
  assign n3799 = (n3309 & n11879) | (n3309 & n3798) | (n11879 & n3798);
  assign n2466 = ~n3796 & n3799;
  assign n2467 = x30 & x43;
  assign n2468 = n2466 & n2467;
  assign n2469 = n2466 | n2467;
  assign n2470 = ~n2468 & n2469;
  assign n2471 = n3331 & n2470;
  assign n2472 = n3331 | n2470;
  assign n2473 = ~n2471 & n2472;
  assign n2474 = x29 & x44;
  assign n2475 = n2473 & n2474;
  assign n2476 = n2473 | n2474;
  assign n2477 = ~n2475 & n2476;
  assign n2478 = n3329 & n2477;
  assign n2479 = n3329 | n2477;
  assign n2480 = ~n2478 & n2479;
  assign n2481 = x28 & x45;
  assign n2482 = n2480 & n2481;
  assign n2483 = n2480 | n2481;
  assign n2484 = ~n2482 & n2483;
  assign n2485 = n3327 & n2484;
  assign n2486 = n3327 | n2484;
  assign n2487 = ~n2485 & n2486;
  assign n2488 = x27 & x46;
  assign n2489 = n2487 & n2488;
  assign n2490 = n2487 | n2488;
  assign n2491 = ~n2489 & n2490;
  assign n2492 = n3325 & n2491;
  assign n2493 = n3325 | n2491;
  assign n2494 = ~n2492 & n2493;
  assign n2495 = x26 & x47;
  assign n2496 = n2494 & n2495;
  assign n2497 = n2494 | n2495;
  assign n2498 = ~n2496 & n2497;
  assign n2499 = n3323 & n2498;
  assign n2500 = n3323 | n2498;
  assign n2501 = ~n2499 & n2500;
  assign n3343 = n2496 | n2498;
  assign n3344 = (n2496 & n3323) | (n2496 & n3343) | (n3323 & n3343);
  assign n3345 = n2489 | n2491;
  assign n3346 = (n2489 & n3325) | (n2489 & n3345) | (n3325 & n3345);
  assign n3347 = n2482 | n2484;
  assign n3348 = (n2482 & n3327) | (n2482 & n3347) | (n3327 & n3347);
  assign n3349 = n2475 | n2477;
  assign n3350 = (n2475 & n3329) | (n2475 & n3349) | (n3329 & n3349);
  assign n2508 = x31 & x43;
  assign n3356 = n2508 & n3788;
  assign n3800 = n2508 & n3788;
  assign n3801 = (n2463 & n2508) | (n2463 & n3800) | (n2508 & n3800);
  assign n3803 = (n2412 & n3356) | (n2412 & n3801) | (n3356 & n3801);
  assign n11880 = n3356 | n3801;
  assign n11881 = (n2414 & n3803) | (n2414 & n11880) | (n3803 & n11880);
  assign n3804 = (n3309 & n11881) | (n3309 & n3803) | (n11881 & n3803);
  assign n3359 = n2508 | n3788;
  assign n3805 = n2508 | n3788;
  assign n3806 = n2463 | n3805;
  assign n3808 = (n2412 & n3359) | (n2412 & n3806) | (n3359 & n3806);
  assign n11882 = n3359 | n3806;
  assign n11883 = (n2414 & n3808) | (n2414 & n11882) | (n3808 & n11882);
  assign n3809 = (n3309 & n11883) | (n3309 & n3808) | (n11883 & n3808);
  assign n2511 = ~n3804 & n3809;
  assign n3811 = n2468 & n2511;
  assign n11884 = (n2470 & n2511) | (n2470 & n3811) | (n2511 & n3811);
  assign n3812 = (n3331 & n11884) | (n3331 & n3811) | (n11884 & n3811);
  assign n3814 = n2468 | n2511;
  assign n11885 = n2470 | n3814;
  assign n3815 = (n3331 & n11885) | (n3331 & n3814) | (n11885 & n3814);
  assign n2514 = ~n3812 & n3815;
  assign n2515 = x30 & x44;
  assign n2516 = n2514 & n2515;
  assign n2517 = n2514 | n2515;
  assign n2518 = ~n2516 & n2517;
  assign n2519 = n3350 & n2518;
  assign n2520 = n3350 | n2518;
  assign n2521 = ~n2519 & n2520;
  assign n2522 = x29 & x45;
  assign n2523 = n2521 & n2522;
  assign n2524 = n2521 | n2522;
  assign n2525 = ~n2523 & n2524;
  assign n2526 = n3348 & n2525;
  assign n2527 = n3348 | n2525;
  assign n2528 = ~n2526 & n2527;
  assign n2529 = x28 & x46;
  assign n2530 = n2528 & n2529;
  assign n2531 = n2528 | n2529;
  assign n2532 = ~n2530 & n2531;
  assign n2533 = n3346 & n2532;
  assign n2534 = n3346 | n2532;
  assign n2535 = ~n2533 & n2534;
  assign n2536 = x27 & x47;
  assign n2537 = n2535 & n2536;
  assign n2538 = n2535 | n2536;
  assign n2539 = ~n2537 & n2538;
  assign n2540 = n3344 & n2539;
  assign n2541 = n3344 | n2539;
  assign n2542 = ~n2540 & n2541;
  assign n3361 = n2537 | n2539;
  assign n3362 = (n2537 & n3344) | (n2537 & n3361) | (n3344 & n3361);
  assign n3363 = n2530 | n2532;
  assign n3364 = (n2530 & n3346) | (n2530 & n3363) | (n3346 & n3363);
  assign n3365 = n2523 | n2525;
  assign n3366 = (n2523 & n3348) | (n2523 & n3365) | (n3348 & n3365);
  assign n2548 = x31 & x44;
  assign n11886 = n2548 & n11881;
  assign n11887 = n2548 & n3803;
  assign n11888 = (n3309 & n11886) | (n3309 & n11887) | (n11886 & n11887);
  assign n3817 = (n2511 & n2548) | (n2511 & n11888) | (n2548 & n11888);
  assign n11889 = (n2468 & n3817) | (n2468 & n11888) | (n3817 & n11888);
  assign n15563 = n2548 | n11888;
  assign n15564 = (n2511 & n11888) | (n2511 & n15563) | (n11888 & n15563);
  assign n11891 = (n2470 & n11889) | (n2470 & n15564) | (n11889 & n15564);
  assign n3819 = (n2468 & n11888) | (n2468 & n3817) | (n11888 & n3817);
  assign n3820 = (n3331 & n11891) | (n3331 & n3819) | (n11891 & n3819);
  assign n11892 = n2548 | n11881;
  assign n11893 = n2548 | n3803;
  assign n11894 = (n3309 & n11892) | (n3309 & n11893) | (n11892 & n11893);
  assign n3822 = n2511 | n11894;
  assign n11895 = (n2468 & n3822) | (n2468 & n11894) | (n3822 & n11894);
  assign n15565 = n2511 | n11894;
  assign n11897 = (n2470 & n11895) | (n2470 & n15565) | (n11895 & n15565);
  assign n3824 = (n2468 & n11894) | (n2468 & n3822) | (n11894 & n3822);
  assign n3825 = (n3331 & n11897) | (n3331 & n3824) | (n11897 & n3824);
  assign n2551 = ~n3820 & n3825;
  assign n3827 = n2516 & n2551;
  assign n11898 = (n2518 & n2551) | (n2518 & n3827) | (n2551 & n3827);
  assign n3828 = (n3350 & n11898) | (n3350 & n3827) | (n11898 & n3827);
  assign n3830 = n2516 | n2551;
  assign n11899 = n2518 | n3830;
  assign n3831 = (n3350 & n11899) | (n3350 & n3830) | (n11899 & n3830);
  assign n2554 = ~n3828 & n3831;
  assign n2555 = x30 & x45;
  assign n2556 = n2554 & n2555;
  assign n2557 = n2554 | n2555;
  assign n2558 = ~n2556 & n2557;
  assign n2559 = n3366 & n2558;
  assign n2560 = n3366 | n2558;
  assign n2561 = ~n2559 & n2560;
  assign n2562 = x29 & x46;
  assign n2563 = n2561 & n2562;
  assign n2564 = n2561 | n2562;
  assign n2565 = ~n2563 & n2564;
  assign n2566 = n3364 & n2565;
  assign n2567 = n3364 | n2565;
  assign n2568 = ~n2566 & n2567;
  assign n2569 = x28 & x47;
  assign n2570 = n2568 & n2569;
  assign n2571 = n2568 | n2569;
  assign n2572 = ~n2570 & n2571;
  assign n2573 = n3362 & n2572;
  assign n2574 = n3362 | n2572;
  assign n2575 = ~n2573 & n2574;
  assign n3377 = n2570 | n2572;
  assign n3378 = (n2570 & n3362) | (n2570 & n3377) | (n3362 & n3377);
  assign n3379 = n2563 | n2565;
  assign n3380 = (n2563 & n3364) | (n2563 & n3379) | (n3364 & n3379);
  assign n2580 = x31 & x45;
  assign n11900 = n2580 & n11891;
  assign n11901 = n2580 & n3819;
  assign n11902 = (n3331 & n11900) | (n3331 & n11901) | (n11900 & n11901);
  assign n3833 = (n2551 & n2580) | (n2551 & n11902) | (n2580 & n11902);
  assign n11903 = (n2516 & n3833) | (n2516 & n11902) | (n3833 & n11902);
  assign n15566 = n2580 | n11902;
  assign n15567 = (n2551 & n11902) | (n2551 & n15566) | (n11902 & n15566);
  assign n11905 = (n2518 & n11903) | (n2518 & n15567) | (n11903 & n15567);
  assign n3835 = (n2516 & n11902) | (n2516 & n3833) | (n11902 & n3833);
  assign n3836 = (n3350 & n11905) | (n3350 & n3835) | (n11905 & n3835);
  assign n11906 = n2580 | n11891;
  assign n11907 = n2580 | n3819;
  assign n11908 = (n3331 & n11906) | (n3331 & n11907) | (n11906 & n11907);
  assign n3838 = n2551 | n11908;
  assign n11909 = (n2516 & n3838) | (n2516 & n11908) | (n3838 & n11908);
  assign n15568 = n2551 | n11908;
  assign n11911 = (n2518 & n11909) | (n2518 & n15568) | (n11909 & n15568);
  assign n3840 = (n2516 & n11908) | (n2516 & n3838) | (n11908 & n3838);
  assign n3841 = (n3350 & n11911) | (n3350 & n3840) | (n11911 & n3840);
  assign n2583 = ~n3836 & n3841;
  assign n3843 = n2556 & n2583;
  assign n11912 = (n2558 & n2583) | (n2558 & n3843) | (n2583 & n3843);
  assign n3844 = (n3366 & n11912) | (n3366 & n3843) | (n11912 & n3843);
  assign n3846 = n2556 | n2583;
  assign n11913 = n2558 | n3846;
  assign n3847 = (n3366 & n11913) | (n3366 & n3846) | (n11913 & n3846);
  assign n2586 = ~n3844 & n3847;
  assign n2587 = x30 & x46;
  assign n2588 = n2586 & n2587;
  assign n2589 = n2586 | n2587;
  assign n2590 = ~n2588 & n2589;
  assign n2591 = n3380 & n2590;
  assign n2592 = n3380 | n2590;
  assign n2593 = ~n2591 & n2592;
  assign n2594 = x29 & x47;
  assign n2595 = n2593 & n2594;
  assign n2596 = n2593 | n2594;
  assign n2597 = ~n2595 & n2596;
  assign n2598 = n3378 & n2597;
  assign n2599 = n3378 | n2597;
  assign n2600 = ~n2598 & n2599;
  assign n3391 = n2595 | n2597;
  assign n3392 = (n2595 & n3378) | (n2595 & n3391) | (n3378 & n3391);
  assign n2604 = x31 & x46;
  assign n11914 = n2604 & n11905;
  assign n11915 = n2604 & n3835;
  assign n11916 = (n3350 & n11914) | (n3350 & n11915) | (n11914 & n11915);
  assign n3849 = (n2583 & n2604) | (n2583 & n11916) | (n2604 & n11916);
  assign n11917 = (n2556 & n3849) | (n2556 & n11916) | (n3849 & n11916);
  assign n15569 = n2604 | n11916;
  assign n15570 = (n2583 & n11916) | (n2583 & n15569) | (n11916 & n15569);
  assign n11919 = (n2558 & n11917) | (n2558 & n15570) | (n11917 & n15570);
  assign n3851 = (n2556 & n11916) | (n2556 & n3849) | (n11916 & n3849);
  assign n3852 = (n3366 & n11919) | (n3366 & n3851) | (n11919 & n3851);
  assign n11920 = n2604 | n11905;
  assign n11921 = n2604 | n3835;
  assign n11922 = (n3350 & n11920) | (n3350 & n11921) | (n11920 & n11921);
  assign n3854 = n2583 | n11922;
  assign n11923 = (n2556 & n3854) | (n2556 & n11922) | (n3854 & n11922);
  assign n15571 = n2583 | n11922;
  assign n11925 = (n2558 & n11923) | (n2558 & n15571) | (n11923 & n15571);
  assign n3856 = (n2556 & n11922) | (n2556 & n3854) | (n11922 & n3854);
  assign n3857 = (n3366 & n11925) | (n3366 & n3856) | (n11925 & n3856);
  assign n2607 = ~n3852 & n3857;
  assign n3859 = n2588 & n2607;
  assign n11926 = (n2590 & n2607) | (n2590 & n3859) | (n2607 & n3859);
  assign n3860 = (n3380 & n11926) | (n3380 & n3859) | (n11926 & n3859);
  assign n3862 = n2588 | n2607;
  assign n11927 = n2590 | n3862;
  assign n3863 = (n3380 & n11927) | (n3380 & n3862) | (n11927 & n3862);
  assign n2610 = ~n3860 & n3863;
  assign n2611 = x30 & x47;
  assign n2612 = n2610 & n2611;
  assign n2613 = n2610 | n2611;
  assign n2614 = ~n2612 & n2613;
  assign n2615 = n3392 & n2614;
  assign n2616 = n3392 | n2614;
  assign n2617 = ~n2615 & n2616;
  assign n2620 = x31 & x47;
  assign n11928 = n2620 & n11919;
  assign n11929 = n2620 & n3851;
  assign n11930 = (n3366 & n11928) | (n3366 & n11929) | (n11928 & n11929);
  assign n3865 = (n2607 & n2620) | (n2607 & n11930) | (n2620 & n11930);
  assign n11931 = (n2588 & n3865) | (n2588 & n11930) | (n3865 & n11930);
  assign n15572 = n2620 | n11930;
  assign n15573 = (n2607 & n11930) | (n2607 & n15572) | (n11930 & n15572);
  assign n11933 = (n2590 & n11931) | (n2590 & n15573) | (n11931 & n15573);
  assign n3867 = (n2588 & n11930) | (n2588 & n3865) | (n11930 & n3865);
  assign n3868 = (n3380 & n11933) | (n3380 & n3867) | (n11933 & n3867);
  assign n11934 = n2620 | n11919;
  assign n11935 = n2620 | n3851;
  assign n11936 = (n3366 & n11934) | (n3366 & n11935) | (n11934 & n11935);
  assign n3870 = n2607 | n11936;
  assign n11937 = (n2588 & n3870) | (n2588 & n11936) | (n3870 & n11936);
  assign n15574 = n2607 | n11936;
  assign n11939 = (n2590 & n11937) | (n2590 & n15574) | (n11937 & n15574);
  assign n3872 = (n2588 & n11936) | (n2588 & n3870) | (n11936 & n3870);
  assign n3873 = (n3380 & n11939) | (n3380 & n3872) | (n11939 & n3872);
  assign n2623 = ~n3868 & n3873;
  assign n3875 = n2612 & n2623;
  assign n11940 = (n2614 & n2623) | (n2614 & n3875) | (n2623 & n3875);
  assign n3876 = (n3392 & n11940) | (n3392 & n3875) | (n11940 & n3875);
  assign n3878 = n2612 | n2623;
  assign n11941 = n2614 | n3878;
  assign n3879 = (n3392 & n11941) | (n3392 & n3878) | (n11941 & n3878);
  assign n2626 = ~n3876 & n3879;
  assign n3413 = n2623 | n3868;
  assign n3881 = (n2612 & n3413) | (n2612 & n3868) | (n3413 & n3868);
  assign n15575 = n2623 | n3868;
  assign n11943 = (n2614 & n3881) | (n2614 & n15575) | (n3881 & n15575);
  assign n3882 = (n3392 & n11943) | (n3392 & n3881) | (n11943 & n3881);
  assign n3947 = x48 & x80;
  assign n3948 = x49 & x80;
  assign n3949 = x48 & x81;
  assign n3950 = n3948 & n3949;
  assign n3951 = n3948 | n3949;
  assign n3952 = ~n3950 & n3951;
  assign n3953 = x50 & x80;
  assign n3954 = x49 & x81;
  assign n3955 = n3953 & n3954;
  assign n3956 = n3953 | n3954;
  assign n3957 = ~n3955 & n3956;
  assign n3958 = n3950 & n3957;
  assign n3959 = n3950 | n3957;
  assign n3960 = ~n3958 & n3959;
  assign n3961 = x48 & x82;
  assign n3962 = n3960 & n3961;
  assign n3963 = n3960 | n3961;
  assign n3964 = ~n3962 & n3963;
  assign n11944 = n3950 | n3955;
  assign n11945 = (n3955 & n3957) | (n3955 & n11944) | (n3957 & n11944);
  assign n3966 = x51 & x80;
  assign n3967 = x50 & x81;
  assign n3968 = n3966 & n3967;
  assign n3969 = n3966 | n3967;
  assign n3970 = ~n3968 & n3969;
  assign n3971 = n11945 & n3970;
  assign n3972 = n11945 | n3970;
  assign n3973 = ~n3971 & n3972;
  assign n3974 = x49 & x82;
  assign n3975 = n3973 & n3974;
  assign n3976 = n3973 | n3974;
  assign n3977 = ~n3975 & n3976;
  assign n3978 = n3962 & n3977;
  assign n3979 = n3962 | n3977;
  assign n3980 = ~n3978 & n3979;
  assign n3981 = x48 & x83;
  assign n3982 = n3980 & n3981;
  assign n3983 = n3980 | n3981;
  assign n3984 = ~n3982 & n3983;
  assign n11946 = n3962 | n3975;
  assign n11947 = (n3975 & n3977) | (n3975 & n11946) | (n3977 & n11946);
  assign n11948 = n3968 | n3970;
  assign n11949 = (n3968 & n11945) | (n3968 & n11948) | (n11945 & n11948);
  assign n3987 = x52 & x80;
  assign n3988 = x51 & x81;
  assign n3989 = n3987 & n3988;
  assign n3990 = n3987 | n3988;
  assign n3991 = ~n3989 & n3990;
  assign n3992 = n11949 & n3991;
  assign n3993 = n11949 | n3991;
  assign n3994 = ~n3992 & n3993;
  assign n3995 = x50 & x82;
  assign n3996 = n3994 & n3995;
  assign n3997 = n3994 | n3995;
  assign n3998 = ~n3996 & n3997;
  assign n3999 = n11947 & n3998;
  assign n4000 = n11947 | n3998;
  assign n4001 = ~n3999 & n4000;
  assign n4002 = x49 & x83;
  assign n4003 = n4001 & n4002;
  assign n4004 = n4001 | n4002;
  assign n4005 = ~n4003 & n4004;
  assign n4006 = n3982 & n4005;
  assign n4007 = n3982 | n4005;
  assign n4008 = ~n4006 & n4007;
  assign n4009 = x48 & x84;
  assign n4010 = n4008 & n4009;
  assign n4011 = n4008 | n4009;
  assign n4012 = ~n4010 & n4011;
  assign n11950 = n3982 | n4003;
  assign n11951 = (n4003 & n4005) | (n4003 & n11950) | (n4005 & n11950);
  assign n4016 = x53 & x80;
  assign n4017 = x52 & x81;
  assign n4018 = n4016 & n4017;
  assign n4019 = n4016 | n4017;
  assign n4020 = ~n4018 & n4019;
  assign n11952 = n3989 | n3991;
  assign n11954 = n4020 & n11952;
  assign n11955 = n3989 & n4020;
  assign n11956 = (n11949 & n11954) | (n11949 & n11955) | (n11954 & n11955);
  assign n11957 = n4020 | n11952;
  assign n11958 = n3989 | n4020;
  assign n11959 = (n11949 & n11957) | (n11949 & n11958) | (n11957 & n11958);
  assign n4023 = ~n11956 & n11959;
  assign n4024 = x51 & x82;
  assign n4025 = n4023 & n4024;
  assign n4026 = n4023 | n4024;
  assign n4027 = ~n4025 & n4026;
  assign n11960 = n3996 & n4027;
  assign n11961 = (n3999 & n4027) | (n3999 & n11960) | (n4027 & n11960);
  assign n11962 = n3996 | n4027;
  assign n11963 = n3999 | n11962;
  assign n4030 = ~n11961 & n11963;
  assign n4031 = x50 & x83;
  assign n4032 = n4030 & n4031;
  assign n4033 = n4030 | n4031;
  assign n4034 = ~n4032 & n4033;
  assign n4035 = n11951 & n4034;
  assign n4036 = n11951 | n4034;
  assign n4037 = ~n4035 & n4036;
  assign n4038 = x49 & x84;
  assign n4039 = n4037 & n4038;
  assign n4040 = n4037 | n4038;
  assign n4041 = ~n4039 & n4040;
  assign n4042 = n4010 & n4041;
  assign n4043 = n4010 | n4041;
  assign n4044 = ~n4042 & n4043;
  assign n4045 = x48 & x85;
  assign n4046 = n4044 & n4045;
  assign n4047 = n4044 | n4045;
  assign n4048 = ~n4046 & n4047;
  assign n11964 = n4010 | n4039;
  assign n11965 = (n4039 & n4041) | (n4039 & n11964) | (n4041 & n11964);
  assign n4050 = n4032 | n4035;
  assign n4053 = x54 & x80;
  assign n4054 = x53 & x81;
  assign n4055 = n4053 & n4054;
  assign n4056 = n4053 | n4054;
  assign n4057 = ~n4055 & n4056;
  assign n11966 = n4018 & n4057;
  assign n11967 = (n4057 & n11956) | (n4057 & n11966) | (n11956 & n11966);
  assign n11968 = n4018 | n4057;
  assign n11969 = n11956 | n11968;
  assign n4060 = ~n11967 & n11969;
  assign n4061 = x52 & x82;
  assign n4062 = n4060 & n4061;
  assign n4063 = n4060 | n4061;
  assign n4064 = ~n4062 & n4063;
  assign n11970 = n4025 & n4064;
  assign n11971 = (n4064 & n11961) | (n4064 & n11970) | (n11961 & n11970);
  assign n11972 = n4025 | n4064;
  assign n11973 = n11961 | n11972;
  assign n4067 = ~n11971 & n11973;
  assign n4068 = x51 & x83;
  assign n4069 = n4067 & n4068;
  assign n4070 = n4067 | n4068;
  assign n4071 = ~n4069 & n4070;
  assign n4072 = n4050 & n4071;
  assign n4073 = n4050 | n4071;
  assign n4074 = ~n4072 & n4073;
  assign n4075 = x50 & x84;
  assign n4076 = n4074 & n4075;
  assign n4077 = n4074 | n4075;
  assign n4078 = ~n4076 & n4077;
  assign n4079 = n11965 & n4078;
  assign n4080 = n11965 | n4078;
  assign n4081 = ~n4079 & n4080;
  assign n4082 = x49 & x85;
  assign n4083 = n4081 & n4082;
  assign n4084 = n4081 | n4082;
  assign n4085 = ~n4083 & n4084;
  assign n4086 = n4046 & n4085;
  assign n4087 = n4046 | n4085;
  assign n4088 = ~n4086 & n4087;
  assign n4089 = x48 & x86;
  assign n4090 = n4088 & n4089;
  assign n4091 = n4088 | n4089;
  assign n4092 = ~n4090 & n4091;
  assign n49856 = n4045 | n4082;
  assign n49857 = (n4044 & n4082) | (n4044 & n49856) | (n4082 & n49856);
  assign n15577 = (n4046 & n4081) | (n4046 & n49857) | (n4081 & n49857);
  assign n11975 = (n4083 & n4085) | (n4083 & n15577) | (n4085 & n15577);
  assign n11976 = n4076 | n11965;
  assign n11977 = (n4076 & n4078) | (n4076 & n11976) | (n4078 & n11976);
  assign n11978 = n4069 | n4071;
  assign n11979 = (n4050 & n4069) | (n4050 & n11978) | (n4069 & n11978);
  assign n4098 = x55 & x80;
  assign n4099 = x54 & x81;
  assign n4100 = n4098 & n4099;
  assign n4101 = n4098 | n4099;
  assign n4102 = ~n4100 & n4101;
  assign n15578 = n4018 | n4055;
  assign n15579 = (n4055 & n4057) | (n4055 & n15578) | (n4057 & n15578);
  assign n11983 = n4102 & n15579;
  assign n11981 = n4055 | n4057;
  assign n11984 = n4102 & n11981;
  assign n11985 = (n11956 & n11983) | (n11956 & n11984) | (n11983 & n11984);
  assign n11986 = n4102 | n15579;
  assign n11987 = n4102 | n11981;
  assign n11988 = (n11956 & n11986) | (n11956 & n11987) | (n11986 & n11987);
  assign n4105 = ~n11985 & n11988;
  assign n4106 = x53 & x82;
  assign n4107 = n4105 & n4106;
  assign n4108 = n4105 | n4106;
  assign n4109 = ~n4107 & n4108;
  assign n11989 = n4062 & n4109;
  assign n11990 = (n4109 & n11971) | (n4109 & n11989) | (n11971 & n11989);
  assign n11991 = n4062 | n4109;
  assign n11992 = n11971 | n11991;
  assign n4112 = ~n11990 & n11992;
  assign n4113 = x52 & x83;
  assign n4114 = n4112 & n4113;
  assign n4115 = n4112 | n4113;
  assign n4116 = ~n4114 & n4115;
  assign n4117 = n11979 & n4116;
  assign n4118 = n11979 | n4116;
  assign n4119 = ~n4117 & n4118;
  assign n4120 = x51 & x84;
  assign n4121 = n4119 & n4120;
  assign n4122 = n4119 | n4120;
  assign n4123 = ~n4121 & n4122;
  assign n4124 = n11977 & n4123;
  assign n4125 = n11977 | n4123;
  assign n4126 = ~n4124 & n4125;
  assign n4127 = x50 & x85;
  assign n4128 = n4126 & n4127;
  assign n4129 = n4126 | n4127;
  assign n4130 = ~n4128 & n4129;
  assign n4131 = n11975 & n4130;
  assign n4132 = n11975 | n4130;
  assign n4133 = ~n4131 & n4132;
  assign n4134 = x49 & x86;
  assign n4135 = n4133 & n4134;
  assign n4136 = n4133 | n4134;
  assign n4137 = ~n4135 & n4136;
  assign n4138 = n4090 & n4137;
  assign n4139 = n4090 | n4137;
  assign n4140 = ~n4138 & n4139;
  assign n4141 = x48 & x87;
  assign n4142 = n4140 & n4141;
  assign n4143 = n4140 | n4141;
  assign n4144 = ~n4142 & n4143;
  assign n11993 = n4090 | n4135;
  assign n11994 = (n4135 & n4137) | (n4135 & n11993) | (n4137 & n11993);
  assign n4146 = n4128 | n4131;
  assign n4147 = n4121 | n4124;
  assign n11995 = n4114 | n4116;
  assign n11996 = (n4114 & n11979) | (n4114 & n11995) | (n11979 & n11995);
  assign n4151 = x56 & x80;
  assign n4152 = x55 & x81;
  assign n4153 = n4151 & n4152;
  assign n4154 = n4151 | n4152;
  assign n4155 = ~n4153 & n4154;
  assign n12000 = n4100 & n4155;
  assign n15582 = (n4155 & n11984) | (n4155 & n12000) | (n11984 & n12000);
  assign n15583 = (n4155 & n11983) | (n4155 & n12000) | (n11983 & n12000);
  assign n15584 = (n11956 & n15582) | (n11956 & n15583) | (n15582 & n15583);
  assign n12002 = n4100 | n4155;
  assign n15585 = n11984 | n12002;
  assign n15586 = n11983 | n12002;
  assign n15587 = (n11956 & n15585) | (n11956 & n15586) | (n15585 & n15586);
  assign n4158 = ~n15584 & n15587;
  assign n4159 = x54 & x82;
  assign n4160 = n4158 & n4159;
  assign n4161 = n4158 | n4159;
  assign n4162 = ~n4160 & n4161;
  assign n11998 = n4107 | n4109;
  assign n15588 = n4162 & n11998;
  assign n15580 = n4062 | n4107;
  assign n15581 = (n4107 & n4109) | (n4107 & n15580) | (n4109 & n15580);
  assign n15589 = n4162 & n15581;
  assign n15590 = (n11971 & n15588) | (n11971 & n15589) | (n15588 & n15589);
  assign n15591 = n4162 | n11998;
  assign n15592 = n4162 | n15581;
  assign n15593 = (n11971 & n15591) | (n11971 & n15592) | (n15591 & n15592);
  assign n4165 = ~n15590 & n15593;
  assign n4166 = x53 & x83;
  assign n4167 = n4165 & n4166;
  assign n4168 = n4165 | n4166;
  assign n4169 = ~n4167 & n4168;
  assign n4170 = n11996 & n4169;
  assign n4171 = n11996 | n4169;
  assign n4172 = ~n4170 & n4171;
  assign n4173 = x52 & x84;
  assign n4174 = n4172 & n4173;
  assign n4175 = n4172 | n4173;
  assign n4176 = ~n4174 & n4175;
  assign n4177 = n4147 & n4176;
  assign n4178 = n4147 | n4176;
  assign n4179 = ~n4177 & n4178;
  assign n4180 = x51 & x85;
  assign n4181 = n4179 & n4180;
  assign n4182 = n4179 | n4180;
  assign n4183 = ~n4181 & n4182;
  assign n4184 = n4146 & n4183;
  assign n4185 = n4146 | n4183;
  assign n4186 = ~n4184 & n4185;
  assign n4187 = x50 & x86;
  assign n4188 = n4186 & n4187;
  assign n4189 = n4186 | n4187;
  assign n4190 = ~n4188 & n4189;
  assign n4191 = n11994 & n4190;
  assign n4192 = n11994 | n4190;
  assign n4193 = ~n4191 & n4192;
  assign n4194 = x49 & x87;
  assign n4195 = n4193 & n4194;
  assign n4196 = n4193 | n4194;
  assign n4197 = ~n4195 & n4196;
  assign n4198 = n4142 & n4197;
  assign n4199 = n4142 | n4197;
  assign n4200 = ~n4198 & n4199;
  assign n4201 = x48 & x88;
  assign n4202 = n4200 & n4201;
  assign n4203 = n4200 | n4201;
  assign n4204 = ~n4202 & n4203;
  assign n49858 = n4141 | n4194;
  assign n49859 = (n4140 & n4194) | (n4140 & n49858) | (n4194 & n49858);
  assign n15595 = (n4142 & n4193) | (n4142 & n49859) | (n4193 & n49859);
  assign n12005 = (n4195 & n4197) | (n4195 & n15595) | (n4197 & n15595);
  assign n12006 = n4188 | n11994;
  assign n12007 = (n4188 & n4190) | (n4188 & n12006) | (n4190 & n12006);
  assign n4207 = n4181 | n4184;
  assign n12008 = n4174 | n4176;
  assign n12009 = (n4147 & n4174) | (n4147 & n12008) | (n4174 & n12008);
  assign n11999 = (n11971 & n15581) | (n11971 & n11998) | (n15581 & n11998);
  assign n4212 = x57 & x80;
  assign n4213 = x56 & x81;
  assign n4214 = n4212 & n4213;
  assign n4215 = n4212 | n4213;
  assign n4216 = ~n4214 & n4215;
  assign n15596 = n4100 | n4153;
  assign n15597 = (n4153 & n4155) | (n4153 & n15596) | (n4155 & n15596);
  assign n12017 = n4216 & n15597;
  assign n12015 = n4153 | n4155;
  assign n12018 = n4216 & n12015;
  assign n15598 = (n11984 & n12017) | (n11984 & n12018) | (n12017 & n12018);
  assign n15599 = (n11983 & n12017) | (n11983 & n12018) | (n12017 & n12018);
  assign n15600 = (n11956 & n15598) | (n11956 & n15599) | (n15598 & n15599);
  assign n12020 = n4216 | n15597;
  assign n12021 = n4216 | n12015;
  assign n15601 = (n11984 & n12020) | (n11984 & n12021) | (n12020 & n12021);
  assign n15602 = (n11983 & n12020) | (n11983 & n12021) | (n12020 & n12021);
  assign n15603 = (n11956 & n15601) | (n11956 & n15602) | (n15601 & n15602);
  assign n4219 = ~n15600 & n15603;
  assign n4220 = x55 & x82;
  assign n4221 = n4219 & n4220;
  assign n4222 = n4219 | n4220;
  assign n4223 = ~n4221 & n4222;
  assign n12012 = n4160 | n4162;
  assign n12023 = n4223 & n12012;
  assign n12024 = n4160 & n4223;
  assign n12025 = (n11999 & n12023) | (n11999 & n12024) | (n12023 & n12024);
  assign n12026 = n4223 | n12012;
  assign n12027 = n4160 | n4223;
  assign n12028 = (n11999 & n12026) | (n11999 & n12027) | (n12026 & n12027);
  assign n4226 = ~n12025 & n12028;
  assign n4227 = x54 & x83;
  assign n4228 = n4226 & n4227;
  assign n4229 = n4226 | n4227;
  assign n4230 = ~n4228 & n4229;
  assign n12010 = n4167 | n4169;
  assign n15604 = n4230 & n12010;
  assign n15605 = n4167 & n4230;
  assign n15606 = (n11996 & n15604) | (n11996 & n15605) | (n15604 & n15605);
  assign n15607 = n4230 | n12010;
  assign n15608 = n4167 | n4230;
  assign n15609 = (n11996 & n15607) | (n11996 & n15608) | (n15607 & n15608);
  assign n4233 = ~n15606 & n15609;
  assign n4234 = x53 & x84;
  assign n4235 = n4233 & n4234;
  assign n4236 = n4233 | n4234;
  assign n4237 = ~n4235 & n4236;
  assign n4238 = n12009 & n4237;
  assign n4239 = n12009 | n4237;
  assign n4240 = ~n4238 & n4239;
  assign n4241 = x52 & x85;
  assign n4242 = n4240 & n4241;
  assign n4243 = n4240 | n4241;
  assign n4244 = ~n4242 & n4243;
  assign n4245 = n4207 & n4244;
  assign n4246 = n4207 | n4244;
  assign n4247 = ~n4245 & n4246;
  assign n4248 = x51 & x86;
  assign n4249 = n4247 & n4248;
  assign n4250 = n4247 | n4248;
  assign n4251 = ~n4249 & n4250;
  assign n4252 = n12007 & n4251;
  assign n4253 = n12007 | n4251;
  assign n4254 = ~n4252 & n4253;
  assign n4255 = x50 & x87;
  assign n4256 = n4254 & n4255;
  assign n4257 = n4254 | n4255;
  assign n4258 = ~n4256 & n4257;
  assign n4259 = n12005 & n4258;
  assign n4260 = n12005 | n4258;
  assign n4261 = ~n4259 & n4260;
  assign n4262 = x49 & x88;
  assign n4263 = n4261 & n4262;
  assign n4264 = n4261 | n4262;
  assign n4265 = ~n4263 & n4264;
  assign n4266 = n4202 & n4265;
  assign n4267 = n4202 | n4265;
  assign n4268 = ~n4266 & n4267;
  assign n4269 = x48 & x89;
  assign n4270 = n4268 & n4269;
  assign n4271 = n4268 | n4269;
  assign n4272 = ~n4270 & n4271;
  assign n49860 = n4201 | n4262;
  assign n49861 = (n4200 & n4262) | (n4200 & n49860) | (n4262 & n49860);
  assign n15611 = (n4202 & n4261) | (n4202 & n49861) | (n4261 & n49861);
  assign n12030 = (n4263 & n4265) | (n4263 & n15611) | (n4265 & n15611);
  assign n12031 = n4256 | n12005;
  assign n12032 = (n4256 & n4258) | (n4256 & n12031) | (n4258 & n12031);
  assign n12033 = n4249 | n12007;
  assign n12034 = (n4249 & n4251) | (n4249 & n12033) | (n4251 & n12033);
  assign n12035 = n4242 | n4244;
  assign n12036 = (n4207 & n4242) | (n4207 & n12035) | (n4242 & n12035);
  assign n12011 = (n4167 & n11996) | (n4167 & n12010) | (n11996 & n12010);
  assign n15612 = n4214 | n4216;
  assign n15613 = (n4214 & n15597) | (n4214 & n15612) | (n15597 & n15612);
  assign n15614 = (n4214 & n12015) | (n4214 & n15612) | (n12015 & n15612);
  assign n15615 = (n11984 & n15613) | (n11984 & n15614) | (n15613 & n15614);
  assign n15616 = (n11983 & n15613) | (n11983 & n15614) | (n15613 & n15614);
  assign n15617 = (n11956 & n15615) | (n11956 & n15616) | (n15615 & n15616);
  assign n4281 = x58 & x80;
  assign n4282 = x57 & x81;
  assign n4283 = n4281 & n4282;
  assign n4284 = n4281 | n4282;
  assign n4285 = ~n4283 & n4284;
  assign n4286 = n15617 & n4285;
  assign n4287 = n15617 | n4285;
  assign n4288 = ~n4286 & n4287;
  assign n4289 = x56 & x82;
  assign n4290 = n4288 & n4289;
  assign n4291 = n4288 | n4289;
  assign n4292 = ~n4290 & n4291;
  assign n12044 = n4221 & n4292;
  assign n15618 = (n4292 & n12023) | (n4292 & n12044) | (n12023 & n12044);
  assign n15619 = (n4292 & n12024) | (n4292 & n12044) | (n12024 & n12044);
  assign n15620 = (n11999 & n15618) | (n11999 & n15619) | (n15618 & n15619);
  assign n12046 = n4221 | n4292;
  assign n15621 = n12023 | n12046;
  assign n15622 = n12024 | n12046;
  assign n15623 = (n11999 & n15621) | (n11999 & n15622) | (n15621 & n15622);
  assign n4295 = ~n15620 & n15623;
  assign n4296 = x55 & x83;
  assign n4297 = n4295 & n4296;
  assign n4298 = n4295 | n4296;
  assign n4299 = ~n4297 & n4298;
  assign n12039 = n4228 | n4230;
  assign n12048 = n4299 & n12039;
  assign n12049 = n4228 & n4299;
  assign n12050 = (n12011 & n12048) | (n12011 & n12049) | (n12048 & n12049);
  assign n12051 = n4299 | n12039;
  assign n12052 = n4228 | n4299;
  assign n12053 = (n12011 & n12051) | (n12011 & n12052) | (n12051 & n12052);
  assign n4302 = ~n12050 & n12053;
  assign n4303 = x54 & x84;
  assign n4304 = n4302 & n4303;
  assign n4305 = n4302 | n4303;
  assign n4306 = ~n4304 & n4305;
  assign n12037 = n4235 | n4237;
  assign n15624 = n4306 & n12037;
  assign n15625 = n4235 & n4306;
  assign n15626 = (n12009 & n15624) | (n12009 & n15625) | (n15624 & n15625);
  assign n15627 = n4306 | n12037;
  assign n15628 = n4235 | n4306;
  assign n15629 = (n12009 & n15627) | (n12009 & n15628) | (n15627 & n15628);
  assign n4309 = ~n15626 & n15629;
  assign n4310 = x53 & x85;
  assign n4311 = n4309 & n4310;
  assign n4312 = n4309 | n4310;
  assign n4313 = ~n4311 & n4312;
  assign n4314 = n12036 & n4313;
  assign n4315 = n12036 | n4313;
  assign n4316 = ~n4314 & n4315;
  assign n4317 = x52 & x86;
  assign n4318 = n4316 & n4317;
  assign n4319 = n4316 | n4317;
  assign n4320 = ~n4318 & n4319;
  assign n4321 = n12034 & n4320;
  assign n4322 = n12034 | n4320;
  assign n4323 = ~n4321 & n4322;
  assign n4324 = x51 & x87;
  assign n4325 = n4323 & n4324;
  assign n4326 = n4323 | n4324;
  assign n4327 = ~n4325 & n4326;
  assign n4328 = n12032 & n4327;
  assign n4329 = n12032 | n4327;
  assign n4330 = ~n4328 & n4329;
  assign n4331 = x50 & x88;
  assign n4332 = n4330 & n4331;
  assign n4333 = n4330 | n4331;
  assign n4334 = ~n4332 & n4333;
  assign n4335 = n12030 & n4334;
  assign n4336 = n12030 | n4334;
  assign n4337 = ~n4335 & n4336;
  assign n4338 = x49 & x89;
  assign n4339 = n4337 & n4338;
  assign n4340 = n4337 | n4338;
  assign n4341 = ~n4339 & n4340;
  assign n4342 = n4270 & n4341;
  assign n4343 = n4270 | n4341;
  assign n4344 = ~n4342 & n4343;
  assign n4345 = x48 & x90;
  assign n4346 = n4344 & n4345;
  assign n4347 = n4344 | n4345;
  assign n4348 = ~n4346 & n4347;
  assign n12054 = n4270 | n4339;
  assign n12055 = (n4339 & n4341) | (n4339 & n12054) | (n4341 & n12054);
  assign n4350 = n4332 | n4335;
  assign n4351 = n4325 | n4328;
  assign n12038 = (n4235 & n12009) | (n4235 & n12037) | (n12009 & n12037);
  assign n12061 = n4290 | n4292;
  assign n15630 = n4221 | n4290;
  assign n15631 = (n4290 & n4292) | (n4290 & n15630) | (n4292 & n15630);
  assign n15632 = (n12023 & n12061) | (n12023 & n15631) | (n12061 & n15631);
  assign n15633 = (n12024 & n12061) | (n12024 & n15631) | (n12061 & n15631);
  assign n15634 = (n11999 & n15632) | (n11999 & n15633) | (n15632 & n15633);
  assign n4358 = x59 & x80;
  assign n4359 = x58 & x81;
  assign n4360 = n4358 & n4359;
  assign n4361 = n4358 | n4359;
  assign n4362 = ~n4360 & n4361;
  assign n12063 = n4283 | n4285;
  assign n12065 = n4362 & n12063;
  assign n12066 = n4283 & n4362;
  assign n12067 = (n15617 & n12065) | (n15617 & n12066) | (n12065 & n12066);
  assign n12068 = n4362 | n12063;
  assign n12069 = n4283 | n4362;
  assign n12070 = (n15617 & n12068) | (n15617 & n12069) | (n12068 & n12069);
  assign n4365 = ~n12067 & n12070;
  assign n4366 = x57 & x82;
  assign n4367 = n4365 & n4366;
  assign n4368 = n4365 | n4366;
  assign n4369 = ~n4367 & n4368;
  assign n4370 = n15634 & n4369;
  assign n4371 = n15634 | n4369;
  assign n4372 = ~n4370 & n4371;
  assign n4373 = x56 & x83;
  assign n4374 = n4372 & n4373;
  assign n4375 = n4372 | n4373;
  assign n4376 = ~n4374 & n4375;
  assign n12071 = n4297 & n4376;
  assign n12072 = (n4376 & n12050) | (n4376 & n12071) | (n12050 & n12071);
  assign n12073 = n4297 | n4376;
  assign n12074 = n12050 | n12073;
  assign n4379 = ~n12072 & n12074;
  assign n4380 = x55 & x84;
  assign n4381 = n4379 & n4380;
  assign n4382 = n4379 | n4380;
  assign n4383 = ~n4381 & n4382;
  assign n12058 = n4304 | n4306;
  assign n12075 = n4383 & n12058;
  assign n12076 = n4304 & n4383;
  assign n12077 = (n12038 & n12075) | (n12038 & n12076) | (n12075 & n12076);
  assign n12078 = n4383 | n12058;
  assign n12079 = n4304 | n4383;
  assign n12080 = (n12038 & n12078) | (n12038 & n12079) | (n12078 & n12079);
  assign n4386 = ~n12077 & n12080;
  assign n4387 = x54 & x85;
  assign n4388 = n4386 & n4387;
  assign n4389 = n4386 | n4387;
  assign n4390 = ~n4388 & n4389;
  assign n12056 = n4311 | n4313;
  assign n15635 = n4390 & n12056;
  assign n15636 = n4311 & n4390;
  assign n15637 = (n12036 & n15635) | (n12036 & n15636) | (n15635 & n15636);
  assign n15638 = n4390 | n12056;
  assign n15639 = n4311 | n4390;
  assign n15640 = (n12036 & n15638) | (n12036 & n15639) | (n15638 & n15639);
  assign n4393 = ~n15637 & n15640;
  assign n4394 = x53 & x86;
  assign n4395 = n4393 & n4394;
  assign n4396 = n4393 | n4394;
  assign n4397 = ~n4395 & n4396;
  assign n15641 = n4318 & n4397;
  assign n15642 = (n4321 & n4397) | (n4321 & n15641) | (n4397 & n15641);
  assign n15643 = n4318 | n4397;
  assign n15644 = n4321 | n15643;
  assign n4400 = ~n15642 & n15644;
  assign n4401 = x52 & x87;
  assign n4402 = n4400 & n4401;
  assign n4403 = n4400 | n4401;
  assign n4404 = ~n4402 & n4403;
  assign n4405 = n4351 & n4404;
  assign n4406 = n4351 | n4404;
  assign n4407 = ~n4405 & n4406;
  assign n4408 = x51 & x88;
  assign n4409 = n4407 & n4408;
  assign n4410 = n4407 | n4408;
  assign n4411 = ~n4409 & n4410;
  assign n4412 = n4350 & n4411;
  assign n4413 = n4350 | n4411;
  assign n4414 = ~n4412 & n4413;
  assign n4415 = x50 & x89;
  assign n4416 = n4414 & n4415;
  assign n4417 = n4414 | n4415;
  assign n4418 = ~n4416 & n4417;
  assign n4419 = n12055 & n4418;
  assign n4420 = n12055 | n4418;
  assign n4421 = ~n4419 & n4420;
  assign n4422 = x49 & x90;
  assign n4423 = n4421 & n4422;
  assign n4424 = n4421 | n4422;
  assign n4425 = ~n4423 & n4424;
  assign n4426 = n4346 & n4425;
  assign n4427 = n4346 | n4425;
  assign n4428 = ~n4426 & n4427;
  assign n4429 = x48 & x91;
  assign n4430 = n4428 & n4429;
  assign n4431 = n4428 | n4429;
  assign n4432 = ~n4430 & n4431;
  assign n49862 = n4345 | n4422;
  assign n49863 = (n4344 & n4422) | (n4344 & n49862) | (n4422 & n49862);
  assign n15646 = (n4346 & n4421) | (n4346 & n49863) | (n4421 & n49863);
  assign n12082 = (n4423 & n4425) | (n4423 & n15646) | (n4425 & n15646);
  assign n12083 = n4416 | n12055;
  assign n12084 = (n4416 & n4418) | (n4416 & n12083) | (n4418 & n12083);
  assign n4435 = n4409 | n4412;
  assign n15647 = n4402 | n4404;
  assign n15648 = (n4351 & n4402) | (n4351 & n15647) | (n4402 & n15647);
  assign n4352 = n4318 | n4321;
  assign n12057 = (n4311 & n12036) | (n4311 & n12056) | (n12036 & n12056);
  assign n4443 = x60 & x80;
  assign n4444 = x59 & x81;
  assign n4445 = n4443 & n4444;
  assign n4446 = n4443 | n4444;
  assign n4447 = ~n4445 & n4446;
  assign n15649 = n4360 | n4362;
  assign n15650 = (n4360 & n12063) | (n4360 & n15649) | (n12063 & n15649);
  assign n12094 = n4447 & n15650;
  assign n15651 = n4283 | n4360;
  assign n15652 = (n4360 & n4362) | (n4360 & n15651) | (n4362 & n15651);
  assign n12095 = n4447 & n15652;
  assign n12096 = (n15617 & n12094) | (n15617 & n12095) | (n12094 & n12095);
  assign n12097 = n4447 | n15650;
  assign n12098 = n4447 | n15652;
  assign n12099 = (n15617 & n12097) | (n15617 & n12098) | (n12097 & n12098);
  assign n4450 = ~n12096 & n12099;
  assign n4451 = x58 & x82;
  assign n4452 = n4450 & n4451;
  assign n4453 = n4450 | n4451;
  assign n4454 = ~n4452 & n4453;
  assign n12089 = n4367 | n4369;
  assign n12100 = n4454 & n12089;
  assign n12101 = n4367 & n4454;
  assign n12102 = (n15634 & n12100) | (n15634 & n12101) | (n12100 & n12101);
  assign n12103 = n4454 | n12089;
  assign n12104 = n4367 | n4454;
  assign n12105 = (n15634 & n12103) | (n15634 & n12104) | (n12103 & n12104);
  assign n4457 = ~n12102 & n12105;
  assign n4458 = x57 & x83;
  assign n4459 = n4457 & n4458;
  assign n4460 = n4457 | n4458;
  assign n4461 = ~n4459 & n4460;
  assign n12106 = n4374 & n4461;
  assign n15653 = (n4461 & n12071) | (n4461 & n12106) | (n12071 & n12106);
  assign n15654 = (n4376 & n4461) | (n4376 & n12106) | (n4461 & n12106);
  assign n15655 = (n12050 & n15653) | (n12050 & n15654) | (n15653 & n15654);
  assign n12108 = n4374 | n4461;
  assign n15656 = n12071 | n12108;
  assign n15657 = n4376 | n12108;
  assign n15658 = (n12050 & n15656) | (n12050 & n15657) | (n15656 & n15657);
  assign n4464 = ~n15655 & n15658;
  assign n4465 = x56 & x84;
  assign n4466 = n4464 & n4465;
  assign n4467 = n4464 | n4465;
  assign n4468 = ~n4466 & n4467;
  assign n12110 = n4381 & n4468;
  assign n12111 = (n4468 & n12077) | (n4468 & n12110) | (n12077 & n12110);
  assign n12112 = n4381 | n4468;
  assign n12113 = n12077 | n12112;
  assign n4471 = ~n12111 & n12113;
  assign n4472 = x55 & x85;
  assign n4473 = n4471 & n4472;
  assign n4474 = n4471 | n4472;
  assign n4475 = ~n4473 & n4474;
  assign n12087 = n4388 | n4390;
  assign n12114 = n4475 & n12087;
  assign n12115 = n4388 & n4475;
  assign n12116 = (n12057 & n12114) | (n12057 & n12115) | (n12114 & n12115);
  assign n12117 = n4475 | n12087;
  assign n12118 = n4388 | n4475;
  assign n12119 = (n12057 & n12117) | (n12057 & n12118) | (n12117 & n12118);
  assign n4478 = ~n12116 & n12119;
  assign n4479 = x54 & x86;
  assign n4480 = n4478 & n4479;
  assign n4481 = n4478 | n4479;
  assign n4482 = ~n4480 & n4481;
  assign n12085 = n4395 | n4397;
  assign n15659 = n4482 & n12085;
  assign n15660 = n4395 & n4482;
  assign n15661 = (n4352 & n15659) | (n4352 & n15660) | (n15659 & n15660);
  assign n15662 = n4482 | n12085;
  assign n15663 = n4395 | n4482;
  assign n15664 = (n4352 & n15662) | (n4352 & n15663) | (n15662 & n15663);
  assign n4485 = ~n15661 & n15664;
  assign n4486 = x53 & x87;
  assign n4487 = n4485 & n4486;
  assign n4488 = n4485 | n4486;
  assign n4489 = ~n4487 & n4488;
  assign n4490 = n15648 & n4489;
  assign n4491 = n15648 | n4489;
  assign n4492 = ~n4490 & n4491;
  assign n4493 = x52 & x88;
  assign n4494 = n4492 & n4493;
  assign n4495 = n4492 | n4493;
  assign n4496 = ~n4494 & n4495;
  assign n4497 = n4435 & n4496;
  assign n4498 = n4435 | n4496;
  assign n4499 = ~n4497 & n4498;
  assign n4500 = x51 & x89;
  assign n4501 = n4499 & n4500;
  assign n4502 = n4499 | n4500;
  assign n4503 = ~n4501 & n4502;
  assign n4504 = n12084 & n4503;
  assign n4505 = n12084 | n4503;
  assign n4506 = ~n4504 & n4505;
  assign n4507 = x50 & x90;
  assign n4508 = n4506 & n4507;
  assign n4509 = n4506 | n4507;
  assign n4510 = ~n4508 & n4509;
  assign n4511 = n12082 & n4510;
  assign n4512 = n12082 | n4510;
  assign n4513 = ~n4511 & n4512;
  assign n4514 = x49 & x91;
  assign n4515 = n4513 & n4514;
  assign n4516 = n4513 | n4514;
  assign n4517 = ~n4515 & n4516;
  assign n4518 = n4430 & n4517;
  assign n4519 = n4430 | n4517;
  assign n4520 = ~n4518 & n4519;
  assign n4521 = x48 & x92;
  assign n4522 = n4520 & n4521;
  assign n4523 = n4520 | n4521;
  assign n4524 = ~n4522 & n4523;
  assign n49864 = n4429 | n4514;
  assign n49865 = (n4428 & n4514) | (n4428 & n49864) | (n4514 & n49864);
  assign n15666 = (n4430 & n4513) | (n4430 & n49865) | (n4513 & n49865);
  assign n12121 = (n4515 & n4517) | (n4515 & n15666) | (n4517 & n15666);
  assign n12122 = n4508 | n12082;
  assign n12123 = (n4508 & n4510) | (n4508 & n12122) | (n4510 & n12122);
  assign n12124 = n4501 | n12084;
  assign n12125 = (n4501 & n4503) | (n4501 & n12124) | (n4503 & n12124);
  assign n15667 = n4494 | n4496;
  assign n15668 = (n4435 & n4494) | (n4435 & n15667) | (n4494 & n15667);
  assign n12126 = n4487 | n4489;
  assign n12127 = (n15648 & n4487) | (n15648 & n12126) | (n4487 & n12126);
  assign n12086 = (n4352 & n4395) | (n4352 & n12085) | (n4395 & n12085);
  assign n12131 = n4459 | n4461;
  assign n15669 = n4374 | n4459;
  assign n15670 = (n4459 & n4461) | (n4459 & n15669) | (n4461 & n15669);
  assign n15671 = (n12071 & n12131) | (n12071 & n15670) | (n12131 & n15670);
  assign n15672 = (n4376 & n12131) | (n4376 & n15670) | (n12131 & n15670);
  assign n15673 = (n12050 & n15671) | (n12050 & n15672) | (n15671 & n15672);
  assign n4536 = x61 & x80;
  assign n4537 = x60 & x81;
  assign n4538 = n4536 & n4537;
  assign n4539 = n4536 | n4537;
  assign n4540 = ~n4538 & n4539;
  assign n15678 = n4445 | n4447;
  assign n49866 = n4540 & n15678;
  assign n49867 = n4445 & n4540;
  assign n49868 = (n15650 & n49866) | (n15650 & n49867) | (n49866 & n49867);
  assign n15680 = (n4445 & n15652) | (n4445 & n15678) | (n15652 & n15678);
  assign n15682 = n4540 & n15680;
  assign n15683 = (n15617 & n49868) | (n15617 & n15682) | (n49868 & n15682);
  assign n49869 = n4540 | n15678;
  assign n49870 = n4445 | n4540;
  assign n49871 = (n15650 & n49869) | (n15650 & n49870) | (n49869 & n49870);
  assign n15685 = n4540 | n15680;
  assign n15686 = (n15617 & n49871) | (n15617 & n15685) | (n49871 & n15685);
  assign n4543 = ~n15683 & n15686;
  assign n4544 = x59 & x82;
  assign n4545 = n4543 & n4544;
  assign n4546 = n4543 | n4544;
  assign n4547 = ~n4545 & n4546;
  assign n15674 = n4452 | n4454;
  assign n15675 = (n4452 & n12089) | (n4452 & n15674) | (n12089 & n15674);
  assign n15687 = n4547 & n15675;
  assign n15676 = n4367 | n4452;
  assign n15677 = (n4452 & n4454) | (n4452 & n15676) | (n4454 & n15676);
  assign n15688 = n4547 & n15677;
  assign n15689 = (n15634 & n15687) | (n15634 & n15688) | (n15687 & n15688);
  assign n15690 = n4547 | n15675;
  assign n15691 = n4547 | n15677;
  assign n15692 = (n15634 & n15690) | (n15634 & n15691) | (n15690 & n15691);
  assign n4550 = ~n15689 & n15692;
  assign n4551 = x58 & x83;
  assign n4552 = n4550 & n4551;
  assign n4553 = n4550 | n4551;
  assign n4554 = ~n4552 & n4553;
  assign n4555 = n15673 & n4554;
  assign n4556 = n15673 | n4554;
  assign n4557 = ~n4555 & n4556;
  assign n4558 = x57 & x84;
  assign n4559 = n4557 & n4558;
  assign n4560 = n4557 | n4558;
  assign n4561 = ~n4559 & n4560;
  assign n12139 = n4466 & n4561;
  assign n12140 = (n4561 & n12111) | (n4561 & n12139) | (n12111 & n12139);
  assign n12141 = n4466 | n4561;
  assign n12142 = n12111 | n12141;
  assign n4564 = ~n12140 & n12142;
  assign n4565 = x56 & x85;
  assign n4566 = n4564 & n4565;
  assign n4567 = n4564 | n4565;
  assign n4568 = ~n4566 & n4567;
  assign n12143 = n4473 & n4568;
  assign n12144 = (n4568 & n12116) | (n4568 & n12143) | (n12116 & n12143);
  assign n12145 = n4473 | n4568;
  assign n12146 = n12116 | n12145;
  assign n4571 = ~n12144 & n12146;
  assign n4572 = x55 & x86;
  assign n4573 = n4571 & n4572;
  assign n4574 = n4571 | n4572;
  assign n4575 = ~n4573 & n4574;
  assign n12128 = n4480 | n4482;
  assign n12147 = n4575 & n12128;
  assign n12148 = n4480 & n4575;
  assign n12149 = (n12086 & n12147) | (n12086 & n12148) | (n12147 & n12148);
  assign n12150 = n4575 | n12128;
  assign n12151 = n4480 | n4575;
  assign n12152 = (n12086 & n12150) | (n12086 & n12151) | (n12150 & n12151);
  assign n4578 = ~n12149 & n12152;
  assign n4579 = x54 & x87;
  assign n4580 = n4578 & n4579;
  assign n4581 = n4578 | n4579;
  assign n4582 = ~n4580 & n4581;
  assign n4583 = n12127 & n4582;
  assign n4584 = n12127 | n4582;
  assign n4585 = ~n4583 & n4584;
  assign n4586 = x53 & x88;
  assign n4587 = n4585 & n4586;
  assign n4588 = n4585 | n4586;
  assign n4589 = ~n4587 & n4588;
  assign n4590 = n15668 & n4589;
  assign n4591 = n15668 | n4589;
  assign n4592 = ~n4590 & n4591;
  assign n4593 = x52 & x89;
  assign n4594 = n4592 & n4593;
  assign n4595 = n4592 | n4593;
  assign n4596 = ~n4594 & n4595;
  assign n4597 = n12125 & n4596;
  assign n4598 = n12125 | n4596;
  assign n4599 = ~n4597 & n4598;
  assign n4600 = x51 & x90;
  assign n4601 = n4599 & n4600;
  assign n4602 = n4599 | n4600;
  assign n4603 = ~n4601 & n4602;
  assign n4604 = n12123 & n4603;
  assign n4605 = n12123 | n4603;
  assign n4606 = ~n4604 & n4605;
  assign n4607 = x50 & x91;
  assign n4608 = n4606 & n4607;
  assign n4609 = n4606 | n4607;
  assign n4610 = ~n4608 & n4609;
  assign n4611 = n12121 & n4610;
  assign n4612 = n12121 | n4610;
  assign n4613 = ~n4611 & n4612;
  assign n4614 = x49 & x92;
  assign n4615 = n4613 & n4614;
  assign n4616 = n4613 | n4614;
  assign n4617 = ~n4615 & n4616;
  assign n4618 = n4522 & n4617;
  assign n4619 = n4522 | n4617;
  assign n4620 = ~n4618 & n4619;
  assign n4621 = x48 & x93;
  assign n4622 = n4620 & n4621;
  assign n4623 = n4620 | n4621;
  assign n4624 = ~n4622 & n4623;
  assign n12153 = n4522 | n4615;
  assign n12154 = (n4615 & n4617) | (n4615 & n12153) | (n4617 & n12153);
  assign n12155 = n4608 | n12121;
  assign n12156 = (n4608 & n4610) | (n4608 & n12155) | (n4610 & n12155);
  assign n12157 = n4601 | n12123;
  assign n12158 = (n4601 & n4603) | (n4601 & n12157) | (n4603 & n12157);
  assign n12159 = n4594 | n12125;
  assign n12160 = (n4594 & n4596) | (n4594 & n12159) | (n4596 & n12159);
  assign n12161 = n4587 | n4589;
  assign n12162 = (n15668 & n4587) | (n15668 & n12161) | (n4587 & n12161);
  assign n4637 = x62 & x80;
  assign n4638 = x61 & x81;
  assign n4639 = n4637 & n4638;
  assign n4640 = n4637 | n4638;
  assign n4641 = ~n4639 & n4640;
  assign n12169 = n4538 | n4540;
  assign n12171 = n4641 & n12169;
  assign n12172 = n4538 & n4641;
  assign n15679 = (n4445 & n15650) | (n4445 & n15678) | (n15650 & n15678);
  assign n15693 = (n12171 & n12172) | (n12171 & n15679) | (n12172 & n15679);
  assign n15694 = (n12171 & n12172) | (n12171 & n15680) | (n12172 & n15680);
  assign n15695 = (n15617 & n15693) | (n15617 & n15694) | (n15693 & n15694);
  assign n12174 = n4641 | n12169;
  assign n12175 = n4538 | n4641;
  assign n15696 = (n12174 & n12175) | (n12174 & n15679) | (n12175 & n15679);
  assign n15697 = (n12174 & n12175) | (n12174 & n15680) | (n12175 & n15680);
  assign n15698 = (n15617 & n15696) | (n15617 & n15697) | (n15696 & n15697);
  assign n4644 = ~n15695 & n15698;
  assign n4645 = x60 & x82;
  assign n4646 = n4644 & n4645;
  assign n4647 = n4644 | n4645;
  assign n4648 = ~n4646 & n4647;
  assign n12167 = n4545 | n4547;
  assign n12177 = n4648 & n12167;
  assign n12178 = n4545 & n4648;
  assign n15699 = (n12177 & n12178) | (n12177 & n15675) | (n12178 & n15675);
  assign n15700 = (n12177 & n12178) | (n12177 & n15677) | (n12178 & n15677);
  assign n15701 = (n15634 & n15699) | (n15634 & n15700) | (n15699 & n15700);
  assign n12180 = n4648 | n12167;
  assign n12181 = n4545 | n4648;
  assign n15702 = (n12180 & n12181) | (n12180 & n15675) | (n12181 & n15675);
  assign n15703 = (n12180 & n12181) | (n12180 & n15677) | (n12181 & n15677);
  assign n15704 = (n15634 & n15702) | (n15634 & n15703) | (n15702 & n15703);
  assign n4651 = ~n15701 & n15704;
  assign n4652 = x59 & x83;
  assign n4653 = n4651 & n4652;
  assign n4654 = n4651 | n4652;
  assign n4655 = ~n4653 & n4654;
  assign n12165 = n4552 | n4554;
  assign n12183 = n4655 & n12165;
  assign n12184 = n4552 & n4655;
  assign n12185 = (n15673 & n12183) | (n15673 & n12184) | (n12183 & n12184);
  assign n12186 = n4655 | n12165;
  assign n12187 = n4552 | n4655;
  assign n12188 = (n15673 & n12186) | (n15673 & n12187) | (n12186 & n12187);
  assign n4658 = ~n12185 & n12188;
  assign n4659 = x58 & x84;
  assign n4660 = n4658 & n4659;
  assign n4661 = n4658 | n4659;
  assign n4662 = ~n4660 & n4661;
  assign n12189 = n4559 & n4662;
  assign n15705 = (n4662 & n12139) | (n4662 & n12189) | (n12139 & n12189);
  assign n15706 = (n4561 & n4662) | (n4561 & n12189) | (n4662 & n12189);
  assign n15707 = (n12111 & n15705) | (n12111 & n15706) | (n15705 & n15706);
  assign n12191 = n4559 | n4662;
  assign n15708 = n12139 | n12191;
  assign n15709 = n4561 | n12191;
  assign n15710 = (n12111 & n15708) | (n12111 & n15709) | (n15708 & n15709);
  assign n4665 = ~n15707 & n15710;
  assign n4666 = x57 & x85;
  assign n4667 = n4665 & n4666;
  assign n4668 = n4665 | n4666;
  assign n4669 = ~n4667 & n4668;
  assign n12193 = n4566 & n4669;
  assign n12194 = (n4669 & n12144) | (n4669 & n12193) | (n12144 & n12193);
  assign n12195 = n4566 | n4669;
  assign n12196 = n12144 | n12195;
  assign n4672 = ~n12194 & n12196;
  assign n4673 = x56 & x86;
  assign n4674 = n4672 & n4673;
  assign n4675 = n4672 | n4673;
  assign n4676 = ~n4674 & n4675;
  assign n12197 = n4573 & n4676;
  assign n12198 = (n4676 & n12149) | (n4676 & n12197) | (n12149 & n12197);
  assign n12199 = n4573 | n4676;
  assign n12200 = n12149 | n12199;
  assign n4679 = ~n12198 & n12200;
  assign n4680 = x55 & x87;
  assign n4681 = n4679 & n4680;
  assign n4682 = n4679 | n4680;
  assign n4683 = ~n4681 & n4682;
  assign n12163 = n4580 | n4582;
  assign n12201 = n4683 & n12163;
  assign n12202 = n4580 & n4683;
  assign n12203 = (n12127 & n12201) | (n12127 & n12202) | (n12201 & n12202);
  assign n12204 = n4683 | n12163;
  assign n12205 = n4580 | n4683;
  assign n12206 = (n12127 & n12204) | (n12127 & n12205) | (n12204 & n12205);
  assign n4686 = ~n12203 & n12206;
  assign n4687 = x54 & x88;
  assign n4688 = n4686 & n4687;
  assign n4689 = n4686 | n4687;
  assign n4690 = ~n4688 & n4689;
  assign n4691 = n12162 & n4690;
  assign n4692 = n12162 | n4690;
  assign n4693 = ~n4691 & n4692;
  assign n4694 = x53 & x89;
  assign n4695 = n4693 & n4694;
  assign n4696 = n4693 | n4694;
  assign n4697 = ~n4695 & n4696;
  assign n4698 = n12160 & n4697;
  assign n4699 = n12160 | n4697;
  assign n4700 = ~n4698 & n4699;
  assign n4701 = x52 & x90;
  assign n4702 = n4700 & n4701;
  assign n4703 = n4700 | n4701;
  assign n4704 = ~n4702 & n4703;
  assign n4705 = n12158 & n4704;
  assign n4706 = n12158 | n4704;
  assign n4707 = ~n4705 & n4706;
  assign n4708 = x51 & x91;
  assign n4709 = n4707 & n4708;
  assign n4710 = n4707 | n4708;
  assign n4711 = ~n4709 & n4710;
  assign n4712 = n12156 & n4711;
  assign n4713 = n12156 | n4711;
  assign n4714 = ~n4712 & n4713;
  assign n4715 = x50 & x92;
  assign n4716 = n4714 & n4715;
  assign n4717 = n4714 | n4715;
  assign n4718 = ~n4716 & n4717;
  assign n4719 = n12154 & n4718;
  assign n4720 = n12154 | n4718;
  assign n4721 = ~n4719 & n4720;
  assign n4722 = x49 & x93;
  assign n4723 = n4721 & n4722;
  assign n4724 = n4721 | n4722;
  assign n4725 = ~n4723 & n4724;
  assign n4726 = n4622 & n4725;
  assign n4727 = n4622 | n4725;
  assign n4728 = ~n4726 & n4727;
  assign n4729 = x48 & x94;
  assign n4730 = n4728 & n4729;
  assign n4731 = n4728 | n4729;
  assign n4732 = ~n4730 & n4731;
  assign n49872 = n4621 | n4722;
  assign n49873 = (n4620 & n4722) | (n4620 & n49872) | (n4722 & n49872);
  assign n15712 = (n4622 & n4721) | (n4622 & n49873) | (n4721 & n49873);
  assign n12208 = (n4723 & n4725) | (n4723 & n15712) | (n4725 & n15712);
  assign n15713 = n4716 | n12154;
  assign n15714 = (n4716 & n4718) | (n4716 & n15713) | (n4718 & n15713);
  assign n4735 = n4709 | n4712;
  assign n4736 = n4702 | n4705;
  assign n12212 = n4660 | n4662;
  assign n15715 = n4559 | n4660;
  assign n15716 = (n4660 & n4662) | (n4660 & n15715) | (n4662 & n15715);
  assign n15717 = (n12139 & n12212) | (n12139 & n15716) | (n12212 & n15716);
  assign n15718 = (n4561 & n12212) | (n4561 & n15716) | (n12212 & n15716);
  assign n15719 = (n12111 & n15717) | (n12111 & n15718) | (n15717 & n15718);
  assign n15720 = n4646 | n4648;
  assign n15721 = (n4646 & n12167) | (n4646 & n15720) | (n12167 & n15720);
  assign n15722 = n4545 | n4646;
  assign n15723 = (n4646 & n4648) | (n4646 & n15722) | (n4648 & n15722);
  assign n15724 = (n15675 & n15721) | (n15675 & n15723) | (n15721 & n15723);
  assign n15725 = (n15677 & n15721) | (n15677 & n15723) | (n15721 & n15723);
  assign n15726 = (n15634 & n15724) | (n15634 & n15725) | (n15724 & n15725);
  assign n4746 = x63 & x80;
  assign n4747 = x62 & x81;
  assign n4748 = n4746 & n4747;
  assign n4749 = n4746 | n4747;
  assign n4750 = ~n4748 & n4749;
  assign n15727 = n4639 | n4641;
  assign n15728 = (n4639 & n12169) | (n4639 & n15727) | (n12169 & n15727);
  assign n12220 = n4750 & n15728;
  assign n15729 = n4538 | n4639;
  assign n15730 = (n4639 & n4641) | (n4639 & n15729) | (n4641 & n15729);
  assign n12221 = n4750 & n15730;
  assign n15731 = (n12220 & n12221) | (n12220 & n15679) | (n12221 & n15679);
  assign n15732 = (n12220 & n12221) | (n12220 & n15680) | (n12221 & n15680);
  assign n15733 = (n15617 & n15731) | (n15617 & n15732) | (n15731 & n15732);
  assign n12223 = n4750 | n15728;
  assign n12224 = n4750 | n15730;
  assign n15734 = (n12223 & n12224) | (n12223 & n15679) | (n12224 & n15679);
  assign n15735 = (n12223 & n12224) | (n12223 & n15680) | (n12224 & n15680);
  assign n15736 = (n15617 & n15734) | (n15617 & n15735) | (n15734 & n15735);
  assign n4753 = ~n15733 & n15736;
  assign n4754 = x61 & x82;
  assign n4755 = n4753 & n4754;
  assign n4756 = n4753 | n4754;
  assign n4757 = ~n4755 & n4756;
  assign n4758 = n15726 & n4757;
  assign n4759 = n15726 | n4757;
  assign n4760 = ~n4758 & n4759;
  assign n4761 = x60 & x83;
  assign n4762 = n4760 & n4761;
  assign n4763 = n4760 | n4761;
  assign n4764 = ~n4762 & n4763;
  assign n12226 = n4653 & n4764;
  assign n15737 = (n4764 & n12183) | (n4764 & n12226) | (n12183 & n12226);
  assign n15738 = (n4764 & n12184) | (n4764 & n12226) | (n12184 & n12226);
  assign n15739 = (n15673 & n15737) | (n15673 & n15738) | (n15737 & n15738);
  assign n12228 = n4653 | n4764;
  assign n15740 = n12183 | n12228;
  assign n15741 = n12184 | n12228;
  assign n15742 = (n15673 & n15740) | (n15673 & n15741) | (n15740 & n15741);
  assign n4767 = ~n15739 & n15742;
  assign n4768 = x59 & x84;
  assign n4769 = n4767 & n4768;
  assign n4770 = n4767 | n4768;
  assign n4771 = ~n4769 & n4770;
  assign n4772 = n15719 & n4771;
  assign n4773 = n15719 | n4771;
  assign n4774 = ~n4772 & n4773;
  assign n4775 = x58 & x85;
  assign n4776 = n4774 & n4775;
  assign n4777 = n4774 | n4775;
  assign n4778 = ~n4776 & n4777;
  assign n12230 = n4667 & n4778;
  assign n12231 = (n4778 & n12194) | (n4778 & n12230) | (n12194 & n12230);
  assign n12232 = n4667 | n4778;
  assign n12233 = n12194 | n12232;
  assign n4781 = ~n12231 & n12233;
  assign n4782 = x57 & x86;
  assign n4783 = n4781 & n4782;
  assign n4784 = n4781 | n4782;
  assign n4785 = ~n4783 & n4784;
  assign n12234 = n4674 & n4785;
  assign n12235 = (n4785 & n12198) | (n4785 & n12234) | (n12198 & n12234);
  assign n12236 = n4674 | n4785;
  assign n12237 = n12198 | n12236;
  assign n4788 = ~n12235 & n12237;
  assign n4789 = x56 & x87;
  assign n4790 = n4788 & n4789;
  assign n4791 = n4788 | n4789;
  assign n4792 = ~n4790 & n4791;
  assign n12238 = n4681 & n4792;
  assign n12239 = (n4792 & n12203) | (n4792 & n12238) | (n12203 & n12238);
  assign n12240 = n4681 | n4792;
  assign n12241 = n12203 | n12240;
  assign n4795 = ~n12239 & n12241;
  assign n4796 = x55 & x88;
  assign n4797 = n4795 & n4796;
  assign n4798 = n4795 | n4796;
  assign n4799 = ~n4797 & n4798;
  assign n12209 = n4688 | n4690;
  assign n12242 = n4799 & n12209;
  assign n12243 = n4688 & n4799;
  assign n12244 = (n12162 & n12242) | (n12162 & n12243) | (n12242 & n12243);
  assign n12245 = n4799 | n12209;
  assign n12246 = n4688 | n4799;
  assign n12247 = (n12162 & n12245) | (n12162 & n12246) | (n12245 & n12246);
  assign n4802 = ~n12244 & n12247;
  assign n4803 = x54 & x89;
  assign n4804 = n4802 & n4803;
  assign n4805 = n4802 | n4803;
  assign n4806 = ~n4804 & n4805;
  assign n12248 = n4695 & n4806;
  assign n12249 = (n4698 & n4806) | (n4698 & n12248) | (n4806 & n12248);
  assign n12250 = n4695 | n4806;
  assign n12251 = n4698 | n12250;
  assign n4809 = ~n12249 & n12251;
  assign n4810 = x53 & x90;
  assign n4811 = n4809 & n4810;
  assign n4812 = n4809 | n4810;
  assign n4813 = ~n4811 & n4812;
  assign n4814 = n4736 & n4813;
  assign n4815 = n4736 | n4813;
  assign n4816 = ~n4814 & n4815;
  assign n4817 = x52 & x91;
  assign n4818 = n4816 & n4817;
  assign n4819 = n4816 | n4817;
  assign n4820 = ~n4818 & n4819;
  assign n4821 = n4735 & n4820;
  assign n4822 = n4735 | n4820;
  assign n4823 = ~n4821 & n4822;
  assign n4824 = x51 & x92;
  assign n4825 = n4823 & n4824;
  assign n4826 = n4823 | n4824;
  assign n4827 = ~n4825 & n4826;
  assign n4828 = n15714 & n4827;
  assign n4829 = n15714 | n4827;
  assign n4830 = ~n4828 & n4829;
  assign n4831 = x50 & x93;
  assign n4832 = n4830 & n4831;
  assign n4833 = n4830 | n4831;
  assign n4834 = ~n4832 & n4833;
  assign n4835 = n12208 & n4834;
  assign n4836 = n12208 | n4834;
  assign n4837 = ~n4835 & n4836;
  assign n4838 = x49 & x94;
  assign n4839 = n4837 & n4838;
  assign n4840 = n4837 | n4838;
  assign n4841 = ~n4839 & n4840;
  assign n4842 = n4730 & n4841;
  assign n4843 = n4730 | n4841;
  assign n4844 = ~n4842 & n4843;
  assign n4845 = x48 & x95;
  assign n4846 = n4844 & n4845;
  assign n4847 = n4844 | n4845;
  assign n4848 = ~n4846 & n4847;
  assign n49874 = n4729 | n4838;
  assign n49875 = (n4728 & n4838) | (n4728 & n49874) | (n4838 & n49874);
  assign n15744 = (n4730 & n4837) | (n4730 & n49875) | (n4837 & n49875);
  assign n12253 = (n4839 & n4841) | (n4839 & n15744) | (n4841 & n15744);
  assign n12254 = n4832 | n12208;
  assign n12255 = (n4832 & n4834) | (n4832 & n12254) | (n4834 & n12254);
  assign n15745 = n4825 | n15714;
  assign n15746 = (n4825 & n4827) | (n4825 & n15745) | (n4827 & n15745);
  assign n4852 = n4818 | n4821;
  assign n12256 = n4811 | n4813;
  assign n12257 = (n4736 & n4811) | (n4736 & n12256) | (n4811 & n12256);
  assign n12261 = n4762 | n4764;
  assign n15747 = n4653 | n4762;
  assign n15748 = (n4762 & n4764) | (n4762 & n15747) | (n4764 & n15747);
  assign n15749 = (n12183 & n12261) | (n12183 & n15748) | (n12261 & n15748);
  assign n15750 = (n12184 & n12261) | (n12184 & n15748) | (n12261 & n15748);
  assign n15751 = (n15673 & n15749) | (n15673 & n15750) | (n15749 & n15750);
  assign n4863 = x64 & x80;
  assign n4864 = x63 & x81;
  assign n4865 = n4863 & n4864;
  assign n4866 = n4863 | n4864;
  assign n4867 = ~n4865 & n4866;
  assign n15752 = n4748 | n4750;
  assign n15757 = (n4748 & n15730) | (n4748 & n15752) | (n15730 & n15752);
  assign n12269 = n4867 & n15757;
  assign n15754 = n4867 & n15752;
  assign n15755 = n4748 & n4867;
  assign n15756 = (n15728 & n15754) | (n15728 & n15755) | (n15754 & n15755);
  assign n15758 = (n12269 & n15679) | (n12269 & n15756) | (n15679 & n15756);
  assign n15759 = (n12269 & n15680) | (n12269 & n15756) | (n15680 & n15756);
  assign n15760 = (n15617 & n15758) | (n15617 & n15759) | (n15758 & n15759);
  assign n12272 = n4867 | n15757;
  assign n15761 = n4867 | n15752;
  assign n15762 = n4748 | n4867;
  assign n15763 = (n15728 & n15761) | (n15728 & n15762) | (n15761 & n15762);
  assign n15764 = (n12272 & n15679) | (n12272 & n15763) | (n15679 & n15763);
  assign n15765 = (n12272 & n15680) | (n12272 & n15763) | (n15680 & n15763);
  assign n15766 = (n15617 & n15764) | (n15617 & n15765) | (n15764 & n15765);
  assign n4870 = ~n15760 & n15766;
  assign n4871 = x62 & x82;
  assign n4872 = n4870 & n4871;
  assign n4873 = n4870 | n4871;
  assign n4874 = ~n4872 & n4873;
  assign n12263 = n4755 | n4757;
  assign n12274 = n4874 & n12263;
  assign n12275 = n4755 & n4874;
  assign n12276 = (n15726 & n12274) | (n15726 & n12275) | (n12274 & n12275);
  assign n12277 = n4874 | n12263;
  assign n12278 = n4755 | n4874;
  assign n12279 = (n15726 & n12277) | (n15726 & n12278) | (n12277 & n12278);
  assign n4877 = ~n12276 & n12279;
  assign n4878 = x61 & x83;
  assign n4879 = n4877 & n4878;
  assign n4880 = n4877 | n4878;
  assign n4881 = ~n4879 & n4880;
  assign n4882 = n15751 & n4881;
  assign n4883 = n15751 | n4881;
  assign n4884 = ~n4882 & n4883;
  assign n4885 = x60 & x84;
  assign n4886 = n4884 & n4885;
  assign n4887 = n4884 | n4885;
  assign n4888 = ~n4886 & n4887;
  assign n12258 = n4769 | n4771;
  assign n12280 = n4888 & n12258;
  assign n12281 = n4769 & n4888;
  assign n12282 = (n15719 & n12280) | (n15719 & n12281) | (n12280 & n12281);
  assign n12283 = n4888 | n12258;
  assign n12284 = n4769 | n4888;
  assign n12285 = (n15719 & n12283) | (n15719 & n12284) | (n12283 & n12284);
  assign n4891 = ~n12282 & n12285;
  assign n4892 = x59 & x85;
  assign n4893 = n4891 & n4892;
  assign n4894 = n4891 | n4892;
  assign n4895 = ~n4893 & n4894;
  assign n12286 = n4776 & n4895;
  assign n15767 = (n4895 & n12230) | (n4895 & n12286) | (n12230 & n12286);
  assign n15768 = (n4778 & n4895) | (n4778 & n12286) | (n4895 & n12286);
  assign n15769 = (n12194 & n15767) | (n12194 & n15768) | (n15767 & n15768);
  assign n12288 = n4776 | n4895;
  assign n15770 = n12230 | n12288;
  assign n15771 = n4778 | n12288;
  assign n15772 = (n12194 & n15770) | (n12194 & n15771) | (n15770 & n15771);
  assign n4898 = ~n15769 & n15772;
  assign n4899 = x58 & x86;
  assign n4900 = n4898 & n4899;
  assign n4901 = n4898 | n4899;
  assign n4902 = ~n4900 & n4901;
  assign n12290 = n4783 & n4902;
  assign n12291 = (n4902 & n12235) | (n4902 & n12290) | (n12235 & n12290);
  assign n12292 = n4783 | n4902;
  assign n12293 = n12235 | n12292;
  assign n4905 = ~n12291 & n12293;
  assign n4906 = x57 & x87;
  assign n4907 = n4905 & n4906;
  assign n4908 = n4905 | n4906;
  assign n4909 = ~n4907 & n4908;
  assign n12294 = n4790 & n4909;
  assign n12295 = (n4909 & n12239) | (n4909 & n12294) | (n12239 & n12294);
  assign n12296 = n4790 | n4909;
  assign n12297 = n12239 | n12296;
  assign n4912 = ~n12295 & n12297;
  assign n4913 = x56 & x88;
  assign n4914 = n4912 & n4913;
  assign n4915 = n4912 | n4913;
  assign n4916 = ~n4914 & n4915;
  assign n12298 = n4797 & n4916;
  assign n12299 = (n4916 & n12244) | (n4916 & n12298) | (n12244 & n12298);
  assign n12300 = n4797 | n4916;
  assign n12301 = n12244 | n12300;
  assign n4919 = ~n12299 & n12301;
  assign n4920 = x55 & x89;
  assign n4921 = n4919 & n4920;
  assign n4922 = n4919 | n4920;
  assign n4923 = ~n4921 & n4922;
  assign n12302 = n4804 & n4923;
  assign n12303 = (n4923 & n12249) | (n4923 & n12302) | (n12249 & n12302);
  assign n12304 = n4804 | n4923;
  assign n12305 = n12249 | n12304;
  assign n4926 = ~n12303 & n12305;
  assign n4927 = x54 & x90;
  assign n4928 = n4926 & n4927;
  assign n4929 = n4926 | n4927;
  assign n4930 = ~n4928 & n4929;
  assign n4931 = n12257 & n4930;
  assign n4932 = n12257 | n4930;
  assign n4933 = ~n4931 & n4932;
  assign n4934 = x53 & x91;
  assign n4935 = n4933 & n4934;
  assign n4936 = n4933 | n4934;
  assign n4937 = ~n4935 & n4936;
  assign n4938 = n4852 & n4937;
  assign n4939 = n4852 | n4937;
  assign n4940 = ~n4938 & n4939;
  assign n4941 = x52 & x92;
  assign n4942 = n4940 & n4941;
  assign n4943 = n4940 | n4941;
  assign n4944 = ~n4942 & n4943;
  assign n4945 = n15746 & n4944;
  assign n4946 = n15746 | n4944;
  assign n4947 = ~n4945 & n4946;
  assign n4948 = x51 & x93;
  assign n4949 = n4947 & n4948;
  assign n4950 = n4947 | n4948;
  assign n4951 = ~n4949 & n4950;
  assign n4952 = n12255 & n4951;
  assign n4953 = n12255 | n4951;
  assign n4954 = ~n4952 & n4953;
  assign n4955 = x50 & x94;
  assign n4956 = n4954 & n4955;
  assign n4957 = n4954 | n4955;
  assign n4958 = ~n4956 & n4957;
  assign n4959 = n12253 & n4958;
  assign n4960 = n12253 | n4958;
  assign n4961 = ~n4959 & n4960;
  assign n4962 = x49 & x95;
  assign n4963 = n4961 & n4962;
  assign n4964 = n4961 | n4962;
  assign n4965 = ~n4963 & n4964;
  assign n4966 = n4846 & n4965;
  assign n4967 = n4846 | n4965;
  assign n4968 = ~n4966 & n4967;
  assign n4969 = x48 & x96;
  assign n4970 = n4968 & n4969;
  assign n4971 = n4968 | n4969;
  assign n4972 = ~n4970 & n4971;
  assign n49876 = n4845 | n4962;
  assign n49877 = (n4844 & n4962) | (n4844 & n49876) | (n4962 & n49876);
  assign n15774 = (n4846 & n4961) | (n4846 & n49877) | (n4961 & n49877);
  assign n12307 = (n4963 & n4965) | (n4963 & n15774) | (n4965 & n15774);
  assign n12308 = n4956 | n12253;
  assign n12309 = (n4956 & n4958) | (n4956 & n12308) | (n4958 & n12308);
  assign n12310 = n4949 | n12255;
  assign n12311 = (n4949 & n4951) | (n4949 & n12310) | (n4951 & n12310);
  assign n15775 = n4942 | n15746;
  assign n15776 = (n4942 & n4944) | (n4942 & n15775) | (n4944 & n15775);
  assign n12312 = n4935 | n4937;
  assign n12313 = (n4852 & n4935) | (n4852 & n12312) | (n4935 & n12312);
  assign n12314 = n4928 | n4930;
  assign n12315 = (n4928 & n12257) | (n4928 & n12314) | (n12257 & n12314);
  assign n12317 = n4893 | n4895;
  assign n15777 = n4776 | n4893;
  assign n15778 = (n4893 & n4895) | (n4893 & n15777) | (n4895 & n15777);
  assign n15779 = (n12230 & n12317) | (n12230 & n15778) | (n12317 & n15778);
  assign n15780 = (n4778 & n12317) | (n4778 & n15778) | (n12317 & n15778);
  assign n15781 = (n12194 & n15779) | (n12194 & n15780) | (n15779 & n15780);
  assign n4988 = x65 & x80;
  assign n4989 = x64 & x81;
  assign n4990 = n4988 & n4989;
  assign n4991 = n4988 | n4989;
  assign n4992 = ~n4990 & n4991;
  assign n12324 = n4865 & n4992;
  assign n12325 = (n4992 & n15760) | (n4992 & n12324) | (n15760 & n12324);
  assign n12326 = n4865 | n4992;
  assign n12327 = n15760 | n12326;
  assign n4995 = ~n12325 & n12327;
  assign n4996 = x63 & x82;
  assign n4997 = n4995 & n4996;
  assign n4998 = n4995 | n4996;
  assign n4999 = ~n4997 & n4998;
  assign n15782 = n4872 | n4874;
  assign n15783 = (n4872 & n12263) | (n4872 & n15782) | (n12263 & n15782);
  assign n12328 = n4999 & n15783;
  assign n15784 = n4755 | n4872;
  assign n15785 = (n4872 & n4874) | (n4872 & n15784) | (n4874 & n15784);
  assign n12329 = n4999 & n15785;
  assign n12330 = (n15726 & n12328) | (n15726 & n12329) | (n12328 & n12329);
  assign n12331 = n4999 | n15783;
  assign n12332 = n4999 | n15785;
  assign n12333 = (n15726 & n12331) | (n15726 & n12332) | (n12331 & n12332);
  assign n5002 = ~n12330 & n12333;
  assign n5003 = x62 & x83;
  assign n5004 = n5002 & n5003;
  assign n5005 = n5002 | n5003;
  assign n5006 = ~n5004 & n5005;
  assign n12319 = n4879 | n4881;
  assign n12334 = n5006 & n12319;
  assign n12335 = n4879 & n5006;
  assign n12336 = (n15751 & n12334) | (n15751 & n12335) | (n12334 & n12335);
  assign n12337 = n5006 | n12319;
  assign n12338 = n4879 | n5006;
  assign n12339 = (n15751 & n12337) | (n15751 & n12338) | (n12337 & n12338);
  assign n5009 = ~n12336 & n12339;
  assign n5010 = x61 & x84;
  assign n5011 = n5009 & n5010;
  assign n5012 = n5009 | n5010;
  assign n5013 = ~n5011 & n5012;
  assign n12340 = n4886 & n5013;
  assign n15786 = (n5013 & n12281) | (n5013 & n12340) | (n12281 & n12340);
  assign n15787 = (n5013 & n12280) | (n5013 & n12340) | (n12280 & n12340);
  assign n15788 = (n15719 & n15786) | (n15719 & n15787) | (n15786 & n15787);
  assign n12342 = n4886 | n5013;
  assign n15789 = n12281 | n12342;
  assign n15790 = n12280 | n12342;
  assign n15791 = (n15719 & n15789) | (n15719 & n15790) | (n15789 & n15790);
  assign n5016 = ~n15788 & n15791;
  assign n5017 = x60 & x85;
  assign n5018 = n5016 & n5017;
  assign n5019 = n5016 | n5017;
  assign n5020 = ~n5018 & n5019;
  assign n5021 = n15781 & n5020;
  assign n5022 = n15781 | n5020;
  assign n5023 = ~n5021 & n5022;
  assign n5024 = x59 & x86;
  assign n5025 = n5023 & n5024;
  assign n5026 = n5023 | n5024;
  assign n5027 = ~n5025 & n5026;
  assign n12344 = n4900 & n5027;
  assign n12345 = (n5027 & n12291) | (n5027 & n12344) | (n12291 & n12344);
  assign n12346 = n4900 | n5027;
  assign n12347 = n12291 | n12346;
  assign n5030 = ~n12345 & n12347;
  assign n5031 = x58 & x87;
  assign n5032 = n5030 & n5031;
  assign n5033 = n5030 | n5031;
  assign n5034 = ~n5032 & n5033;
  assign n12348 = n4907 & n5034;
  assign n12349 = (n5034 & n12295) | (n5034 & n12348) | (n12295 & n12348);
  assign n12350 = n4907 | n5034;
  assign n12351 = n12295 | n12350;
  assign n5037 = ~n12349 & n12351;
  assign n5038 = x57 & x88;
  assign n5039 = n5037 & n5038;
  assign n5040 = n5037 | n5038;
  assign n5041 = ~n5039 & n5040;
  assign n12352 = n4914 & n5041;
  assign n12353 = (n5041 & n12299) | (n5041 & n12352) | (n12299 & n12352);
  assign n12354 = n4914 | n5041;
  assign n12355 = n12299 | n12354;
  assign n5044 = ~n12353 & n12355;
  assign n5045 = x56 & x89;
  assign n5046 = n5044 & n5045;
  assign n5047 = n5044 | n5045;
  assign n5048 = ~n5046 & n5047;
  assign n12356 = n4921 & n5048;
  assign n12357 = (n5048 & n12303) | (n5048 & n12356) | (n12303 & n12356);
  assign n12358 = n4921 | n5048;
  assign n12359 = n12303 | n12358;
  assign n5051 = ~n12357 & n12359;
  assign n5052 = x55 & x90;
  assign n5053 = n5051 & n5052;
  assign n5054 = n5051 | n5052;
  assign n5055 = ~n5053 & n5054;
  assign n5056 = n12315 & n5055;
  assign n5057 = n12315 | n5055;
  assign n5058 = ~n5056 & n5057;
  assign n5059 = x54 & x91;
  assign n5060 = n5058 & n5059;
  assign n5061 = n5058 | n5059;
  assign n5062 = ~n5060 & n5061;
  assign n5063 = n12313 & n5062;
  assign n5064 = n12313 | n5062;
  assign n5065 = ~n5063 & n5064;
  assign n5066 = x53 & x92;
  assign n5067 = n5065 & n5066;
  assign n5068 = n5065 | n5066;
  assign n5069 = ~n5067 & n5068;
  assign n5070 = n15776 & n5069;
  assign n5071 = n15776 | n5069;
  assign n5072 = ~n5070 & n5071;
  assign n5073 = x52 & x93;
  assign n5074 = n5072 & n5073;
  assign n5075 = n5072 | n5073;
  assign n5076 = ~n5074 & n5075;
  assign n5077 = n12311 & n5076;
  assign n5078 = n12311 | n5076;
  assign n5079 = ~n5077 & n5078;
  assign n5080 = x51 & x94;
  assign n5081 = n5079 & n5080;
  assign n5082 = n5079 | n5080;
  assign n5083 = ~n5081 & n5082;
  assign n5084 = n12309 & n5083;
  assign n5085 = n12309 | n5083;
  assign n5086 = ~n5084 & n5085;
  assign n5087 = x50 & x95;
  assign n5088 = n5086 & n5087;
  assign n5089 = n5086 | n5087;
  assign n5090 = ~n5088 & n5089;
  assign n5091 = n12307 & n5090;
  assign n5092 = n12307 | n5090;
  assign n5093 = ~n5091 & n5092;
  assign n5094 = x49 & x96;
  assign n5095 = n5093 & n5094;
  assign n5096 = n5093 | n5094;
  assign n5097 = ~n5095 & n5096;
  assign n5098 = n4970 & n5097;
  assign n5099 = n4970 | n5097;
  assign n5100 = ~n5098 & n5099;
  assign n5101 = x48 & x97;
  assign n5102 = n5100 & n5101;
  assign n5103 = n5100 | n5101;
  assign n5104 = ~n5102 & n5103;
  assign n12360 = n4970 | n5095;
  assign n12361 = (n5095 & n5097) | (n5095 & n12360) | (n5097 & n12360);
  assign n12362 = n5088 | n12307;
  assign n12363 = (n5088 & n5090) | (n5088 & n12362) | (n5090 & n12362);
  assign n12364 = n5081 | n12309;
  assign n12365 = (n5081 & n5083) | (n5081 & n12364) | (n5083 & n12364);
  assign n12366 = n5074 | n12311;
  assign n12367 = (n5074 & n5076) | (n5074 & n12366) | (n5076 & n12366);
  assign n12368 = n5067 | n5069;
  assign n12369 = (n15776 & n5067) | (n15776 & n12368) | (n5067 & n12368);
  assign n12370 = n5060 | n5062;
  assign n12371 = (n5060 & n12313) | (n5060 & n12370) | (n12313 & n12370);
  assign n12372 = n5053 | n5055;
  assign n12373 = (n5053 & n12315) | (n5053 & n12372) | (n12315 & n12372);
  assign n12377 = n5011 | n5013;
  assign n15792 = n4886 | n5011;
  assign n15793 = (n5011 & n5013) | (n5011 & n15792) | (n5013 & n15792);
  assign n15794 = (n12281 & n12377) | (n12281 & n15793) | (n12377 & n15793);
  assign n15795 = (n12280 & n12377) | (n12280 & n15793) | (n12377 & n15793);
  assign n15796 = (n15719 & n15794) | (n15719 & n15795) | (n15794 & n15795);
  assign n5121 = x66 & x80;
  assign n5122 = x65 & x81;
  assign n5123 = n5121 & n5122;
  assign n5124 = n5121 | n5122;
  assign n5125 = ~n5123 & n5124;
  assign n15801 = n4865 | n4990;
  assign n15802 = (n4990 & n4992) | (n4990 & n15801) | (n4992 & n15801);
  assign n12385 = n5125 & n15802;
  assign n12383 = n4990 | n4992;
  assign n12386 = n5125 & n12383;
  assign n12387 = (n15760 & n12385) | (n15760 & n12386) | (n12385 & n12386);
  assign n12388 = n5125 | n15802;
  assign n12389 = n5125 | n12383;
  assign n12390 = (n15760 & n12388) | (n15760 & n12389) | (n12388 & n12389);
  assign n5128 = ~n12387 & n12390;
  assign n5129 = x64 & x82;
  assign n5130 = n5128 & n5129;
  assign n5131 = n5128 | n5129;
  assign n5132 = ~n5130 & n5131;
  assign n12391 = n4997 & n5132;
  assign n15803 = (n5132 & n12328) | (n5132 & n12391) | (n12328 & n12391);
  assign n15804 = (n5132 & n12329) | (n5132 & n12391) | (n12329 & n12391);
  assign n15805 = (n15726 & n15803) | (n15726 & n15804) | (n15803 & n15804);
  assign n12393 = n4997 | n5132;
  assign n15806 = n12328 | n12393;
  assign n15807 = n12329 | n12393;
  assign n15808 = (n15726 & n15806) | (n15726 & n15807) | (n15806 & n15807);
  assign n5135 = ~n15805 & n15808;
  assign n5136 = x63 & x83;
  assign n5137 = n5135 & n5136;
  assign n5138 = n5135 | n5136;
  assign n5139 = ~n5137 & n5138;
  assign n15797 = n5004 | n5006;
  assign n15798 = (n5004 & n12319) | (n5004 & n15797) | (n12319 & n15797);
  assign n15809 = n5139 & n15798;
  assign n15799 = n4879 | n5004;
  assign n15800 = (n5004 & n5006) | (n5004 & n15799) | (n5006 & n15799);
  assign n15810 = n5139 & n15800;
  assign n15811 = (n15751 & n15809) | (n15751 & n15810) | (n15809 & n15810);
  assign n15812 = n5139 | n15798;
  assign n15813 = n5139 | n15800;
  assign n15814 = (n15751 & n15812) | (n15751 & n15813) | (n15812 & n15813);
  assign n5142 = ~n15811 & n15814;
  assign n5143 = x62 & x84;
  assign n5144 = n5142 & n5143;
  assign n5145 = n5142 | n5143;
  assign n5146 = ~n5144 & n5145;
  assign n5147 = n15796 & n5146;
  assign n5148 = n15796 | n5146;
  assign n5149 = ~n5147 & n5148;
  assign n5150 = x61 & x85;
  assign n5151 = n5149 & n5150;
  assign n5152 = n5149 | n5150;
  assign n5153 = ~n5151 & n5152;
  assign n12374 = n5018 | n5020;
  assign n12395 = n5153 & n12374;
  assign n12396 = n5018 & n5153;
  assign n12397 = (n15781 & n12395) | (n15781 & n12396) | (n12395 & n12396);
  assign n12398 = n5153 | n12374;
  assign n12399 = n5018 | n5153;
  assign n12400 = (n15781 & n12398) | (n15781 & n12399) | (n12398 & n12399);
  assign n5156 = ~n12397 & n12400;
  assign n5157 = x60 & x86;
  assign n5158 = n5156 & n5157;
  assign n5159 = n5156 | n5157;
  assign n5160 = ~n5158 & n5159;
  assign n12401 = n5025 & n5160;
  assign n15815 = (n5160 & n12344) | (n5160 & n12401) | (n12344 & n12401);
  assign n15816 = (n5027 & n5160) | (n5027 & n12401) | (n5160 & n12401);
  assign n15817 = (n12291 & n15815) | (n12291 & n15816) | (n15815 & n15816);
  assign n12403 = n5025 | n5160;
  assign n15818 = n12344 | n12403;
  assign n15819 = n5027 | n12403;
  assign n15820 = (n12291 & n15818) | (n12291 & n15819) | (n15818 & n15819);
  assign n5163 = ~n15817 & n15820;
  assign n5164 = x59 & x87;
  assign n5165 = n5163 & n5164;
  assign n5166 = n5163 | n5164;
  assign n5167 = ~n5165 & n5166;
  assign n12405 = n5032 & n5167;
  assign n12406 = (n5167 & n12349) | (n5167 & n12405) | (n12349 & n12405);
  assign n12407 = n5032 | n5167;
  assign n12408 = n12349 | n12407;
  assign n5170 = ~n12406 & n12408;
  assign n5171 = x58 & x88;
  assign n5172 = n5170 & n5171;
  assign n5173 = n5170 | n5171;
  assign n5174 = ~n5172 & n5173;
  assign n12409 = n5039 & n5174;
  assign n12410 = (n5174 & n12353) | (n5174 & n12409) | (n12353 & n12409);
  assign n12411 = n5039 | n5174;
  assign n12412 = n12353 | n12411;
  assign n5177 = ~n12410 & n12412;
  assign n5178 = x57 & x89;
  assign n5179 = n5177 & n5178;
  assign n5180 = n5177 | n5178;
  assign n5181 = ~n5179 & n5180;
  assign n12413 = n5046 & n5181;
  assign n12414 = (n5181 & n12357) | (n5181 & n12413) | (n12357 & n12413);
  assign n12415 = n5046 | n5181;
  assign n12416 = n12357 | n12415;
  assign n5184 = ~n12414 & n12416;
  assign n5185 = x56 & x90;
  assign n5186 = n5184 & n5185;
  assign n5187 = n5184 | n5185;
  assign n5188 = ~n5186 & n5187;
  assign n5189 = n12373 & n5188;
  assign n5190 = n12373 | n5188;
  assign n5191 = ~n5189 & n5190;
  assign n5192 = x55 & x91;
  assign n5193 = n5191 & n5192;
  assign n5194 = n5191 | n5192;
  assign n5195 = ~n5193 & n5194;
  assign n5196 = n12371 & n5195;
  assign n5197 = n12371 | n5195;
  assign n5198 = ~n5196 & n5197;
  assign n5199 = x54 & x92;
  assign n5200 = n5198 & n5199;
  assign n5201 = n5198 | n5199;
  assign n5202 = ~n5200 & n5201;
  assign n5203 = n12369 & n5202;
  assign n5204 = n12369 | n5202;
  assign n5205 = ~n5203 & n5204;
  assign n5206 = x53 & x93;
  assign n5207 = n5205 & n5206;
  assign n5208 = n5205 | n5206;
  assign n5209 = ~n5207 & n5208;
  assign n5210 = n12367 & n5209;
  assign n5211 = n12367 | n5209;
  assign n5212 = ~n5210 & n5211;
  assign n5213 = x52 & x94;
  assign n5214 = n5212 & n5213;
  assign n5215 = n5212 | n5213;
  assign n5216 = ~n5214 & n5215;
  assign n5217 = n12365 & n5216;
  assign n5218 = n12365 | n5216;
  assign n5219 = ~n5217 & n5218;
  assign n5220 = x51 & x95;
  assign n5221 = n5219 & n5220;
  assign n5222 = n5219 | n5220;
  assign n5223 = ~n5221 & n5222;
  assign n5224 = n12363 & n5223;
  assign n5225 = n12363 | n5223;
  assign n5226 = ~n5224 & n5225;
  assign n5227 = x50 & x96;
  assign n5228 = n5226 & n5227;
  assign n5229 = n5226 | n5227;
  assign n5230 = ~n5228 & n5229;
  assign n5231 = n12361 & n5230;
  assign n5232 = n12361 | n5230;
  assign n5233 = ~n5231 & n5232;
  assign n5234 = x49 & x97;
  assign n5235 = n5233 & n5234;
  assign n5236 = n5233 | n5234;
  assign n5237 = ~n5235 & n5236;
  assign n5238 = n5102 & n5237;
  assign n5239 = n5102 | n5237;
  assign n5240 = ~n5238 & n5239;
  assign n5241 = x48 & x98;
  assign n5242 = n5240 & n5241;
  assign n5243 = n5240 | n5241;
  assign n5244 = ~n5242 & n5243;
  assign n49878 = n5101 | n5234;
  assign n49879 = (n5100 & n5234) | (n5100 & n49878) | (n5234 & n49878);
  assign n15822 = (n5102 & n5233) | (n5102 & n49879) | (n5233 & n49879);
  assign n12418 = (n5235 & n5237) | (n5235 & n15822) | (n5237 & n15822);
  assign n15823 = n5228 | n12361;
  assign n15824 = (n5228 & n5230) | (n5228 & n15823) | (n5230 & n15823);
  assign n5247 = n5221 | n5224;
  assign n5248 = n5214 | n5217;
  assign n5249 = n5207 | n5210;
  assign n12419 = n5200 | n5202;
  assign n12420 = (n5200 & n12369) | (n5200 & n12419) | (n12369 & n12419);
  assign n12421 = n5193 | n5195;
  assign n12422 = (n5193 & n12371) | (n5193 & n12421) | (n12371 & n12421);
  assign n12423 = n5186 | n5188;
  assign n12424 = (n5186 & n12373) | (n5186 & n12423) | (n12373 & n12423);
  assign n12426 = n5158 | n5160;
  assign n15825 = n5025 | n5158;
  assign n15826 = (n5158 & n5160) | (n5158 & n15825) | (n5160 & n15825);
  assign n15827 = (n12344 & n12426) | (n12344 & n15826) | (n12426 & n15826);
  assign n15828 = (n5027 & n12426) | (n5027 & n15826) | (n12426 & n15826);
  assign n15829 = (n12291 & n15827) | (n12291 & n15828) | (n15827 & n15828);
  assign n5262 = x67 & x80;
  assign n5263 = x66 & x81;
  assign n5264 = n5262 & n5263;
  assign n5265 = n5262 | n5263;
  assign n5266 = ~n5264 & n5265;
  assign n15830 = n5123 | n5125;
  assign n15831 = (n5123 & n15802) | (n5123 & n15830) | (n15802 & n15830);
  assign n12438 = n5266 & n15831;
  assign n15832 = (n5123 & n12383) | (n5123 & n15830) | (n12383 & n15830);
  assign n12439 = n5266 & n15832;
  assign n12440 = (n15760 & n12438) | (n15760 & n12439) | (n12438 & n12439);
  assign n12441 = n5266 | n15831;
  assign n12442 = n5266 | n15832;
  assign n12443 = (n15760 & n12441) | (n15760 & n12442) | (n12441 & n12442);
  assign n5269 = ~n12440 & n12443;
  assign n5270 = x65 & x82;
  assign n5271 = n5269 & n5270;
  assign n5272 = n5269 | n5270;
  assign n5273 = ~n5271 & n5272;
  assign n15833 = n4997 | n5130;
  assign n15834 = (n5130 & n5132) | (n5130 & n15833) | (n5132 & n15833);
  assign n12444 = n5273 & n15834;
  assign n12433 = n5130 | n5132;
  assign n12445 = n5273 & n12433;
  assign n15835 = (n12328 & n12444) | (n12328 & n12445) | (n12444 & n12445);
  assign n15836 = (n12329 & n12444) | (n12329 & n12445) | (n12444 & n12445);
  assign n15837 = (n15726 & n15835) | (n15726 & n15836) | (n15835 & n15836);
  assign n12447 = n5273 | n15834;
  assign n12448 = n5273 | n12433;
  assign n15838 = (n12328 & n12447) | (n12328 & n12448) | (n12447 & n12448);
  assign n15839 = (n12329 & n12447) | (n12329 & n12448) | (n12447 & n12448);
  assign n15840 = (n15726 & n15838) | (n15726 & n15839) | (n15838 & n15839);
  assign n5276 = ~n15837 & n15840;
  assign n5277 = x64 & x83;
  assign n5278 = n5276 & n5277;
  assign n5279 = n5276 | n5277;
  assign n5280 = ~n5278 & n5279;
  assign n12430 = n5137 | n5139;
  assign n12450 = n5280 & n12430;
  assign n12451 = n5137 & n5280;
  assign n15841 = (n12450 & n12451) | (n12450 & n15798) | (n12451 & n15798);
  assign n15842 = (n12450 & n12451) | (n12450 & n15800) | (n12451 & n15800);
  assign n15843 = (n15751 & n15841) | (n15751 & n15842) | (n15841 & n15842);
  assign n12453 = n5280 | n12430;
  assign n12454 = n5137 | n5280;
  assign n15844 = (n12453 & n12454) | (n12453 & n15798) | (n12454 & n15798);
  assign n15845 = (n12453 & n12454) | (n12453 & n15800) | (n12454 & n15800);
  assign n15846 = (n15751 & n15844) | (n15751 & n15845) | (n15844 & n15845);
  assign n5283 = ~n15843 & n15846;
  assign n5284 = x63 & x84;
  assign n5285 = n5283 & n5284;
  assign n5286 = n5283 | n5284;
  assign n5287 = ~n5285 & n5286;
  assign n12428 = n5144 | n5146;
  assign n12456 = n5287 & n12428;
  assign n12457 = n5144 & n5287;
  assign n12458 = (n15796 & n12456) | (n15796 & n12457) | (n12456 & n12457);
  assign n12459 = n5287 | n12428;
  assign n12460 = n5144 | n5287;
  assign n12461 = (n15796 & n12459) | (n15796 & n12460) | (n12459 & n12460);
  assign n5290 = ~n12458 & n12461;
  assign n5291 = x62 & x85;
  assign n5292 = n5290 & n5291;
  assign n5293 = n5290 | n5291;
  assign n5294 = ~n5292 & n5293;
  assign n12462 = n5151 & n5294;
  assign n15847 = (n5294 & n12396) | (n5294 & n12462) | (n12396 & n12462);
  assign n15848 = (n5294 & n12395) | (n5294 & n12462) | (n12395 & n12462);
  assign n15849 = (n15781 & n15847) | (n15781 & n15848) | (n15847 & n15848);
  assign n12464 = n5151 | n5294;
  assign n15850 = n12396 | n12464;
  assign n15851 = n12395 | n12464;
  assign n15852 = (n15781 & n15850) | (n15781 & n15851) | (n15850 & n15851);
  assign n5297 = ~n15849 & n15852;
  assign n5298 = x61 & x86;
  assign n5299 = n5297 & n5298;
  assign n5300 = n5297 | n5298;
  assign n5301 = ~n5299 & n5300;
  assign n5302 = n15829 & n5301;
  assign n5303 = n15829 | n5301;
  assign n5304 = ~n5302 & n5303;
  assign n5305 = x60 & x87;
  assign n5306 = n5304 & n5305;
  assign n5307 = n5304 | n5305;
  assign n5308 = ~n5306 & n5307;
  assign n12466 = n5165 & n5308;
  assign n12467 = (n5308 & n12406) | (n5308 & n12466) | (n12406 & n12466);
  assign n12468 = n5165 | n5308;
  assign n12469 = n12406 | n12468;
  assign n5311 = ~n12467 & n12469;
  assign n5312 = x59 & x88;
  assign n5313 = n5311 & n5312;
  assign n5314 = n5311 | n5312;
  assign n5315 = ~n5313 & n5314;
  assign n12470 = n5172 & n5315;
  assign n12471 = (n5315 & n12410) | (n5315 & n12470) | (n12410 & n12470);
  assign n12472 = n5172 | n5315;
  assign n12473 = n12410 | n12472;
  assign n5318 = ~n12471 & n12473;
  assign n5319 = x58 & x89;
  assign n5320 = n5318 & n5319;
  assign n5321 = n5318 | n5319;
  assign n5322 = ~n5320 & n5321;
  assign n12474 = n5179 & n5322;
  assign n12475 = (n5322 & n12414) | (n5322 & n12474) | (n12414 & n12474);
  assign n12476 = n5179 | n5322;
  assign n12477 = n12414 | n12476;
  assign n5325 = ~n12475 & n12477;
  assign n5326 = x57 & x90;
  assign n5327 = n5325 & n5326;
  assign n5328 = n5325 | n5326;
  assign n5329 = ~n5327 & n5328;
  assign n5330 = n12424 & n5329;
  assign n5331 = n12424 | n5329;
  assign n5332 = ~n5330 & n5331;
  assign n5333 = x56 & x91;
  assign n5334 = n5332 & n5333;
  assign n5335 = n5332 | n5333;
  assign n5336 = ~n5334 & n5335;
  assign n5337 = n12422 & n5336;
  assign n5338 = n12422 | n5336;
  assign n5339 = ~n5337 & n5338;
  assign n5340 = x55 & x92;
  assign n5341 = n5339 & n5340;
  assign n5342 = n5339 | n5340;
  assign n5343 = ~n5341 & n5342;
  assign n5344 = n12420 & n5343;
  assign n5345 = n12420 | n5343;
  assign n5346 = ~n5344 & n5345;
  assign n5347 = x54 & x93;
  assign n5348 = n5346 & n5347;
  assign n5349 = n5346 | n5347;
  assign n5350 = ~n5348 & n5349;
  assign n5351 = n5249 & n5350;
  assign n5352 = n5249 | n5350;
  assign n5353 = ~n5351 & n5352;
  assign n5354 = x53 & x94;
  assign n5355 = n5353 & n5354;
  assign n5356 = n5353 | n5354;
  assign n5357 = ~n5355 & n5356;
  assign n5358 = n5248 & n5357;
  assign n5359 = n5248 | n5357;
  assign n5360 = ~n5358 & n5359;
  assign n5361 = x52 & x95;
  assign n5362 = n5360 & n5361;
  assign n5363 = n5360 | n5361;
  assign n5364 = ~n5362 & n5363;
  assign n5365 = n5247 & n5364;
  assign n5366 = n5247 | n5364;
  assign n5367 = ~n5365 & n5366;
  assign n5368 = x51 & x96;
  assign n5369 = n5367 & n5368;
  assign n5370 = n5367 | n5368;
  assign n5371 = ~n5369 & n5370;
  assign n5372 = n15824 & n5371;
  assign n5373 = n15824 | n5371;
  assign n5374 = ~n5372 & n5373;
  assign n5375 = x50 & x97;
  assign n5376 = n5374 & n5375;
  assign n5377 = n5374 | n5375;
  assign n5378 = ~n5376 & n5377;
  assign n5379 = n12418 & n5378;
  assign n5380 = n12418 | n5378;
  assign n5381 = ~n5379 & n5380;
  assign n5382 = x49 & x98;
  assign n5383 = n5381 & n5382;
  assign n5384 = n5381 | n5382;
  assign n5385 = ~n5383 & n5384;
  assign n5386 = n5242 & n5385;
  assign n5387 = n5242 | n5385;
  assign n5388 = ~n5386 & n5387;
  assign n5389 = x48 & x99;
  assign n5390 = n5388 & n5389;
  assign n5391 = n5388 | n5389;
  assign n5392 = ~n5390 & n5391;
  assign n49880 = n5241 | n5382;
  assign n49881 = (n5240 & n5382) | (n5240 & n49880) | (n5382 & n49880);
  assign n15854 = (n5242 & n5381) | (n5242 & n49881) | (n5381 & n49881);
  assign n12479 = (n5383 & n5385) | (n5383 & n15854) | (n5385 & n15854);
  assign n12480 = n5376 | n12418;
  assign n12481 = (n5376 & n5378) | (n5376 & n12480) | (n5378 & n12480);
  assign n15855 = n5369 | n15824;
  assign n15856 = (n5369 & n5371) | (n5369 & n15855) | (n5371 & n15855);
  assign n5396 = n5362 | n5365;
  assign n5397 = n5355 | n5358;
  assign n12482 = n5348 | n5350;
  assign n12483 = (n5249 & n5348) | (n5249 & n12482) | (n5348 & n12482);
  assign n12484 = n5341 | n5343;
  assign n12485 = (n5341 & n12420) | (n5341 & n12484) | (n12420 & n12484);
  assign n12486 = n5334 | n5336;
  assign n12487 = (n5334 & n12422) | (n5334 & n12486) | (n12422 & n12486);
  assign n12488 = n5327 | n5329;
  assign n12489 = (n5327 & n12424) | (n5327 & n12488) | (n12424 & n12488);
  assign n12493 = n5292 | n5294;
  assign n15857 = n5151 | n5292;
  assign n15858 = (n5292 & n5294) | (n5292 & n15857) | (n5294 & n15857);
  assign n15859 = (n12396 & n12493) | (n12396 & n15858) | (n12493 & n15858);
  assign n15860 = (n12395 & n12493) | (n12395 & n15858) | (n12493 & n15858);
  assign n15861 = (n15781 & n15859) | (n15781 & n15860) | (n15859 & n15860);
  assign n15862 = n5278 | n5280;
  assign n15863 = (n5278 & n12430) | (n5278 & n15862) | (n12430 & n15862);
  assign n15864 = n5137 | n5278;
  assign n15865 = (n5278 & n5280) | (n5278 & n15864) | (n5280 & n15864);
  assign n15866 = (n15798 & n15863) | (n15798 & n15865) | (n15863 & n15865);
  assign n15867 = (n15800 & n15863) | (n15800 & n15865) | (n15863 & n15865);
  assign n15868 = (n15751 & n15866) | (n15751 & n15867) | (n15866 & n15867);
  assign n15869 = n5271 | n5273;
  assign n15870 = (n5271 & n15834) | (n5271 & n15869) | (n15834 & n15869);
  assign n15871 = (n5271 & n12433) | (n5271 & n15869) | (n12433 & n15869);
  assign n15872 = (n12328 & n15870) | (n12328 & n15871) | (n15870 & n15871);
  assign n15873 = (n12329 & n15870) | (n12329 & n15871) | (n15870 & n15871);
  assign n15874 = (n15726 & n15872) | (n15726 & n15873) | (n15872 & n15873);
  assign n5411 = x68 & x80;
  assign n5412 = x67 & x81;
  assign n5413 = n5411 & n5412;
  assign n5414 = n5411 | n5412;
  assign n5415 = ~n5413 & n5414;
  assign n15875 = n5264 | n5266;
  assign n15877 = n5415 & n15875;
  assign n15878 = n5264 & n5415;
  assign n15879 = (n15831 & n15877) | (n15831 & n15878) | (n15877 & n15878);
  assign n15881 = (n15832 & n15877) | (n15832 & n15878) | (n15877 & n15878);
  assign n12506 = (n15760 & n15879) | (n15760 & n15881) | (n15879 & n15881);
  assign n15882 = n5415 | n15875;
  assign n15883 = n5264 | n5415;
  assign n15884 = (n15831 & n15882) | (n15831 & n15883) | (n15882 & n15883);
  assign n15885 = (n15832 & n15882) | (n15832 & n15883) | (n15882 & n15883);
  assign n12509 = (n15760 & n15884) | (n15760 & n15885) | (n15884 & n15885);
  assign n5418 = ~n12506 & n12509;
  assign n5419 = x66 & x82;
  assign n5420 = n5418 & n5419;
  assign n5421 = n5418 | n5419;
  assign n5422 = ~n5420 & n5421;
  assign n5423 = n15874 & n5422;
  assign n5424 = n15874 | n5422;
  assign n5425 = ~n5423 & n5424;
  assign n5426 = x65 & x83;
  assign n5427 = n5425 & n5426;
  assign n5428 = n5425 | n5426;
  assign n5429 = ~n5427 & n5428;
  assign n5430 = n15868 & n5429;
  assign n5431 = n15868 | n5429;
  assign n5432 = ~n5430 & n5431;
  assign n5433 = x64 & x84;
  assign n5434 = n5432 & n5433;
  assign n5435 = n5432 | n5433;
  assign n5436 = ~n5434 & n5435;
  assign n12510 = n5285 & n5436;
  assign n15886 = (n5436 & n12456) | (n5436 & n12510) | (n12456 & n12510);
  assign n15887 = (n5436 & n12457) | (n5436 & n12510) | (n12457 & n12510);
  assign n15888 = (n15796 & n15886) | (n15796 & n15887) | (n15886 & n15887);
  assign n12512 = n5285 | n5436;
  assign n15889 = n12456 | n12512;
  assign n15890 = n12457 | n12512;
  assign n15891 = (n15796 & n15889) | (n15796 & n15890) | (n15889 & n15890);
  assign n5439 = ~n15888 & n15891;
  assign n5440 = x63 & x85;
  assign n5441 = n5439 & n5440;
  assign n5442 = n5439 | n5440;
  assign n5443 = ~n5441 & n5442;
  assign n5444 = n15861 & n5443;
  assign n5445 = n15861 | n5443;
  assign n5446 = ~n5444 & n5445;
  assign n5447 = x62 & x86;
  assign n5448 = n5446 & n5447;
  assign n5449 = n5446 | n5447;
  assign n5450 = ~n5448 & n5449;
  assign n12490 = n5299 | n5301;
  assign n12514 = n5450 & n12490;
  assign n12515 = n5299 & n5450;
  assign n12516 = (n15829 & n12514) | (n15829 & n12515) | (n12514 & n12515);
  assign n12517 = n5450 | n12490;
  assign n12518 = n5299 | n5450;
  assign n12519 = (n15829 & n12517) | (n15829 & n12518) | (n12517 & n12518);
  assign n5453 = ~n12516 & n12519;
  assign n5454 = x61 & x87;
  assign n5455 = n5453 & n5454;
  assign n5456 = n5453 | n5454;
  assign n5457 = ~n5455 & n5456;
  assign n12520 = n5306 & n5457;
  assign n15892 = (n5457 & n12466) | (n5457 & n12520) | (n12466 & n12520);
  assign n15893 = (n5308 & n5457) | (n5308 & n12520) | (n5457 & n12520);
  assign n15894 = (n12406 & n15892) | (n12406 & n15893) | (n15892 & n15893);
  assign n12522 = n5306 | n5457;
  assign n15895 = n12466 | n12522;
  assign n15896 = n5308 | n12522;
  assign n15897 = (n12406 & n15895) | (n12406 & n15896) | (n15895 & n15896);
  assign n5460 = ~n15894 & n15897;
  assign n5461 = x60 & x88;
  assign n5462 = n5460 & n5461;
  assign n5463 = n5460 | n5461;
  assign n5464 = ~n5462 & n5463;
  assign n12524 = n5313 & n5464;
  assign n12525 = (n5464 & n12471) | (n5464 & n12524) | (n12471 & n12524);
  assign n12526 = n5313 | n5464;
  assign n12527 = n12471 | n12526;
  assign n5467 = ~n12525 & n12527;
  assign n5468 = x59 & x89;
  assign n5469 = n5467 & n5468;
  assign n5470 = n5467 | n5468;
  assign n5471 = ~n5469 & n5470;
  assign n12528 = n5320 & n5471;
  assign n12529 = (n5471 & n12475) | (n5471 & n12528) | (n12475 & n12528);
  assign n12530 = n5320 | n5471;
  assign n12531 = n12475 | n12530;
  assign n5474 = ~n12529 & n12531;
  assign n5475 = x58 & x90;
  assign n5476 = n5474 & n5475;
  assign n5477 = n5474 | n5475;
  assign n5478 = ~n5476 & n5477;
  assign n5479 = n12489 & n5478;
  assign n5480 = n12489 | n5478;
  assign n5481 = ~n5479 & n5480;
  assign n5482 = x57 & x91;
  assign n5483 = n5481 & n5482;
  assign n5484 = n5481 | n5482;
  assign n5485 = ~n5483 & n5484;
  assign n5486 = n12487 & n5485;
  assign n5487 = n12487 | n5485;
  assign n5488 = ~n5486 & n5487;
  assign n5489 = x56 & x92;
  assign n5490 = n5488 & n5489;
  assign n5491 = n5488 | n5489;
  assign n5492 = ~n5490 & n5491;
  assign n5493 = n12485 & n5492;
  assign n5494 = n12485 | n5492;
  assign n5495 = ~n5493 & n5494;
  assign n5496 = x55 & x93;
  assign n5497 = n5495 & n5496;
  assign n5498 = n5495 | n5496;
  assign n5499 = ~n5497 & n5498;
  assign n5500 = n12483 & n5499;
  assign n5501 = n12483 | n5499;
  assign n5502 = ~n5500 & n5501;
  assign n5503 = x54 & x94;
  assign n5504 = n5502 & n5503;
  assign n5505 = n5502 | n5503;
  assign n5506 = ~n5504 & n5505;
  assign n5507 = n5397 & n5506;
  assign n5508 = n5397 | n5506;
  assign n5509 = ~n5507 & n5508;
  assign n5510 = x53 & x95;
  assign n5511 = n5509 & n5510;
  assign n5512 = n5509 | n5510;
  assign n5513 = ~n5511 & n5512;
  assign n5514 = n5396 & n5513;
  assign n5515 = n5396 | n5513;
  assign n5516 = ~n5514 & n5515;
  assign n5517 = x52 & x96;
  assign n5518 = n5516 & n5517;
  assign n5519 = n5516 | n5517;
  assign n5520 = ~n5518 & n5519;
  assign n5521 = n15856 & n5520;
  assign n5522 = n15856 | n5520;
  assign n5523 = ~n5521 & n5522;
  assign n5524 = x51 & x97;
  assign n5525 = n5523 & n5524;
  assign n5526 = n5523 | n5524;
  assign n5527 = ~n5525 & n5526;
  assign n5528 = n12481 & n5527;
  assign n5529 = n12481 | n5527;
  assign n5530 = ~n5528 & n5529;
  assign n5531 = x50 & x98;
  assign n5532 = n5530 & n5531;
  assign n5533 = n5530 | n5531;
  assign n5534 = ~n5532 & n5533;
  assign n5535 = n12479 & n5534;
  assign n5536 = n12479 | n5534;
  assign n5537 = ~n5535 & n5536;
  assign n5538 = x49 & x99;
  assign n5539 = n5537 & n5538;
  assign n5540 = n5537 | n5538;
  assign n5541 = ~n5539 & n5540;
  assign n5542 = n5390 & n5541;
  assign n5543 = n5390 | n5541;
  assign n5544 = ~n5542 & n5543;
  assign n5545 = x48 & x100;
  assign n5546 = n5544 & n5545;
  assign n5547 = n5544 | n5545;
  assign n5548 = ~n5546 & n5547;
  assign n49882 = n5389 | n5538;
  assign n49883 = (n5388 & n5538) | (n5388 & n49882) | (n5538 & n49882);
  assign n15899 = (n5390 & n5537) | (n5390 & n49883) | (n5537 & n49883);
  assign n12533 = (n5539 & n5541) | (n5539 & n15899) | (n5541 & n15899);
  assign n12534 = n5532 | n12479;
  assign n12535 = (n5532 & n5534) | (n5532 & n12534) | (n5534 & n12534);
  assign n12536 = n5525 | n12481;
  assign n12537 = (n5525 & n5527) | (n5525 & n12536) | (n5527 & n12536);
  assign n15900 = n5518 | n15856;
  assign n15901 = (n5518 & n5520) | (n5518 & n15900) | (n5520 & n15900);
  assign n5553 = n5511 | n5514;
  assign n12538 = n5504 | n5506;
  assign n12539 = (n5397 & n5504) | (n5397 & n12538) | (n5504 & n12538);
  assign n12540 = n5497 | n5499;
  assign n12541 = (n5497 & n12483) | (n5497 & n12540) | (n12483 & n12540);
  assign n12542 = n5490 | n5492;
  assign n12543 = (n5490 & n12485) | (n5490 & n12542) | (n12485 & n12542);
  assign n12544 = n5483 | n5485;
  assign n12545 = (n5483 & n12487) | (n5483 & n12544) | (n12487 & n12544);
  assign n12546 = n5476 | n5478;
  assign n12547 = (n5476 & n12489) | (n5476 & n12546) | (n12489 & n12546);
  assign n12549 = n5455 | n5457;
  assign n15902 = n5306 | n5455;
  assign n15903 = (n5455 & n5457) | (n5455 & n15902) | (n5457 & n15902);
  assign n15904 = (n12466 & n12549) | (n12466 & n15903) | (n12549 & n15903);
  assign n15905 = (n5308 & n12549) | (n5308 & n15903) | (n12549 & n15903);
  assign n15906 = (n12406 & n15904) | (n12406 & n15905) | (n15904 & n15905);
  assign n12554 = n5434 | n5436;
  assign n15907 = n5285 | n5434;
  assign n15908 = (n5434 & n5436) | (n5434 & n15907) | (n5436 & n15907);
  assign n15909 = (n12456 & n12554) | (n12456 & n15908) | (n12554 & n15908);
  assign n15910 = (n12457 & n12554) | (n12457 & n15908) | (n12554 & n15908);
  assign n15911 = (n15796 & n15909) | (n15796 & n15910) | (n15909 & n15910);
  assign n5568 = x69 & x80;
  assign n5569 = x68 & x81;
  assign n5570 = n5568 & n5569;
  assign n5571 = n5568 | n5569;
  assign n5572 = ~n5570 & n5571;
  assign n12560 = n5413 & n5572;
  assign n15912 = (n5572 & n12560) | (n5572 & n15881) | (n12560 & n15881);
  assign n15913 = (n5572 & n12560) | (n5572 & n15879) | (n12560 & n15879);
  assign n15914 = (n15760 & n15912) | (n15760 & n15913) | (n15912 & n15913);
  assign n12562 = n5413 | n5572;
  assign n15915 = n12562 | n15881;
  assign n15916 = n12562 | n15879;
  assign n15917 = (n15760 & n15915) | (n15760 & n15916) | (n15915 & n15916);
  assign n5575 = ~n15914 & n15917;
  assign n5576 = x67 & x82;
  assign n5577 = n5575 & n5576;
  assign n5578 = n5575 | n5576;
  assign n5579 = ~n5577 & n5578;
  assign n12558 = n5420 | n5422;
  assign n12564 = n5579 & n12558;
  assign n12565 = n5420 & n5579;
  assign n12566 = (n15874 & n12564) | (n15874 & n12565) | (n12564 & n12565);
  assign n12567 = n5579 | n12558;
  assign n12568 = n5420 | n5579;
  assign n12569 = (n15874 & n12567) | (n15874 & n12568) | (n12567 & n12568);
  assign n5582 = ~n12566 & n12569;
  assign n5583 = x66 & x83;
  assign n5584 = n5582 & n5583;
  assign n5585 = n5582 | n5583;
  assign n5586 = ~n5584 & n5585;
  assign n12556 = n5427 | n5429;
  assign n12570 = n5586 & n12556;
  assign n12571 = n5427 & n5586;
  assign n12572 = (n15868 & n12570) | (n15868 & n12571) | (n12570 & n12571);
  assign n12573 = n5586 | n12556;
  assign n12574 = n5427 | n5586;
  assign n12575 = (n15868 & n12573) | (n15868 & n12574) | (n12573 & n12574);
  assign n5589 = ~n12572 & n12575;
  assign n5590 = x65 & x84;
  assign n5591 = n5589 & n5590;
  assign n5592 = n5589 | n5590;
  assign n5593 = ~n5591 & n5592;
  assign n5594 = n15911 & n5593;
  assign n5595 = n15911 | n5593;
  assign n5596 = ~n5594 & n5595;
  assign n5597 = x64 & x85;
  assign n5598 = n5596 & n5597;
  assign n5599 = n5596 | n5597;
  assign n5600 = ~n5598 & n5599;
  assign n12551 = n5441 | n5443;
  assign n12576 = n5600 & n12551;
  assign n12577 = n5441 & n5600;
  assign n12578 = (n15861 & n12576) | (n15861 & n12577) | (n12576 & n12577);
  assign n12579 = n5600 | n12551;
  assign n12580 = n5441 | n5600;
  assign n12581 = (n15861 & n12579) | (n15861 & n12580) | (n12579 & n12580);
  assign n5603 = ~n12578 & n12581;
  assign n5604 = x63 & x86;
  assign n5605 = n5603 & n5604;
  assign n5606 = n5603 | n5604;
  assign n5607 = ~n5605 & n5606;
  assign n12582 = n5448 & n5607;
  assign n15918 = (n5607 & n12515) | (n5607 & n12582) | (n12515 & n12582);
  assign n15919 = (n5607 & n12514) | (n5607 & n12582) | (n12514 & n12582);
  assign n15920 = (n15829 & n15918) | (n15829 & n15919) | (n15918 & n15919);
  assign n12584 = n5448 | n5607;
  assign n15921 = n12515 | n12584;
  assign n15922 = n12514 | n12584;
  assign n15923 = (n15829 & n15921) | (n15829 & n15922) | (n15921 & n15922);
  assign n5610 = ~n15920 & n15923;
  assign n5611 = x62 & x87;
  assign n5612 = n5610 & n5611;
  assign n5613 = n5610 | n5611;
  assign n5614 = ~n5612 & n5613;
  assign n5615 = n15906 & n5614;
  assign n5616 = n15906 | n5614;
  assign n5617 = ~n5615 & n5616;
  assign n5618 = x61 & x88;
  assign n5619 = n5617 & n5618;
  assign n5620 = n5617 | n5618;
  assign n5621 = ~n5619 & n5620;
  assign n12586 = n5462 & n5621;
  assign n12587 = (n5621 & n12525) | (n5621 & n12586) | (n12525 & n12586);
  assign n12588 = n5462 | n5621;
  assign n12589 = n12525 | n12588;
  assign n5624 = ~n12587 & n12589;
  assign n5625 = x60 & x89;
  assign n5626 = n5624 & n5625;
  assign n5627 = n5624 | n5625;
  assign n5628 = ~n5626 & n5627;
  assign n12590 = n5469 & n5628;
  assign n12591 = (n5628 & n12529) | (n5628 & n12590) | (n12529 & n12590);
  assign n12592 = n5469 | n5628;
  assign n12593 = n12529 | n12592;
  assign n5631 = ~n12591 & n12593;
  assign n5632 = x59 & x90;
  assign n5633 = n5631 & n5632;
  assign n5634 = n5631 | n5632;
  assign n5635 = ~n5633 & n5634;
  assign n5636 = n12547 & n5635;
  assign n5637 = n12547 | n5635;
  assign n5638 = ~n5636 & n5637;
  assign n5639 = x58 & x91;
  assign n5640 = n5638 & n5639;
  assign n5641 = n5638 | n5639;
  assign n5642 = ~n5640 & n5641;
  assign n5643 = n12545 & n5642;
  assign n5644 = n12545 | n5642;
  assign n5645 = ~n5643 & n5644;
  assign n5646 = x57 & x92;
  assign n5647 = n5645 & n5646;
  assign n5648 = n5645 | n5646;
  assign n5649 = ~n5647 & n5648;
  assign n5650 = n12543 & n5649;
  assign n5651 = n12543 | n5649;
  assign n5652 = ~n5650 & n5651;
  assign n5653 = x56 & x93;
  assign n5654 = n5652 & n5653;
  assign n5655 = n5652 | n5653;
  assign n5656 = ~n5654 & n5655;
  assign n5657 = n12541 & n5656;
  assign n5658 = n12541 | n5656;
  assign n5659 = ~n5657 & n5658;
  assign n5660 = x55 & x94;
  assign n5661 = n5659 & n5660;
  assign n5662 = n5659 | n5660;
  assign n5663 = ~n5661 & n5662;
  assign n5664 = n12539 & n5663;
  assign n5665 = n12539 | n5663;
  assign n5666 = ~n5664 & n5665;
  assign n5667 = x54 & x95;
  assign n5668 = n5666 & n5667;
  assign n5669 = n5666 | n5667;
  assign n5670 = ~n5668 & n5669;
  assign n5671 = n5553 & n5670;
  assign n5672 = n5553 | n5670;
  assign n5673 = ~n5671 & n5672;
  assign n5674 = x53 & x96;
  assign n5675 = n5673 & n5674;
  assign n5676 = n5673 | n5674;
  assign n5677 = ~n5675 & n5676;
  assign n5678 = n15901 & n5677;
  assign n5679 = n15901 | n5677;
  assign n5680 = ~n5678 & n5679;
  assign n5681 = x52 & x97;
  assign n5682 = n5680 & n5681;
  assign n5683 = n5680 | n5681;
  assign n5684 = ~n5682 & n5683;
  assign n5685 = n12537 & n5684;
  assign n5686 = n12537 | n5684;
  assign n5687 = ~n5685 & n5686;
  assign n5688 = x51 & x98;
  assign n5689 = n5687 & n5688;
  assign n5690 = n5687 | n5688;
  assign n5691 = ~n5689 & n5690;
  assign n5692 = n12535 & n5691;
  assign n5693 = n12535 | n5691;
  assign n5694 = ~n5692 & n5693;
  assign n5695 = x50 & x99;
  assign n5696 = n5694 & n5695;
  assign n5697 = n5694 | n5695;
  assign n5698 = ~n5696 & n5697;
  assign n5699 = n12533 & n5698;
  assign n5700 = n12533 | n5698;
  assign n5701 = ~n5699 & n5700;
  assign n5702 = x49 & x100;
  assign n5703 = n5701 & n5702;
  assign n5704 = n5701 | n5702;
  assign n5705 = ~n5703 & n5704;
  assign n5706 = n5546 & n5705;
  assign n5707 = n5546 | n5705;
  assign n5708 = ~n5706 & n5707;
  assign n5709 = x48 & x101;
  assign n5710 = n5708 & n5709;
  assign n5711 = n5708 | n5709;
  assign n5712 = ~n5710 & n5711;
  assign n49884 = n5545 | n5702;
  assign n49885 = (n5544 & n5702) | (n5544 & n49884) | (n5702 & n49884);
  assign n15925 = (n5546 & n5701) | (n5546 & n49885) | (n5701 & n49885);
  assign n12595 = (n5703 & n5705) | (n5703 & n15925) | (n5705 & n15925);
  assign n12596 = n5696 | n12533;
  assign n12597 = (n5696 & n5698) | (n5696 & n12596) | (n5698 & n12596);
  assign n12598 = n5689 | n12535;
  assign n12599 = (n5689 & n5691) | (n5689 & n12598) | (n5691 & n12598);
  assign n12600 = n5682 | n12537;
  assign n12601 = (n5682 & n5684) | (n5682 & n12600) | (n5684 & n12600);
  assign n15926 = n5675 | n15901;
  assign n15927 = (n5675 & n5677) | (n5675 & n15926) | (n5677 & n15926);
  assign n12602 = n5668 | n5670;
  assign n12603 = (n5553 & n5668) | (n5553 & n12602) | (n5668 & n12602);
  assign n12604 = n5661 | n5663;
  assign n12605 = (n5661 & n12539) | (n5661 & n12604) | (n12539 & n12604);
  assign n12606 = n5654 | n5656;
  assign n12607 = (n5654 & n12541) | (n5654 & n12606) | (n12541 & n12606);
  assign n12608 = n5647 | n5649;
  assign n12609 = (n5647 & n12543) | (n5647 & n12608) | (n12543 & n12608);
  assign n12610 = n5640 | n5642;
  assign n12611 = (n5640 & n12545) | (n5640 & n12610) | (n12545 & n12610);
  assign n12612 = n5633 | n5635;
  assign n12613 = (n5633 & n12547) | (n5633 & n12612) | (n12547 & n12612);
  assign n12617 = n5605 | n5607;
  assign n15928 = n5448 | n5605;
  assign n15929 = (n5605 & n5607) | (n5605 & n15928) | (n5607 & n15928);
  assign n15930 = (n12515 & n12617) | (n12515 & n15929) | (n12617 & n15929);
  assign n15931 = (n12514 & n12617) | (n12514 & n15929) | (n12617 & n15929);
  assign n15932 = (n15829 & n15930) | (n15829 & n15931) | (n15930 & n15931);
  assign n5733 = x70 & x80;
  assign n5734 = x69 & x81;
  assign n5735 = n5733 & n5734;
  assign n5736 = n5733 | n5734;
  assign n5737 = ~n5735 & n5736;
  assign n15937 = n5413 | n5570;
  assign n15938 = (n5570 & n5572) | (n5570 & n15937) | (n5572 & n15937);
  assign n12630 = n5737 & n15938;
  assign n12628 = n5570 | n5572;
  assign n12631 = n5737 & n12628;
  assign n15939 = (n12630 & n12631) | (n12630 & n15881) | (n12631 & n15881);
  assign n15940 = (n12630 & n12631) | (n12630 & n15879) | (n12631 & n15879);
  assign n15941 = (n15760 & n15939) | (n15760 & n15940) | (n15939 & n15940);
  assign n12633 = n5737 | n15938;
  assign n12634 = n5737 | n12628;
  assign n15942 = (n12633 & n12634) | (n12633 & n15881) | (n12634 & n15881);
  assign n15943 = (n12633 & n12634) | (n12633 & n15879) | (n12634 & n15879);
  assign n15944 = (n15760 & n15942) | (n15760 & n15943) | (n15942 & n15943);
  assign n5740 = ~n15941 & n15944;
  assign n5741 = x68 & x82;
  assign n5742 = n5740 & n5741;
  assign n5743 = n5740 | n5741;
  assign n5744 = ~n5742 & n5743;
  assign n15945 = n5577 | n5579;
  assign n15946 = (n5577 & n12558) | (n5577 & n15945) | (n12558 & n15945);
  assign n12636 = n5744 & n15946;
  assign n15947 = n5420 | n5577;
  assign n15948 = (n5577 & n5579) | (n5577 & n15947) | (n5579 & n15947);
  assign n12637 = n5744 & n15948;
  assign n12638 = (n15874 & n12636) | (n15874 & n12637) | (n12636 & n12637);
  assign n12639 = n5744 | n15946;
  assign n12640 = n5744 | n15948;
  assign n12641 = (n15874 & n12639) | (n15874 & n12640) | (n12639 & n12640);
  assign n5747 = ~n12638 & n12641;
  assign n5748 = x67 & x83;
  assign n5749 = n5747 & n5748;
  assign n5750 = n5747 | n5748;
  assign n5751 = ~n5749 & n5750;
  assign n15933 = n5584 | n5586;
  assign n15934 = (n5584 & n12556) | (n5584 & n15933) | (n12556 & n15933);
  assign n15949 = n5751 & n15934;
  assign n15935 = n5427 | n5584;
  assign n15936 = (n5584 & n5586) | (n5584 & n15935) | (n5586 & n15935);
  assign n15950 = n5751 & n15936;
  assign n15951 = (n15868 & n15949) | (n15868 & n15950) | (n15949 & n15950);
  assign n15952 = n5751 | n15934;
  assign n15953 = n5751 | n15936;
  assign n15954 = (n15868 & n15952) | (n15868 & n15953) | (n15952 & n15953);
  assign n5754 = ~n15951 & n15954;
  assign n5755 = x66 & x84;
  assign n5756 = n5754 & n5755;
  assign n5757 = n5754 | n5755;
  assign n5758 = ~n5756 & n5757;
  assign n12619 = n5591 | n5593;
  assign n12642 = n5758 & n12619;
  assign n12643 = n5591 & n5758;
  assign n12644 = (n15911 & n12642) | (n15911 & n12643) | (n12642 & n12643);
  assign n12645 = n5758 | n12619;
  assign n12646 = n5591 | n5758;
  assign n12647 = (n15911 & n12645) | (n15911 & n12646) | (n12645 & n12646);
  assign n5761 = ~n12644 & n12647;
  assign n5762 = x65 & x85;
  assign n5763 = n5761 & n5762;
  assign n5764 = n5761 | n5762;
  assign n5765 = ~n5763 & n5764;
  assign n12648 = n5598 & n5765;
  assign n15955 = (n5765 & n12577) | (n5765 & n12648) | (n12577 & n12648);
  assign n15956 = (n5765 & n12576) | (n5765 & n12648) | (n12576 & n12648);
  assign n15957 = (n15861 & n15955) | (n15861 & n15956) | (n15955 & n15956);
  assign n12650 = n5598 | n5765;
  assign n15958 = n12577 | n12650;
  assign n15959 = n12576 | n12650;
  assign n15960 = (n15861 & n15958) | (n15861 & n15959) | (n15958 & n15959);
  assign n5768 = ~n15957 & n15960;
  assign n5769 = x64 & x86;
  assign n5770 = n5768 & n5769;
  assign n5771 = n5768 | n5769;
  assign n5772 = ~n5770 & n5771;
  assign n5773 = n15932 & n5772;
  assign n5774 = n15932 | n5772;
  assign n5775 = ~n5773 & n5774;
  assign n5776 = x63 & x87;
  assign n5777 = n5775 & n5776;
  assign n5778 = n5775 | n5776;
  assign n5779 = ~n5777 & n5778;
  assign n12614 = n5612 | n5614;
  assign n12652 = n5779 & n12614;
  assign n12653 = n5612 & n5779;
  assign n12654 = (n15906 & n12652) | (n15906 & n12653) | (n12652 & n12653);
  assign n12655 = n5779 | n12614;
  assign n12656 = n5612 | n5779;
  assign n12657 = (n15906 & n12655) | (n15906 & n12656) | (n12655 & n12656);
  assign n5782 = ~n12654 & n12657;
  assign n5783 = x62 & x88;
  assign n5784 = n5782 & n5783;
  assign n5785 = n5782 | n5783;
  assign n5786 = ~n5784 & n5785;
  assign n12658 = n5619 & n5786;
  assign n15961 = (n5786 & n12586) | (n5786 & n12658) | (n12586 & n12658);
  assign n15962 = (n5621 & n5786) | (n5621 & n12658) | (n5786 & n12658);
  assign n15963 = (n12525 & n15961) | (n12525 & n15962) | (n15961 & n15962);
  assign n12660 = n5619 | n5786;
  assign n15964 = n12586 | n12660;
  assign n15965 = n5621 | n12660;
  assign n15966 = (n12525 & n15964) | (n12525 & n15965) | (n15964 & n15965);
  assign n5789 = ~n15963 & n15966;
  assign n5790 = x61 & x89;
  assign n5791 = n5789 & n5790;
  assign n5792 = n5789 | n5790;
  assign n5793 = ~n5791 & n5792;
  assign n12662 = n5626 & n5793;
  assign n12663 = (n5793 & n12591) | (n5793 & n12662) | (n12591 & n12662);
  assign n12664 = n5626 | n5793;
  assign n12665 = n12591 | n12664;
  assign n5796 = ~n12663 & n12665;
  assign n5797 = x60 & x90;
  assign n5798 = n5796 & n5797;
  assign n5799 = n5796 | n5797;
  assign n5800 = ~n5798 & n5799;
  assign n5801 = n12613 & n5800;
  assign n5802 = n12613 | n5800;
  assign n5803 = ~n5801 & n5802;
  assign n5804 = x59 & x91;
  assign n5805 = n5803 & n5804;
  assign n5806 = n5803 | n5804;
  assign n5807 = ~n5805 & n5806;
  assign n5808 = n12611 & n5807;
  assign n5809 = n12611 | n5807;
  assign n5810 = ~n5808 & n5809;
  assign n5811 = x58 & x92;
  assign n5812 = n5810 & n5811;
  assign n5813 = n5810 | n5811;
  assign n5814 = ~n5812 & n5813;
  assign n5815 = n12609 & n5814;
  assign n5816 = n12609 | n5814;
  assign n5817 = ~n5815 & n5816;
  assign n5818 = x57 & x93;
  assign n5819 = n5817 & n5818;
  assign n5820 = n5817 | n5818;
  assign n5821 = ~n5819 & n5820;
  assign n5822 = n12607 & n5821;
  assign n5823 = n12607 | n5821;
  assign n5824 = ~n5822 & n5823;
  assign n5825 = x56 & x94;
  assign n5826 = n5824 & n5825;
  assign n5827 = n5824 | n5825;
  assign n5828 = ~n5826 & n5827;
  assign n5829 = n12605 & n5828;
  assign n5830 = n12605 | n5828;
  assign n5831 = ~n5829 & n5830;
  assign n5832 = x55 & x95;
  assign n5833 = n5831 & n5832;
  assign n5834 = n5831 | n5832;
  assign n5835 = ~n5833 & n5834;
  assign n5836 = n12603 & n5835;
  assign n5837 = n12603 | n5835;
  assign n5838 = ~n5836 & n5837;
  assign n5839 = x54 & x96;
  assign n5840 = n5838 & n5839;
  assign n5841 = n5838 | n5839;
  assign n5842 = ~n5840 & n5841;
  assign n5843 = n15927 & n5842;
  assign n5844 = n15927 | n5842;
  assign n5845 = ~n5843 & n5844;
  assign n5846 = x53 & x97;
  assign n5847 = n5845 & n5846;
  assign n5848 = n5845 | n5846;
  assign n5849 = ~n5847 & n5848;
  assign n5850 = n12601 & n5849;
  assign n5851 = n12601 | n5849;
  assign n5852 = ~n5850 & n5851;
  assign n5853 = x52 & x98;
  assign n5854 = n5852 & n5853;
  assign n5855 = n5852 | n5853;
  assign n5856 = ~n5854 & n5855;
  assign n5857 = n12599 & n5856;
  assign n5858 = n12599 | n5856;
  assign n5859 = ~n5857 & n5858;
  assign n5860 = x51 & x99;
  assign n5861 = n5859 & n5860;
  assign n5862 = n5859 | n5860;
  assign n5863 = ~n5861 & n5862;
  assign n5864 = n12597 & n5863;
  assign n5865 = n12597 | n5863;
  assign n5866 = ~n5864 & n5865;
  assign n5867 = x50 & x100;
  assign n5868 = n5866 & n5867;
  assign n5869 = n5866 | n5867;
  assign n5870 = ~n5868 & n5869;
  assign n5871 = n12595 & n5870;
  assign n5872 = n12595 | n5870;
  assign n5873 = ~n5871 & n5872;
  assign n5874 = x49 & x101;
  assign n5875 = n5873 & n5874;
  assign n5876 = n5873 | n5874;
  assign n5877 = ~n5875 & n5876;
  assign n5878 = n5710 & n5877;
  assign n5879 = n5710 | n5877;
  assign n5880 = ~n5878 & n5879;
  assign n5881 = x48 & x102;
  assign n5882 = n5880 & n5881;
  assign n5883 = n5880 | n5881;
  assign n5884 = ~n5882 & n5883;
  assign n12666 = n5710 | n5875;
  assign n12667 = (n5875 & n5877) | (n5875 & n12666) | (n5877 & n12666);
  assign n12668 = n5868 | n12595;
  assign n12669 = (n5868 & n5870) | (n5868 & n12668) | (n5870 & n12668);
  assign n12670 = n5861 | n12597;
  assign n12671 = (n5861 & n5863) | (n5861 & n12670) | (n5863 & n12670);
  assign n12672 = n5854 | n12599;
  assign n12673 = (n5854 & n5856) | (n5854 & n12672) | (n5856 & n12672);
  assign n12674 = n5847 | n12601;
  assign n12675 = (n5847 & n5849) | (n5847 & n12674) | (n5849 & n12674);
  assign n12676 = n5840 | n5842;
  assign n12677 = (n15927 & n5840) | (n15927 & n12676) | (n5840 & n12676);
  assign n12678 = n5833 | n5835;
  assign n12679 = (n5833 & n12603) | (n5833 & n12678) | (n12603 & n12678);
  assign n12680 = n5826 | n5828;
  assign n12681 = (n5826 & n12605) | (n5826 & n12680) | (n12605 & n12680);
  assign n12682 = n5819 | n5821;
  assign n12683 = (n5819 & n12607) | (n5819 & n12682) | (n12607 & n12682);
  assign n12684 = n5812 | n5814;
  assign n12685 = (n5812 & n12609) | (n5812 & n12684) | (n12609 & n12684);
  assign n12686 = n5805 | n5807;
  assign n12687 = (n5805 & n12611) | (n5805 & n12686) | (n12611 & n12686);
  assign n12688 = n5798 | n5800;
  assign n12689 = (n5798 & n12613) | (n5798 & n12688) | (n12613 & n12688);
  assign n12691 = n5784 | n5786;
  assign n15967 = n5619 | n5784;
  assign n15968 = (n5784 & n5786) | (n5784 & n15967) | (n5786 & n15967);
  assign n15969 = (n12586 & n12691) | (n12586 & n15968) | (n12691 & n15968);
  assign n15970 = (n5621 & n12691) | (n5621 & n15968) | (n12691 & n15968);
  assign n15971 = (n12525 & n15969) | (n12525 & n15970) | (n15969 & n15970);
  assign n12696 = n5763 | n5765;
  assign n15972 = n5598 | n5763;
  assign n15973 = (n5763 & n5765) | (n5763 & n15972) | (n5765 & n15972);
  assign n15974 = (n12577 & n12696) | (n12577 & n15973) | (n12696 & n15973);
  assign n15975 = (n12576 & n12696) | (n12576 & n15973) | (n12696 & n15973);
  assign n15976 = (n15861 & n15974) | (n15861 & n15975) | (n15974 & n15975);
  assign n5906 = x71 & x80;
  assign n5907 = x70 & x81;
  assign n5908 = n5906 & n5907;
  assign n5909 = n5906 | n5907;
  assign n5910 = ~n5908 & n5909;
  assign n15984 = n5735 | n5737;
  assign n15985 = (n5735 & n15938) | (n5735 & n15984) | (n15938 & n15984);
  assign n12709 = n5910 & n15985;
  assign n15986 = (n5735 & n12628) | (n5735 & n15984) | (n12628 & n15984);
  assign n12710 = n5910 & n15986;
  assign n15987 = (n12709 & n12710) | (n12709 & n15881) | (n12710 & n15881);
  assign n15988 = (n12709 & n12710) | (n12709 & n15879) | (n12710 & n15879);
  assign n15989 = (n15760 & n15987) | (n15760 & n15988) | (n15987 & n15988);
  assign n12712 = n5910 | n15985;
  assign n12713 = n5910 | n15986;
  assign n15990 = (n12712 & n12713) | (n12712 & n15881) | (n12713 & n15881);
  assign n15991 = (n12712 & n12713) | (n12712 & n15879) | (n12713 & n15879);
  assign n15992 = (n15760 & n15990) | (n15760 & n15991) | (n15990 & n15991);
  assign n5913 = ~n15989 & n15992;
  assign n5914 = x69 & x82;
  assign n5915 = n5913 & n5914;
  assign n5916 = n5913 | n5914;
  assign n5917 = ~n5915 & n5916;
  assign n15981 = n5742 | n5744;
  assign n49886 = n5917 & n15981;
  assign n49887 = n5742 & n5917;
  assign n49888 = (n15946 & n49886) | (n15946 & n49887) | (n49886 & n49887);
  assign n15982 = (n5742 & n15948) | (n5742 & n15981) | (n15948 & n15981);
  assign n15994 = n5917 & n15982;
  assign n15995 = (n15874 & n49888) | (n15874 & n15994) | (n49888 & n15994);
  assign n49889 = n5917 | n15981;
  assign n49890 = n5742 | n5917;
  assign n49891 = (n15946 & n49889) | (n15946 & n49890) | (n49889 & n49890);
  assign n15997 = n5917 | n15982;
  assign n15998 = (n15874 & n49891) | (n15874 & n15997) | (n49891 & n15997);
  assign n5920 = ~n15995 & n15998;
  assign n5921 = x68 & x83;
  assign n5922 = n5920 & n5921;
  assign n5923 = n5920 | n5921;
  assign n5924 = ~n5922 & n5923;
  assign n12701 = n5749 | n5751;
  assign n12715 = n5924 & n12701;
  assign n12716 = n5749 & n5924;
  assign n15999 = (n12715 & n12716) | (n12715 & n15934) | (n12716 & n15934);
  assign n16000 = (n12715 & n12716) | (n12715 & n15936) | (n12716 & n15936);
  assign n16001 = (n15868 & n15999) | (n15868 & n16000) | (n15999 & n16000);
  assign n12718 = n5924 | n12701;
  assign n12719 = n5749 | n5924;
  assign n16002 = (n12718 & n12719) | (n12718 & n15934) | (n12719 & n15934);
  assign n16003 = (n12718 & n12719) | (n12718 & n15936) | (n12719 & n15936);
  assign n16004 = (n15868 & n16002) | (n15868 & n16003) | (n16002 & n16003);
  assign n5927 = ~n16001 & n16004;
  assign n5928 = x67 & x84;
  assign n5929 = n5927 & n5928;
  assign n5930 = n5927 | n5928;
  assign n5931 = ~n5929 & n5930;
  assign n15979 = n5756 | n5758;
  assign n15980 = (n5756 & n12619) | (n5756 & n15979) | (n12619 & n15979);
  assign n16005 = n5931 & n15980;
  assign n15977 = n5591 | n5756;
  assign n15978 = (n5756 & n5758) | (n5756 & n15977) | (n5758 & n15977);
  assign n16006 = n5931 & n15978;
  assign n16007 = (n15911 & n16005) | (n15911 & n16006) | (n16005 & n16006);
  assign n16008 = n5931 | n15980;
  assign n16009 = n5931 | n15978;
  assign n16010 = (n15911 & n16008) | (n15911 & n16009) | (n16008 & n16009);
  assign n5934 = ~n16007 & n16010;
  assign n5935 = x66 & x85;
  assign n5936 = n5934 & n5935;
  assign n5937 = n5934 | n5935;
  assign n5938 = ~n5936 & n5937;
  assign n5939 = n15976 & n5938;
  assign n5940 = n15976 | n5938;
  assign n5941 = ~n5939 & n5940;
  assign n5942 = x65 & x86;
  assign n5943 = n5941 & n5942;
  assign n5944 = n5941 | n5942;
  assign n5945 = ~n5943 & n5944;
  assign n12693 = n5770 | n5772;
  assign n12721 = n5945 & n12693;
  assign n12722 = n5770 & n5945;
  assign n12723 = (n15932 & n12721) | (n15932 & n12722) | (n12721 & n12722);
  assign n12724 = n5945 | n12693;
  assign n12725 = n5770 | n5945;
  assign n12726 = (n15932 & n12724) | (n15932 & n12725) | (n12724 & n12725);
  assign n5948 = ~n12723 & n12726;
  assign n5949 = x64 & x87;
  assign n5950 = n5948 & n5949;
  assign n5951 = n5948 | n5949;
  assign n5952 = ~n5950 & n5951;
  assign n12727 = n5777 & n5952;
  assign n16011 = (n5952 & n12653) | (n5952 & n12727) | (n12653 & n12727);
  assign n16012 = (n5952 & n12652) | (n5952 & n12727) | (n12652 & n12727);
  assign n16013 = (n15906 & n16011) | (n15906 & n16012) | (n16011 & n16012);
  assign n12729 = n5777 | n5952;
  assign n16014 = n12653 | n12729;
  assign n16015 = n12652 | n12729;
  assign n16016 = (n15906 & n16014) | (n15906 & n16015) | (n16014 & n16015);
  assign n5955 = ~n16013 & n16016;
  assign n5956 = x63 & x88;
  assign n5957 = n5955 & n5956;
  assign n5958 = n5955 | n5956;
  assign n5959 = ~n5957 & n5958;
  assign n5960 = n15971 & n5959;
  assign n5961 = n15971 | n5959;
  assign n5962 = ~n5960 & n5961;
  assign n5963 = x62 & x89;
  assign n5964 = n5962 & n5963;
  assign n5965 = n5962 | n5963;
  assign n5966 = ~n5964 & n5965;
  assign n12731 = n5791 & n5966;
  assign n12732 = (n5966 & n12663) | (n5966 & n12731) | (n12663 & n12731);
  assign n12733 = n5791 | n5966;
  assign n12734 = n12663 | n12733;
  assign n5969 = ~n12732 & n12734;
  assign n5970 = x61 & x90;
  assign n5971 = n5969 & n5970;
  assign n5972 = n5969 | n5970;
  assign n5973 = ~n5971 & n5972;
  assign n5974 = n12689 & n5973;
  assign n5975 = n12689 | n5973;
  assign n5976 = ~n5974 & n5975;
  assign n5977 = x60 & x91;
  assign n5978 = n5976 & n5977;
  assign n5979 = n5976 | n5977;
  assign n5980 = ~n5978 & n5979;
  assign n5981 = n12687 & n5980;
  assign n5982 = n12687 | n5980;
  assign n5983 = ~n5981 & n5982;
  assign n5984 = x59 & x92;
  assign n5985 = n5983 & n5984;
  assign n5986 = n5983 | n5984;
  assign n5987 = ~n5985 & n5986;
  assign n5988 = n12685 & n5987;
  assign n5989 = n12685 | n5987;
  assign n5990 = ~n5988 & n5989;
  assign n5991 = x58 & x93;
  assign n5992 = n5990 & n5991;
  assign n5993 = n5990 | n5991;
  assign n5994 = ~n5992 & n5993;
  assign n5995 = n12683 & n5994;
  assign n5996 = n12683 | n5994;
  assign n5997 = ~n5995 & n5996;
  assign n5998 = x57 & x94;
  assign n5999 = n5997 & n5998;
  assign n6000 = n5997 | n5998;
  assign n6001 = ~n5999 & n6000;
  assign n6002 = n12681 & n6001;
  assign n6003 = n12681 | n6001;
  assign n6004 = ~n6002 & n6003;
  assign n6005 = x56 & x95;
  assign n6006 = n6004 & n6005;
  assign n6007 = n6004 | n6005;
  assign n6008 = ~n6006 & n6007;
  assign n6009 = n12679 & n6008;
  assign n6010 = n12679 | n6008;
  assign n6011 = ~n6009 & n6010;
  assign n6012 = x55 & x96;
  assign n6013 = n6011 & n6012;
  assign n6014 = n6011 | n6012;
  assign n6015 = ~n6013 & n6014;
  assign n6016 = n12677 & n6015;
  assign n6017 = n12677 | n6015;
  assign n6018 = ~n6016 & n6017;
  assign n6019 = x54 & x97;
  assign n6020 = n6018 & n6019;
  assign n6021 = n6018 | n6019;
  assign n6022 = ~n6020 & n6021;
  assign n6023 = n12675 & n6022;
  assign n6024 = n12675 | n6022;
  assign n6025 = ~n6023 & n6024;
  assign n6026 = x53 & x98;
  assign n6027 = n6025 & n6026;
  assign n6028 = n6025 | n6026;
  assign n6029 = ~n6027 & n6028;
  assign n6030 = n12673 & n6029;
  assign n6031 = n12673 | n6029;
  assign n6032 = ~n6030 & n6031;
  assign n6033 = x52 & x99;
  assign n6034 = n6032 & n6033;
  assign n6035 = n6032 | n6033;
  assign n6036 = ~n6034 & n6035;
  assign n6037 = n12671 & n6036;
  assign n6038 = n12671 | n6036;
  assign n6039 = ~n6037 & n6038;
  assign n6040 = x51 & x100;
  assign n6041 = n6039 & n6040;
  assign n6042 = n6039 | n6040;
  assign n6043 = ~n6041 & n6042;
  assign n6044 = n12669 & n6043;
  assign n6045 = n12669 | n6043;
  assign n6046 = ~n6044 & n6045;
  assign n6047 = x50 & x101;
  assign n6048 = n6046 & n6047;
  assign n6049 = n6046 | n6047;
  assign n6050 = ~n6048 & n6049;
  assign n6051 = n12667 & n6050;
  assign n6052 = n12667 | n6050;
  assign n6053 = ~n6051 & n6052;
  assign n6054 = x49 & x102;
  assign n6055 = n6053 & n6054;
  assign n6056 = n6053 | n6054;
  assign n6057 = ~n6055 & n6056;
  assign n6058 = n5882 & n6057;
  assign n6059 = n5882 | n6057;
  assign n6060 = ~n6058 & n6059;
  assign n6061 = x48 & x103;
  assign n6062 = n6060 & n6061;
  assign n6063 = n6060 | n6061;
  assign n6064 = ~n6062 & n6063;
  assign n49892 = n5881 | n6054;
  assign n49893 = (n5880 & n6054) | (n5880 & n49892) | (n6054 & n49892);
  assign n16018 = (n5882 & n6053) | (n5882 & n49893) | (n6053 & n49893);
  assign n12736 = (n6055 & n6057) | (n6055 & n16018) | (n6057 & n16018);
  assign n16019 = n6048 | n12667;
  assign n16020 = (n6048 & n6050) | (n6048 & n16019) | (n6050 & n16019);
  assign n6067 = n6041 | n6044;
  assign n6068 = n6034 | n6037;
  assign n6069 = n6027 | n6030;
  assign n6070 = n6020 | n6023;
  assign n12737 = n6013 | n6015;
  assign n12738 = (n6013 & n12677) | (n6013 & n12737) | (n12677 & n12737);
  assign n12739 = n6006 | n6008;
  assign n12740 = (n6006 & n12679) | (n6006 & n12739) | (n12679 & n12739);
  assign n12741 = n5999 | n6001;
  assign n12742 = (n5999 & n12681) | (n5999 & n12741) | (n12681 & n12741);
  assign n12743 = n5992 | n5994;
  assign n12744 = (n5992 & n12683) | (n5992 & n12743) | (n12683 & n12743);
  assign n12745 = n5985 | n5987;
  assign n12746 = (n5985 & n12685) | (n5985 & n12745) | (n12685 & n12745);
  assign n12747 = n5978 | n5980;
  assign n12748 = (n5978 & n12687) | (n5978 & n12747) | (n12687 & n12747);
  assign n12749 = n5971 | n5973;
  assign n12750 = (n5971 & n12689) | (n5971 & n12749) | (n12689 & n12749);
  assign n12754 = n5950 | n5952;
  assign n16021 = n5777 | n5950;
  assign n16022 = (n5950 & n5952) | (n5950 & n16021) | (n5952 & n16021);
  assign n16023 = (n12653 & n12754) | (n12653 & n16022) | (n12754 & n16022);
  assign n16024 = (n12652 & n12754) | (n12652 & n16022) | (n12754 & n16022);
  assign n16025 = (n15906 & n16023) | (n15906 & n16024) | (n16023 & n16024);
  assign n12623 = (n15868 & n15934) | (n15868 & n15936) | (n15934 & n15936);
  assign n6087 = x72 & x80;
  assign n6088 = x71 & x81;
  assign n6089 = n6087 & n6088;
  assign n6090 = n6087 | n6088;
  assign n6091 = ~n6089 & n6090;
  assign n16026 = n5908 | n5910;
  assign n16028 = n6091 & n16026;
  assign n16029 = n5908 & n6091;
  assign n16030 = (n15985 & n16028) | (n15985 & n16029) | (n16028 & n16029);
  assign n16032 = (n15986 & n16028) | (n15986 & n16029) | (n16028 & n16029);
  assign n16033 = (n15881 & n16030) | (n15881 & n16032) | (n16030 & n16032);
  assign n16034 = (n15879 & n16030) | (n15879 & n16032) | (n16030 & n16032);
  assign n16035 = (n15760 & n16033) | (n15760 & n16034) | (n16033 & n16034);
  assign n16036 = n6091 | n16026;
  assign n16037 = n5908 | n6091;
  assign n16038 = (n15985 & n16036) | (n15985 & n16037) | (n16036 & n16037);
  assign n16039 = (n15986 & n16036) | (n15986 & n16037) | (n16036 & n16037);
  assign n16040 = (n15881 & n16038) | (n15881 & n16039) | (n16038 & n16039);
  assign n16041 = (n15879 & n16038) | (n15879 & n16039) | (n16038 & n16039);
  assign n16042 = (n15760 & n16040) | (n15760 & n16041) | (n16040 & n16041);
  assign n6094 = ~n16035 & n16042;
  assign n6095 = x70 & x82;
  assign n6096 = n6094 & n6095;
  assign n6097 = n6094 | n6095;
  assign n6098 = ~n6096 & n6097;
  assign n12763 = n5915 | n5917;
  assign n12774 = n6098 & n12763;
  assign n12775 = n5915 & n6098;
  assign n15983 = (n5742 & n15946) | (n5742 & n15981) | (n15946 & n15981);
  assign n16043 = (n12774 & n12775) | (n12774 & n15983) | (n12775 & n15983);
  assign n16044 = (n12774 & n12775) | (n12774 & n15982) | (n12775 & n15982);
  assign n16045 = (n15874 & n16043) | (n15874 & n16044) | (n16043 & n16044);
  assign n12777 = n6098 | n12763;
  assign n12778 = n5915 | n6098;
  assign n16046 = (n12777 & n12778) | (n12777 & n15983) | (n12778 & n15983);
  assign n16047 = (n12777 & n12778) | (n12777 & n15982) | (n12778 & n15982);
  assign n16048 = (n15874 & n16046) | (n15874 & n16047) | (n16046 & n16047);
  assign n6101 = ~n16045 & n16048;
  assign n6102 = x69 & x83;
  assign n6103 = n6101 & n6102;
  assign n6104 = n6101 | n6102;
  assign n6105 = ~n6103 & n6104;
  assign n16049 = n5922 | n5924;
  assign n16050 = (n5922 & n12701) | (n5922 & n16049) | (n12701 & n16049);
  assign n12780 = n6105 & n16050;
  assign n16051 = n5749 | n5922;
  assign n16052 = (n5922 & n5924) | (n5922 & n16051) | (n5924 & n16051);
  assign n12781 = n6105 & n16052;
  assign n12782 = (n12623 & n12780) | (n12623 & n12781) | (n12780 & n12781);
  assign n12783 = n6105 | n16050;
  assign n12784 = n6105 | n16052;
  assign n12785 = (n12623 & n12783) | (n12623 & n12784) | (n12783 & n12784);
  assign n6108 = ~n12782 & n12785;
  assign n6109 = x68 & x84;
  assign n6110 = n6108 & n6109;
  assign n6111 = n6108 | n6109;
  assign n6112 = ~n6110 & n6111;
  assign n12758 = n5929 | n5931;
  assign n12786 = n6112 & n12758;
  assign n12787 = n5929 & n6112;
  assign n16053 = (n12786 & n12787) | (n12786 & n15980) | (n12787 & n15980);
  assign n16054 = (n12786 & n12787) | (n12786 & n15978) | (n12787 & n15978);
  assign n16055 = (n15911 & n16053) | (n15911 & n16054) | (n16053 & n16054);
  assign n12789 = n6112 | n12758;
  assign n12790 = n5929 | n6112;
  assign n16056 = (n12789 & n12790) | (n12789 & n15980) | (n12790 & n15980);
  assign n16057 = (n12789 & n12790) | (n12789 & n15978) | (n12790 & n15978);
  assign n16058 = (n15911 & n16056) | (n15911 & n16057) | (n16056 & n16057);
  assign n6115 = ~n16055 & n16058;
  assign n6116 = x67 & x85;
  assign n6117 = n6115 & n6116;
  assign n6118 = n6115 | n6116;
  assign n6119 = ~n6117 & n6118;
  assign n12756 = n5936 | n5938;
  assign n12792 = n6119 & n12756;
  assign n12793 = n5936 & n6119;
  assign n12794 = (n15976 & n12792) | (n15976 & n12793) | (n12792 & n12793);
  assign n12795 = n6119 | n12756;
  assign n12796 = n5936 | n6119;
  assign n12797 = (n15976 & n12795) | (n15976 & n12796) | (n12795 & n12796);
  assign n6122 = ~n12794 & n12797;
  assign n6123 = x66 & x86;
  assign n6124 = n6122 & n6123;
  assign n6125 = n6122 | n6123;
  assign n6126 = ~n6124 & n6125;
  assign n12798 = n5943 & n6126;
  assign n16059 = (n6126 & n12722) | (n6126 & n12798) | (n12722 & n12798);
  assign n16060 = (n6126 & n12721) | (n6126 & n12798) | (n12721 & n12798);
  assign n16061 = (n15932 & n16059) | (n15932 & n16060) | (n16059 & n16060);
  assign n12800 = n5943 | n6126;
  assign n16062 = n12722 | n12800;
  assign n16063 = n12721 | n12800;
  assign n16064 = (n15932 & n16062) | (n15932 & n16063) | (n16062 & n16063);
  assign n6129 = ~n16061 & n16064;
  assign n6130 = x65 & x87;
  assign n6131 = n6129 & n6130;
  assign n6132 = n6129 | n6130;
  assign n6133 = ~n6131 & n6132;
  assign n6134 = n16025 & n6133;
  assign n6135 = n16025 | n6133;
  assign n6136 = ~n6134 & n6135;
  assign n6137 = x64 & x88;
  assign n6138 = n6136 & n6137;
  assign n6139 = n6136 | n6137;
  assign n6140 = ~n6138 & n6139;
  assign n12751 = n5957 | n5959;
  assign n12802 = n6140 & n12751;
  assign n12803 = n5957 & n6140;
  assign n12804 = (n15971 & n12802) | (n15971 & n12803) | (n12802 & n12803);
  assign n12805 = n6140 | n12751;
  assign n12806 = n5957 | n6140;
  assign n12807 = (n15971 & n12805) | (n15971 & n12806) | (n12805 & n12806);
  assign n6143 = ~n12804 & n12807;
  assign n6144 = x63 & x89;
  assign n6145 = n6143 & n6144;
  assign n6146 = n6143 | n6144;
  assign n6147 = ~n6145 & n6146;
  assign n12808 = n5964 & n6147;
  assign n16065 = (n6147 & n12731) | (n6147 & n12808) | (n12731 & n12808);
  assign n16066 = (n5966 & n6147) | (n5966 & n12808) | (n6147 & n12808);
  assign n16067 = (n12663 & n16065) | (n12663 & n16066) | (n16065 & n16066);
  assign n12810 = n5964 | n6147;
  assign n16068 = n12731 | n12810;
  assign n16069 = n5966 | n12810;
  assign n16070 = (n12663 & n16068) | (n12663 & n16069) | (n16068 & n16069);
  assign n6150 = ~n16067 & n16070;
  assign n6151 = x62 & x90;
  assign n6152 = n6150 & n6151;
  assign n6153 = n6150 | n6151;
  assign n6154 = ~n6152 & n6153;
  assign n6155 = n12750 & n6154;
  assign n6156 = n12750 | n6154;
  assign n6157 = ~n6155 & n6156;
  assign n6158 = x61 & x91;
  assign n6159 = n6157 & n6158;
  assign n6160 = n6157 | n6158;
  assign n6161 = ~n6159 & n6160;
  assign n6162 = n12748 & n6161;
  assign n6163 = n12748 | n6161;
  assign n6164 = ~n6162 & n6163;
  assign n6165 = x60 & x92;
  assign n6166 = n6164 & n6165;
  assign n6167 = n6164 | n6165;
  assign n6168 = ~n6166 & n6167;
  assign n6169 = n12746 & n6168;
  assign n6170 = n12746 | n6168;
  assign n6171 = ~n6169 & n6170;
  assign n6172 = x59 & x93;
  assign n6173 = n6171 & n6172;
  assign n6174 = n6171 | n6172;
  assign n6175 = ~n6173 & n6174;
  assign n6176 = n12744 & n6175;
  assign n6177 = n12744 | n6175;
  assign n6178 = ~n6176 & n6177;
  assign n6179 = x58 & x94;
  assign n6180 = n6178 & n6179;
  assign n6181 = n6178 | n6179;
  assign n6182 = ~n6180 & n6181;
  assign n6183 = n12742 & n6182;
  assign n6184 = n12742 | n6182;
  assign n6185 = ~n6183 & n6184;
  assign n6186 = x57 & x95;
  assign n6187 = n6185 & n6186;
  assign n6188 = n6185 | n6186;
  assign n6189 = ~n6187 & n6188;
  assign n6190 = n12740 & n6189;
  assign n6191 = n12740 | n6189;
  assign n6192 = ~n6190 & n6191;
  assign n6193 = x56 & x96;
  assign n6194 = n6192 & n6193;
  assign n6195 = n6192 | n6193;
  assign n6196 = ~n6194 & n6195;
  assign n6197 = n12738 & n6196;
  assign n6198 = n12738 | n6196;
  assign n6199 = ~n6197 & n6198;
  assign n6200 = x55 & x97;
  assign n6201 = n6199 & n6200;
  assign n6202 = n6199 | n6200;
  assign n6203 = ~n6201 & n6202;
  assign n6204 = n6070 & n6203;
  assign n6205 = n6070 | n6203;
  assign n6206 = ~n6204 & n6205;
  assign n6207 = x54 & x98;
  assign n6208 = n6206 & n6207;
  assign n6209 = n6206 | n6207;
  assign n6210 = ~n6208 & n6209;
  assign n6211 = n6069 & n6210;
  assign n6212 = n6069 | n6210;
  assign n6213 = ~n6211 & n6212;
  assign n6214 = x53 & x99;
  assign n6215 = n6213 & n6214;
  assign n6216 = n6213 | n6214;
  assign n6217 = ~n6215 & n6216;
  assign n6218 = n6068 & n6217;
  assign n6219 = n6068 | n6217;
  assign n6220 = ~n6218 & n6219;
  assign n6221 = x52 & x100;
  assign n6222 = n6220 & n6221;
  assign n6223 = n6220 | n6221;
  assign n6224 = ~n6222 & n6223;
  assign n6225 = n6067 & n6224;
  assign n6226 = n6067 | n6224;
  assign n6227 = ~n6225 & n6226;
  assign n6228 = x51 & x101;
  assign n6229 = n6227 & n6228;
  assign n6230 = n6227 | n6228;
  assign n6231 = ~n6229 & n6230;
  assign n6232 = n16020 & n6231;
  assign n6233 = n16020 | n6231;
  assign n6234 = ~n6232 & n6233;
  assign n6235 = x50 & x102;
  assign n6236 = n6234 & n6235;
  assign n6237 = n6234 | n6235;
  assign n6238 = ~n6236 & n6237;
  assign n6239 = n12736 & n6238;
  assign n6240 = n12736 | n6238;
  assign n6241 = ~n6239 & n6240;
  assign n6242 = x49 & x103;
  assign n6243 = n6241 & n6242;
  assign n6244 = n6241 | n6242;
  assign n6245 = ~n6243 & n6244;
  assign n6246 = n6062 & n6245;
  assign n6247 = n6062 | n6245;
  assign n6248 = ~n6246 & n6247;
  assign n6249 = x48 & x104;
  assign n6250 = n6248 & n6249;
  assign n6251 = n6248 | n6249;
  assign n6252 = ~n6250 & n6251;
  assign n49894 = n6061 | n6242;
  assign n49895 = (n6060 & n6242) | (n6060 & n49894) | (n6242 & n49894);
  assign n16072 = (n6062 & n6241) | (n6062 & n49895) | (n6241 & n49895);
  assign n12813 = (n6243 & n6245) | (n6243 & n16072) | (n6245 & n16072);
  assign n12814 = n6236 | n12736;
  assign n12815 = (n6236 & n6238) | (n6236 & n12814) | (n6238 & n12814);
  assign n16073 = n6229 | n16020;
  assign n16074 = (n6229 & n6231) | (n6229 & n16073) | (n6231 & n16073);
  assign n6256 = n6222 | n6225;
  assign n6257 = n6215 | n6218;
  assign n6258 = n6208 | n6211;
  assign n12816 = n6201 | n6203;
  assign n12817 = (n6070 & n6201) | (n6070 & n12816) | (n6201 & n12816);
  assign n12818 = n6194 | n6196;
  assign n12819 = (n6194 & n12738) | (n6194 & n12818) | (n12738 & n12818);
  assign n12820 = n6187 | n6189;
  assign n12821 = (n6187 & n12740) | (n6187 & n12820) | (n12740 & n12820);
  assign n12822 = n6180 | n6182;
  assign n12823 = (n6180 & n12742) | (n6180 & n12822) | (n12742 & n12822);
  assign n12824 = n6173 | n6175;
  assign n12825 = (n6173 & n12744) | (n6173 & n12824) | (n12744 & n12824);
  assign n12826 = n6166 | n6168;
  assign n12827 = (n6166 & n12746) | (n6166 & n12826) | (n12746 & n12826);
  assign n12828 = n6159 | n6161;
  assign n12829 = (n6159 & n12748) | (n6159 & n12828) | (n12748 & n12828);
  assign n12833 = n6145 | n6147;
  assign n16075 = n5964 | n6145;
  assign n16076 = (n6145 & n6147) | (n6145 & n16075) | (n6147 & n16075);
  assign n16077 = (n12731 & n12833) | (n12731 & n16076) | (n12833 & n16076);
  assign n16078 = (n5966 & n12833) | (n5966 & n16076) | (n12833 & n16076);
  assign n16079 = (n12663 & n16077) | (n12663 & n16078) | (n16077 & n16078);
  assign n12838 = n6124 | n6126;
  assign n16080 = n5943 | n6124;
  assign n16081 = (n6124 & n6126) | (n6124 & n16080) | (n6126 & n16080);
  assign n16082 = (n12722 & n12838) | (n12722 & n16081) | (n12838 & n16081);
  assign n16083 = (n12721 & n12838) | (n12721 & n16081) | (n12838 & n16081);
  assign n16084 = (n15932 & n16082) | (n15932 & n16083) | (n16082 & n16083);
  assign n12700 = (n15911 & n15978) | (n15911 & n15980) | (n15978 & n15980);
  assign n12846 = n6089 | n16030;
  assign n12847 = n6089 | n16032;
  assign n16087 = (n12846 & n12847) | (n12846 & n15881) | (n12847 & n15881);
  assign n16088 = (n12846 & n12847) | (n12846 & n15879) | (n12847 & n15879);
  assign n16089 = (n15760 & n16087) | (n15760 & n16088) | (n16087 & n16088);
  assign n6276 = x73 & x80;
  assign n6277 = x72 & x81;
  assign n6278 = n6276 & n6277;
  assign n6279 = n6276 | n6277;
  assign n6280 = ~n6278 & n6279;
  assign n6281 = n16089 & n6280;
  assign n6282 = n16089 | n6280;
  assign n6283 = ~n6281 & n6282;
  assign n6284 = x71 & x82;
  assign n6285 = n6283 & n6284;
  assign n6286 = n6283 | n6284;
  assign n6287 = ~n6285 & n6286;
  assign n16090 = n6096 | n6098;
  assign n16091 = (n6096 & n12763) | (n6096 & n16090) | (n12763 & n16090);
  assign n12849 = n6287 & n16091;
  assign n16092 = n5915 | n6096;
  assign n16093 = (n6096 & n6098) | (n6096 & n16092) | (n6098 & n16092);
  assign n12850 = n6287 & n16093;
  assign n16094 = (n12849 & n12850) | (n12849 & n15983) | (n12850 & n15983);
  assign n16095 = (n12849 & n12850) | (n12849 & n15982) | (n12850 & n15982);
  assign n16096 = (n15874 & n16094) | (n15874 & n16095) | (n16094 & n16095);
  assign n12852 = n6287 | n16091;
  assign n12853 = n6287 | n16093;
  assign n16097 = (n12852 & n12853) | (n12852 & n15983) | (n12853 & n15983);
  assign n16098 = (n12852 & n12853) | (n12852 & n15982) | (n12853 & n15982);
  assign n16099 = (n15874 & n16097) | (n15874 & n16098) | (n16097 & n16098);
  assign n6290 = ~n16096 & n16099;
  assign n6291 = x70 & x83;
  assign n6292 = n6290 & n6291;
  assign n6293 = n6290 | n6291;
  assign n6294 = ~n6292 & n6293;
  assign n12855 = n6103 & n6294;
  assign n49896 = (n6105 & n6294) | (n6105 & n12855) | (n6294 & n12855);
  assign n49897 = n6294 & n12855;
  assign n49898 = (n16050 & n49896) | (n16050 & n49897) | (n49896 & n49897);
  assign n16101 = (n6294 & n12781) | (n6294 & n12855) | (n12781 & n12855);
  assign n16102 = (n12623 & n49898) | (n12623 & n16101) | (n49898 & n16101);
  assign n12857 = n6103 | n6294;
  assign n49899 = n6105 | n12857;
  assign n49900 = (n12857 & n16050) | (n12857 & n49899) | (n16050 & n49899);
  assign n16104 = n12781 | n12857;
  assign n16105 = (n12623 & n49900) | (n12623 & n16104) | (n49900 & n16104);
  assign n6297 = ~n16102 & n16105;
  assign n6298 = x69 & x84;
  assign n6299 = n6297 & n6298;
  assign n6300 = n6297 | n6298;
  assign n6301 = ~n6299 & n6300;
  assign n49901 = n6110 & n6301;
  assign n49902 = (n6301 & n12786) | (n6301 & n49901) | (n12786 & n49901);
  assign n16085 = n5929 | n6110;
  assign n16086 = (n6110 & n6112) | (n6110 & n16085) | (n6112 & n16085);
  assign n16107 = n6301 & n16086;
  assign n16108 = (n12700 & n49902) | (n12700 & n16107) | (n49902 & n16107);
  assign n49903 = n6110 | n6301;
  assign n49904 = n12786 | n49903;
  assign n16110 = n6301 | n16086;
  assign n16111 = (n12700 & n49904) | (n12700 & n16110) | (n49904 & n16110);
  assign n6304 = ~n16108 & n16111;
  assign n6305 = x68 & x85;
  assign n6306 = n6304 & n6305;
  assign n6307 = n6304 | n6305;
  assign n6308 = ~n6306 & n6307;
  assign n12859 = n6117 & n6308;
  assign n16112 = (n6308 & n12792) | (n6308 & n12859) | (n12792 & n12859);
  assign n16113 = (n6308 & n12793) | (n6308 & n12859) | (n12793 & n12859);
  assign n16114 = (n15976 & n16112) | (n15976 & n16113) | (n16112 & n16113);
  assign n12861 = n6117 | n6308;
  assign n16115 = n12792 | n12861;
  assign n16116 = n12793 | n12861;
  assign n16117 = (n15976 & n16115) | (n15976 & n16116) | (n16115 & n16116);
  assign n6311 = ~n16114 & n16117;
  assign n6312 = x67 & x86;
  assign n6313 = n6311 & n6312;
  assign n6314 = n6311 | n6312;
  assign n6315 = ~n6313 & n6314;
  assign n6316 = n16084 & n6315;
  assign n6317 = n16084 | n6315;
  assign n6318 = ~n6316 & n6317;
  assign n6319 = x66 & x87;
  assign n6320 = n6318 & n6319;
  assign n6321 = n6318 | n6319;
  assign n6322 = ~n6320 & n6321;
  assign n12835 = n6131 | n6133;
  assign n12863 = n6322 & n12835;
  assign n12864 = n6131 & n6322;
  assign n12865 = (n16025 & n12863) | (n16025 & n12864) | (n12863 & n12864);
  assign n12866 = n6322 | n12835;
  assign n12867 = n6131 | n6322;
  assign n12868 = (n16025 & n12866) | (n16025 & n12867) | (n12866 & n12867);
  assign n6325 = ~n12865 & n12868;
  assign n6326 = x65 & x88;
  assign n6327 = n6325 & n6326;
  assign n6328 = n6325 | n6326;
  assign n6329 = ~n6327 & n6328;
  assign n12869 = n6138 & n6329;
  assign n16118 = (n6329 & n12803) | (n6329 & n12869) | (n12803 & n12869);
  assign n16119 = (n6329 & n12802) | (n6329 & n12869) | (n12802 & n12869);
  assign n16120 = (n15971 & n16118) | (n15971 & n16119) | (n16118 & n16119);
  assign n12871 = n6138 | n6329;
  assign n16121 = n12803 | n12871;
  assign n16122 = n12802 | n12871;
  assign n16123 = (n15971 & n16121) | (n15971 & n16122) | (n16121 & n16122);
  assign n6332 = ~n16120 & n16123;
  assign n6333 = x64 & x89;
  assign n6334 = n6332 & n6333;
  assign n6335 = n6332 | n6333;
  assign n6336 = ~n6334 & n6335;
  assign n6337 = n16079 & n6336;
  assign n6338 = n16079 | n6336;
  assign n6339 = ~n6337 & n6338;
  assign n6340 = x63 & x90;
  assign n6341 = n6339 & n6340;
  assign n6342 = n6339 | n6340;
  assign n6343 = ~n6341 & n6342;
  assign n12830 = n6152 | n6154;
  assign n16124 = n6343 & n12830;
  assign n16125 = n6152 & n6343;
  assign n16126 = (n12750 & n16124) | (n12750 & n16125) | (n16124 & n16125);
  assign n16127 = n6343 | n12830;
  assign n16128 = n6152 | n6343;
  assign n16129 = (n12750 & n16127) | (n12750 & n16128) | (n16127 & n16128);
  assign n6346 = ~n16126 & n16129;
  assign n6347 = x62 & x91;
  assign n6348 = n6346 & n6347;
  assign n6349 = n6346 | n6347;
  assign n6350 = ~n6348 & n6349;
  assign n6351 = n12829 & n6350;
  assign n6352 = n12829 | n6350;
  assign n6353 = ~n6351 & n6352;
  assign n6354 = x61 & x92;
  assign n6355 = n6353 & n6354;
  assign n6356 = n6353 | n6354;
  assign n6357 = ~n6355 & n6356;
  assign n6358 = n12827 & n6357;
  assign n6359 = n12827 | n6357;
  assign n6360 = ~n6358 & n6359;
  assign n6361 = x60 & x93;
  assign n6362 = n6360 & n6361;
  assign n6363 = n6360 | n6361;
  assign n6364 = ~n6362 & n6363;
  assign n6365 = n12825 & n6364;
  assign n6366 = n12825 | n6364;
  assign n6367 = ~n6365 & n6366;
  assign n6368 = x59 & x94;
  assign n6369 = n6367 & n6368;
  assign n6370 = n6367 | n6368;
  assign n6371 = ~n6369 & n6370;
  assign n6372 = n12823 & n6371;
  assign n6373 = n12823 | n6371;
  assign n6374 = ~n6372 & n6373;
  assign n6375 = x58 & x95;
  assign n6376 = n6374 & n6375;
  assign n6377 = n6374 | n6375;
  assign n6378 = ~n6376 & n6377;
  assign n6379 = n12821 & n6378;
  assign n6380 = n12821 | n6378;
  assign n6381 = ~n6379 & n6380;
  assign n6382 = x57 & x96;
  assign n6383 = n6381 & n6382;
  assign n6384 = n6381 | n6382;
  assign n6385 = ~n6383 & n6384;
  assign n6386 = n12819 & n6385;
  assign n6387 = n12819 | n6385;
  assign n6388 = ~n6386 & n6387;
  assign n6389 = x56 & x97;
  assign n6390 = n6388 & n6389;
  assign n6391 = n6388 | n6389;
  assign n6392 = ~n6390 & n6391;
  assign n6393 = n12817 & n6392;
  assign n6394 = n12817 | n6392;
  assign n6395 = ~n6393 & n6394;
  assign n6396 = x55 & x98;
  assign n6397 = n6395 & n6396;
  assign n6398 = n6395 | n6396;
  assign n6399 = ~n6397 & n6398;
  assign n6400 = n6258 & n6399;
  assign n6401 = n6258 | n6399;
  assign n6402 = ~n6400 & n6401;
  assign n6403 = x54 & x99;
  assign n6404 = n6402 & n6403;
  assign n6405 = n6402 | n6403;
  assign n6406 = ~n6404 & n6405;
  assign n6407 = n6257 & n6406;
  assign n6408 = n6257 | n6406;
  assign n6409 = ~n6407 & n6408;
  assign n6410 = x53 & x100;
  assign n6411 = n6409 & n6410;
  assign n6412 = n6409 | n6410;
  assign n6413 = ~n6411 & n6412;
  assign n6414 = n6256 & n6413;
  assign n6415 = n6256 | n6413;
  assign n6416 = ~n6414 & n6415;
  assign n6417 = x52 & x101;
  assign n6418 = n6416 & n6417;
  assign n6419 = n6416 | n6417;
  assign n6420 = ~n6418 & n6419;
  assign n6421 = n16074 & n6420;
  assign n6422 = n16074 | n6420;
  assign n6423 = ~n6421 & n6422;
  assign n6424 = x51 & x102;
  assign n6425 = n6423 & n6424;
  assign n6426 = n6423 | n6424;
  assign n6427 = ~n6425 & n6426;
  assign n6428 = n12815 & n6427;
  assign n6429 = n12815 | n6427;
  assign n6430 = ~n6428 & n6429;
  assign n6431 = x50 & x103;
  assign n6432 = n6430 & n6431;
  assign n6433 = n6430 | n6431;
  assign n6434 = ~n6432 & n6433;
  assign n6435 = n12813 & n6434;
  assign n6436 = n12813 | n6434;
  assign n6437 = ~n6435 & n6436;
  assign n6438 = x49 & x104;
  assign n6439 = n6437 & n6438;
  assign n6440 = n6437 | n6438;
  assign n6441 = ~n6439 & n6440;
  assign n6442 = n6250 & n6441;
  assign n6443 = n6250 | n6441;
  assign n6444 = ~n6442 & n6443;
  assign n6445 = x48 & x105;
  assign n6446 = n6444 & n6445;
  assign n6447 = n6444 | n6445;
  assign n6448 = ~n6446 & n6447;
  assign n49905 = n6249 | n6438;
  assign n49906 = (n6248 & n6438) | (n6248 & n49905) | (n6438 & n49905);
  assign n16131 = (n6250 & n6437) | (n6250 & n49906) | (n6437 & n49906);
  assign n12874 = (n6439 & n6441) | (n6439 & n16131) | (n6441 & n16131);
  assign n12875 = n6432 | n12813;
  assign n12876 = (n6432 & n6434) | (n6432 & n12875) | (n6434 & n12875);
  assign n12877 = n6425 | n12815;
  assign n12878 = (n6425 & n6427) | (n6425 & n12877) | (n6427 & n12877);
  assign n16132 = n6418 | n16074;
  assign n16133 = (n6418 & n6420) | (n6418 & n16132) | (n6420 & n16132);
  assign n6453 = n6411 | n6414;
  assign n6454 = n6404 | n6407;
  assign n12879 = n6397 | n6399;
  assign n12880 = (n6258 & n6397) | (n6258 & n12879) | (n6397 & n12879);
  assign n12881 = n6390 | n6392;
  assign n12882 = (n6390 & n12817) | (n6390 & n12881) | (n12817 & n12881);
  assign n12883 = n6383 | n6385;
  assign n12884 = (n6383 & n12819) | (n6383 & n12883) | (n12819 & n12883);
  assign n12885 = n6376 | n6378;
  assign n12886 = (n6376 & n12821) | (n6376 & n12885) | (n12821 & n12885);
  assign n12887 = n6369 | n6371;
  assign n12888 = (n6369 & n12823) | (n6369 & n12887) | (n12823 & n12887);
  assign n12889 = n6362 | n6364;
  assign n12890 = (n6362 & n12825) | (n6362 & n12889) | (n12825 & n12889);
  assign n12891 = n6355 | n6357;
  assign n12892 = (n6355 & n12827) | (n6355 & n12891) | (n12827 & n12891);
  assign n12831 = (n6152 & n12750) | (n6152 & n12830) | (n12750 & n12830);
  assign n12900 = n6327 | n6329;
  assign n16134 = n6138 | n6327;
  assign n16135 = (n6327 & n6329) | (n6327 & n16134) | (n6329 & n16134);
  assign n16136 = (n12803 & n12900) | (n12803 & n16135) | (n12900 & n16135);
  assign n16137 = (n12802 & n12900) | (n12802 & n16135) | (n12900 & n16135);
  assign n16138 = (n15971 & n16136) | (n15971 & n16137) | (n16136 & n16137);
  assign n12905 = n6306 | n6308;
  assign n16139 = n6117 | n6306;
  assign n16140 = (n6306 & n6308) | (n6306 & n16139) | (n6308 & n16139);
  assign n16141 = (n12792 & n12905) | (n12792 & n16140) | (n12905 & n16140);
  assign n16142 = (n12793 & n12905) | (n12793 & n16140) | (n12905 & n16140);
  assign n16143 = (n15976 & n16141) | (n15976 & n16142) | (n16141 & n16142);
  assign n12840 = n6110 | n12786;
  assign n12913 = n6285 | n12850;
  assign n16144 = n6285 | n6287;
  assign n16145 = (n6285 & n16091) | (n6285 & n16144) | (n16091 & n16144);
  assign n16146 = (n12913 & n15983) | (n12913 & n16145) | (n15983 & n16145);
  assign n16147 = (n12913 & n15982) | (n12913 & n16145) | (n15982 & n16145);
  assign n16148 = (n15874 & n16146) | (n15874 & n16147) | (n16146 & n16147);
  assign n6473 = x74 & x80;
  assign n6474 = x73 & x81;
  assign n6475 = n6473 & n6474;
  assign n6476 = n6473 | n6474;
  assign n6477 = ~n6475 & n6476;
  assign n12915 = n6278 | n6280;
  assign n12917 = n6477 & n12915;
  assign n12918 = n6278 & n6477;
  assign n12919 = (n16089 & n12917) | (n16089 & n12918) | (n12917 & n12918);
  assign n12920 = n6477 | n12915;
  assign n12921 = n6278 | n6477;
  assign n12922 = (n16089 & n12920) | (n16089 & n12921) | (n12920 & n12921);
  assign n6480 = ~n12919 & n12922;
  assign n6481 = x72 & x82;
  assign n6482 = n6480 & n6481;
  assign n6483 = n6480 | n6481;
  assign n6484 = ~n6482 & n6483;
  assign n6485 = n16148 & n6484;
  assign n6486 = n16148 | n6484;
  assign n6487 = ~n6485 & n6486;
  assign n6488 = x71 & x83;
  assign n6489 = n6487 & n6488;
  assign n6490 = n6487 | n6488;
  assign n6491 = ~n6489 & n6490;
  assign n16149 = n6103 | n6292;
  assign n16150 = (n6292 & n6294) | (n6292 & n16149) | (n6294 & n16149);
  assign n12923 = n6491 & n16150;
  assign n12910 = n6292 | n6294;
  assign n12924 = n6491 & n12910;
  assign n16151 = (n12780 & n12923) | (n12780 & n12924) | (n12923 & n12924);
  assign n16152 = (n12781 & n12923) | (n12781 & n12924) | (n12923 & n12924);
  assign n16153 = (n12623 & n16151) | (n12623 & n16152) | (n16151 & n16152);
  assign n12926 = n6491 | n16150;
  assign n12927 = n6491 | n12910;
  assign n16154 = (n12780 & n12926) | (n12780 & n12927) | (n12926 & n12927);
  assign n16155 = (n12781 & n12926) | (n12781 & n12927) | (n12926 & n12927);
  assign n16156 = (n12623 & n16154) | (n12623 & n16155) | (n16154 & n16155);
  assign n6494 = ~n16153 & n16156;
  assign n6495 = x70 & x84;
  assign n6496 = n6494 & n6495;
  assign n6497 = n6494 | n6495;
  assign n6498 = ~n6496 & n6497;
  assign n12907 = n6299 | n6301;
  assign n12929 = n6498 & n12907;
  assign n12930 = n6299 & n6498;
  assign n16157 = (n12840 & n12929) | (n12840 & n12930) | (n12929 & n12930);
  assign n16158 = (n12929 & n12930) | (n12929 & n16086) | (n12930 & n16086);
  assign n16159 = (n12700 & n16157) | (n12700 & n16158) | (n16157 & n16158);
  assign n12932 = n6498 | n12907;
  assign n12933 = n6299 | n6498;
  assign n16160 = (n12840 & n12932) | (n12840 & n12933) | (n12932 & n12933);
  assign n16161 = (n12932 & n12933) | (n12932 & n16086) | (n12933 & n16086);
  assign n16162 = (n12700 & n16160) | (n12700 & n16161) | (n16160 & n16161);
  assign n6501 = ~n16159 & n16162;
  assign n6502 = x69 & x85;
  assign n6503 = n6501 & n6502;
  assign n6504 = n6501 | n6502;
  assign n6505 = ~n6503 & n6504;
  assign n6506 = n16143 & n6505;
  assign n6507 = n16143 | n6505;
  assign n6508 = ~n6506 & n6507;
  assign n6509 = x68 & x86;
  assign n6510 = n6508 & n6509;
  assign n6511 = n6508 | n6509;
  assign n6512 = ~n6510 & n6511;
  assign n12902 = n6313 | n6315;
  assign n12935 = n6512 & n12902;
  assign n12936 = n6313 & n6512;
  assign n12937 = (n16084 & n12935) | (n16084 & n12936) | (n12935 & n12936);
  assign n12938 = n6512 | n12902;
  assign n12939 = n6313 | n6512;
  assign n12940 = (n16084 & n12938) | (n16084 & n12939) | (n12938 & n12939);
  assign n6515 = ~n12937 & n12940;
  assign n6516 = x67 & x87;
  assign n6517 = n6515 & n6516;
  assign n6518 = n6515 | n6516;
  assign n6519 = ~n6517 & n6518;
  assign n12941 = n6320 & n6519;
  assign n16163 = (n6519 & n12864) | (n6519 & n12941) | (n12864 & n12941);
  assign n16164 = (n6519 & n12863) | (n6519 & n12941) | (n12863 & n12941);
  assign n16165 = (n16025 & n16163) | (n16025 & n16164) | (n16163 & n16164);
  assign n12943 = n6320 | n6519;
  assign n16166 = n12864 | n12943;
  assign n16167 = n12863 | n12943;
  assign n16168 = (n16025 & n16166) | (n16025 & n16167) | (n16166 & n16167);
  assign n6522 = ~n16165 & n16168;
  assign n6523 = x66 & x88;
  assign n6524 = n6522 & n6523;
  assign n6525 = n6522 | n6523;
  assign n6526 = ~n6524 & n6525;
  assign n6527 = n16138 & n6526;
  assign n6528 = n16138 | n6526;
  assign n6529 = ~n6527 & n6528;
  assign n6530 = x65 & x89;
  assign n6531 = n6529 & n6530;
  assign n6532 = n6529 | n6530;
  assign n6533 = ~n6531 & n6532;
  assign n12897 = n6334 | n6336;
  assign n12945 = n6533 & n12897;
  assign n12946 = n6334 & n6533;
  assign n12947 = (n16079 & n12945) | (n16079 & n12946) | (n12945 & n12946);
  assign n12948 = n6533 | n12897;
  assign n12949 = n6334 | n6533;
  assign n12950 = (n16079 & n12948) | (n16079 & n12949) | (n12948 & n12949);
  assign n6536 = ~n12947 & n12950;
  assign n6537 = x64 & x90;
  assign n6538 = n6536 & n6537;
  assign n6539 = n6536 | n6537;
  assign n6540 = ~n6538 & n6539;
  assign n12895 = n6341 | n6343;
  assign n16169 = n6540 & n12895;
  assign n16170 = n6341 & n6540;
  assign n16171 = (n12831 & n16169) | (n12831 & n16170) | (n16169 & n16170);
  assign n16172 = n6540 | n12895;
  assign n16173 = n6341 | n6540;
  assign n16174 = (n12831 & n16172) | (n12831 & n16173) | (n16172 & n16173);
  assign n6543 = ~n16171 & n16174;
  assign n6544 = x63 & x91;
  assign n6545 = n6543 & n6544;
  assign n6546 = n6543 | n6544;
  assign n6547 = ~n6545 & n6546;
  assign n12893 = n6348 | n6350;
  assign n16175 = n6547 & n12893;
  assign n16176 = n6348 & n6547;
  assign n16177 = (n12829 & n16175) | (n12829 & n16176) | (n16175 & n16176);
  assign n16178 = n6547 | n12893;
  assign n16179 = n6348 | n6547;
  assign n16180 = (n12829 & n16178) | (n12829 & n16179) | (n16178 & n16179);
  assign n6550 = ~n16177 & n16180;
  assign n6551 = x62 & x92;
  assign n6552 = n6550 & n6551;
  assign n6553 = n6550 | n6551;
  assign n6554 = ~n6552 & n6553;
  assign n6555 = n12892 & n6554;
  assign n6556 = n12892 | n6554;
  assign n6557 = ~n6555 & n6556;
  assign n6558 = x61 & x93;
  assign n6559 = n6557 & n6558;
  assign n6560 = n6557 | n6558;
  assign n6561 = ~n6559 & n6560;
  assign n6562 = n12890 & n6561;
  assign n6563 = n12890 | n6561;
  assign n6564 = ~n6562 & n6563;
  assign n6565 = x60 & x94;
  assign n6566 = n6564 & n6565;
  assign n6567 = n6564 | n6565;
  assign n6568 = ~n6566 & n6567;
  assign n6569 = n12888 & n6568;
  assign n6570 = n12888 | n6568;
  assign n6571 = ~n6569 & n6570;
  assign n6572 = x59 & x95;
  assign n6573 = n6571 & n6572;
  assign n6574 = n6571 | n6572;
  assign n6575 = ~n6573 & n6574;
  assign n6576 = n12886 & n6575;
  assign n6577 = n12886 | n6575;
  assign n6578 = ~n6576 & n6577;
  assign n6579 = x58 & x96;
  assign n6580 = n6578 & n6579;
  assign n6581 = n6578 | n6579;
  assign n6582 = ~n6580 & n6581;
  assign n6583 = n12884 & n6582;
  assign n6584 = n12884 | n6582;
  assign n6585 = ~n6583 & n6584;
  assign n6586 = x57 & x97;
  assign n6587 = n6585 & n6586;
  assign n6588 = n6585 | n6586;
  assign n6589 = ~n6587 & n6588;
  assign n6590 = n12882 & n6589;
  assign n6591 = n12882 | n6589;
  assign n6592 = ~n6590 & n6591;
  assign n6593 = x56 & x98;
  assign n6594 = n6592 & n6593;
  assign n6595 = n6592 | n6593;
  assign n6596 = ~n6594 & n6595;
  assign n6597 = n12880 & n6596;
  assign n6598 = n12880 | n6596;
  assign n6599 = ~n6597 & n6598;
  assign n6600 = x55 & x99;
  assign n6601 = n6599 & n6600;
  assign n6602 = n6599 | n6600;
  assign n6603 = ~n6601 & n6602;
  assign n6604 = n6454 & n6603;
  assign n6605 = n6454 | n6603;
  assign n6606 = ~n6604 & n6605;
  assign n6607 = x54 & x100;
  assign n6608 = n6606 & n6607;
  assign n6609 = n6606 | n6607;
  assign n6610 = ~n6608 & n6609;
  assign n6611 = n6453 & n6610;
  assign n6612 = n6453 | n6610;
  assign n6613 = ~n6611 & n6612;
  assign n6614 = x53 & x101;
  assign n6615 = n6613 & n6614;
  assign n6616 = n6613 | n6614;
  assign n6617 = ~n6615 & n6616;
  assign n6618 = n16133 & n6617;
  assign n6619 = n16133 | n6617;
  assign n6620 = ~n6618 & n6619;
  assign n6621 = x52 & x102;
  assign n6622 = n6620 & n6621;
  assign n6623 = n6620 | n6621;
  assign n6624 = ~n6622 & n6623;
  assign n6625 = n12878 & n6624;
  assign n6626 = n12878 | n6624;
  assign n6627 = ~n6625 & n6626;
  assign n6628 = x51 & x103;
  assign n6629 = n6627 & n6628;
  assign n6630 = n6627 | n6628;
  assign n6631 = ~n6629 & n6630;
  assign n6632 = n12876 & n6631;
  assign n6633 = n12876 | n6631;
  assign n6634 = ~n6632 & n6633;
  assign n6635 = x50 & x104;
  assign n6636 = n6634 & n6635;
  assign n6637 = n6634 | n6635;
  assign n6638 = ~n6636 & n6637;
  assign n6639 = n12874 & n6638;
  assign n6640 = n12874 | n6638;
  assign n6641 = ~n6639 & n6640;
  assign n6642 = x49 & x105;
  assign n6643 = n6641 & n6642;
  assign n6644 = n6641 | n6642;
  assign n6645 = ~n6643 & n6644;
  assign n6646 = n6446 & n6645;
  assign n6647 = n6446 | n6645;
  assign n6648 = ~n6646 & n6647;
  assign n6649 = x48 & x106;
  assign n6650 = n6648 & n6649;
  assign n6651 = n6648 | n6649;
  assign n6652 = ~n6650 & n6651;
  assign n49907 = n6445 | n6642;
  assign n49908 = (n6444 & n6642) | (n6444 & n49907) | (n6642 & n49907);
  assign n16182 = (n6446 & n6641) | (n6446 & n49908) | (n6641 & n49908);
  assign n12952 = (n6643 & n6645) | (n6643 & n16182) | (n6645 & n16182);
  assign n12953 = n6636 | n12874;
  assign n12954 = (n6636 & n6638) | (n6636 & n12953) | (n6638 & n12953);
  assign n12955 = n6629 | n12876;
  assign n12956 = (n6629 & n6631) | (n6629 & n12955) | (n6631 & n12955);
  assign n12957 = n6622 | n12878;
  assign n12958 = (n6622 & n6624) | (n6622 & n12957) | (n6624 & n12957);
  assign n16183 = n6615 | n16133;
  assign n16184 = (n6615 & n6617) | (n6615 & n16183) | (n6617 & n16183);
  assign n6658 = n6608 | n6611;
  assign n12959 = n6601 | n6603;
  assign n12960 = (n6454 & n6601) | (n6454 & n12959) | (n6601 & n12959);
  assign n12961 = n6594 | n6596;
  assign n12962 = (n6594 & n12880) | (n6594 & n12961) | (n12880 & n12961);
  assign n12963 = n6587 | n6589;
  assign n12964 = (n6587 & n12882) | (n6587 & n12963) | (n12882 & n12963);
  assign n12965 = n6580 | n6582;
  assign n12966 = (n6580 & n12884) | (n6580 & n12965) | (n12884 & n12965);
  assign n12967 = n6573 | n6575;
  assign n12968 = (n6573 & n12886) | (n6573 & n12967) | (n12886 & n12967);
  assign n12969 = n6566 | n6568;
  assign n12970 = (n6566 & n12888) | (n6566 & n12969) | (n12888 & n12969);
  assign n12971 = n6559 | n6561;
  assign n12972 = (n6559 & n12890) | (n6559 & n12971) | (n12890 & n12971);
  assign n12894 = (n6348 & n12829) | (n6348 & n12893) | (n12829 & n12893);
  assign n12896 = (n6341 & n12831) | (n6341 & n12895) | (n12831 & n12895);
  assign n12982 = n6517 | n6519;
  assign n16185 = n6320 | n6517;
  assign n16186 = (n6517 & n6519) | (n6517 & n16185) | (n6519 & n16185);
  assign n16187 = (n12864 & n12982) | (n12864 & n16186) | (n12982 & n16186);
  assign n16188 = (n12863 & n12982) | (n12863 & n16186) | (n12982 & n16186);
  assign n16189 = (n16025 & n16187) | (n16025 & n16188) | (n16187 & n16188);
  assign n16190 = n6496 | n6498;
  assign n16191 = (n6496 & n12907) | (n6496 & n16190) | (n12907 & n16190);
  assign n16192 = n6299 | n6496;
  assign n16193 = (n6496 & n6498) | (n6496 & n16192) | (n6498 & n16192);
  assign n16194 = (n12840 & n16191) | (n12840 & n16193) | (n16191 & n16193);
  assign n16195 = (n16086 & n16191) | (n16086 & n16193) | (n16191 & n16193);
  assign n16196 = (n12700 & n16194) | (n12700 & n16195) | (n16194 & n16195);
  assign n12989 = n6489 | n12923;
  assign n12990 = n6489 | n12924;
  assign n16197 = (n12780 & n12989) | (n12780 & n12990) | (n12989 & n12990);
  assign n16198 = (n12781 & n12989) | (n12781 & n12990) | (n12989 & n12990);
  assign n16199 = (n12623 & n16197) | (n12623 & n16198) | (n16197 & n16198);
  assign n6678 = x75 & x80;
  assign n6679 = x74 & x81;
  assign n6680 = n6678 & n6679;
  assign n6681 = n6678 | n6679;
  assign n6682 = ~n6680 & n6681;
  assign n16200 = n6475 | n6477;
  assign n16201 = (n6475 & n12915) | (n6475 & n16200) | (n12915 & n16200);
  assign n12997 = n6682 & n16201;
  assign n16202 = n6278 | n6475;
  assign n16203 = (n6475 & n6477) | (n6475 & n16202) | (n6477 & n16202);
  assign n12998 = n6682 & n16203;
  assign n12999 = (n16089 & n12997) | (n16089 & n12998) | (n12997 & n12998);
  assign n13000 = n6682 | n16201;
  assign n13001 = n6682 | n16203;
  assign n13002 = (n16089 & n13000) | (n16089 & n13001) | (n13000 & n13001);
  assign n6685 = ~n12999 & n13002;
  assign n6686 = x73 & x82;
  assign n6687 = n6685 & n6686;
  assign n6688 = n6685 | n6686;
  assign n6689 = ~n6687 & n6688;
  assign n12992 = n6482 | n6484;
  assign n13003 = n6689 & n12992;
  assign n13004 = n6482 & n6689;
  assign n13005 = (n16148 & n13003) | (n16148 & n13004) | (n13003 & n13004);
  assign n13006 = n6689 | n12992;
  assign n13007 = n6482 | n6689;
  assign n13008 = (n16148 & n13006) | (n16148 & n13007) | (n13006 & n13007);
  assign n6692 = ~n13005 & n13008;
  assign n6693 = x72 & x83;
  assign n6694 = n6692 & n6693;
  assign n6695 = n6692 | n6693;
  assign n6696 = ~n6694 & n6695;
  assign n6697 = n16199 & n6696;
  assign n6698 = n16199 | n6696;
  assign n6699 = ~n6697 & n6698;
  assign n6700 = x71 & x84;
  assign n6701 = n6699 & n6700;
  assign n6702 = n6699 | n6700;
  assign n6703 = ~n6701 & n6702;
  assign n6704 = n16196 & n6703;
  assign n6705 = n16196 | n6703;
  assign n6706 = ~n6704 & n6705;
  assign n6707 = x70 & x85;
  assign n6708 = n6706 & n6707;
  assign n6709 = n6706 | n6707;
  assign n6710 = ~n6708 & n6709;
  assign n12984 = n6503 | n6505;
  assign n13009 = n6710 & n12984;
  assign n13010 = n6503 & n6710;
  assign n13011 = (n16143 & n13009) | (n16143 & n13010) | (n13009 & n13010);
  assign n13012 = n6710 | n12984;
  assign n13013 = n6503 | n6710;
  assign n13014 = (n16143 & n13012) | (n16143 & n13013) | (n13012 & n13013);
  assign n6713 = ~n13011 & n13014;
  assign n6714 = x69 & x86;
  assign n6715 = n6713 & n6714;
  assign n6716 = n6713 | n6714;
  assign n6717 = ~n6715 & n6716;
  assign n13015 = n6510 & n6717;
  assign n16204 = (n6717 & n12936) | (n6717 & n13015) | (n12936 & n13015);
  assign n16205 = (n6717 & n12935) | (n6717 & n13015) | (n12935 & n13015);
  assign n16206 = (n16084 & n16204) | (n16084 & n16205) | (n16204 & n16205);
  assign n13017 = n6510 | n6717;
  assign n16207 = n12936 | n13017;
  assign n16208 = n12935 | n13017;
  assign n16209 = (n16084 & n16207) | (n16084 & n16208) | (n16207 & n16208);
  assign n6720 = ~n16206 & n16209;
  assign n6721 = x68 & x87;
  assign n6722 = n6720 & n6721;
  assign n6723 = n6720 | n6721;
  assign n6724 = ~n6722 & n6723;
  assign n6725 = n16189 & n6724;
  assign n6726 = n16189 | n6724;
  assign n6727 = ~n6725 & n6726;
  assign n6728 = x67 & x88;
  assign n6729 = n6727 & n6728;
  assign n6730 = n6727 | n6728;
  assign n6731 = ~n6729 & n6730;
  assign n12979 = n6524 | n6526;
  assign n13019 = n6731 & n12979;
  assign n13020 = n6524 & n6731;
  assign n13021 = (n16138 & n13019) | (n16138 & n13020) | (n13019 & n13020);
  assign n13022 = n6731 | n12979;
  assign n13023 = n6524 | n6731;
  assign n13024 = (n16138 & n13022) | (n16138 & n13023) | (n13022 & n13023);
  assign n6734 = ~n13021 & n13024;
  assign n6735 = x66 & x89;
  assign n6736 = n6734 & n6735;
  assign n6737 = n6734 | n6735;
  assign n6738 = ~n6736 & n6737;
  assign n13025 = n6531 & n6738;
  assign n16210 = (n6738 & n12946) | (n6738 & n13025) | (n12946 & n13025);
  assign n16211 = (n6738 & n12945) | (n6738 & n13025) | (n12945 & n13025);
  assign n16212 = (n16079 & n16210) | (n16079 & n16211) | (n16210 & n16211);
  assign n13027 = n6531 | n6738;
  assign n16213 = n12946 | n13027;
  assign n16214 = n12945 | n13027;
  assign n16215 = (n16079 & n16213) | (n16079 & n16214) | (n16213 & n16214);
  assign n6741 = ~n16212 & n16215;
  assign n6742 = x65 & x90;
  assign n6743 = n6741 & n6742;
  assign n6744 = n6741 | n6742;
  assign n6745 = ~n6743 & n6744;
  assign n12977 = n6538 | n6540;
  assign n13029 = n6745 & n12977;
  assign n13030 = n6538 & n6745;
  assign n13031 = (n12896 & n13029) | (n12896 & n13030) | (n13029 & n13030);
  assign n13032 = n6745 | n12977;
  assign n13033 = n6538 | n6745;
  assign n13034 = (n12896 & n13032) | (n12896 & n13033) | (n13032 & n13033);
  assign n6748 = ~n13031 & n13034;
  assign n6749 = x64 & x91;
  assign n6750 = n6748 & n6749;
  assign n6751 = n6748 | n6749;
  assign n6752 = ~n6750 & n6751;
  assign n12975 = n6545 | n6547;
  assign n16216 = n6752 & n12975;
  assign n16217 = n6545 & n6752;
  assign n16218 = (n12894 & n16216) | (n12894 & n16217) | (n16216 & n16217);
  assign n16219 = n6752 | n12975;
  assign n16220 = n6545 | n6752;
  assign n16221 = (n12894 & n16219) | (n12894 & n16220) | (n16219 & n16220);
  assign n6755 = ~n16218 & n16221;
  assign n6756 = x63 & x92;
  assign n6757 = n6755 & n6756;
  assign n6758 = n6755 | n6756;
  assign n6759 = ~n6757 & n6758;
  assign n12973 = n6552 | n6554;
  assign n16222 = n6759 & n12973;
  assign n16223 = n6552 & n6759;
  assign n16224 = (n12892 & n16222) | (n12892 & n16223) | (n16222 & n16223);
  assign n16225 = n6759 | n12973;
  assign n16226 = n6552 | n6759;
  assign n16227 = (n12892 & n16225) | (n12892 & n16226) | (n16225 & n16226);
  assign n6762 = ~n16224 & n16227;
  assign n6763 = x62 & x93;
  assign n6764 = n6762 & n6763;
  assign n6765 = n6762 | n6763;
  assign n6766 = ~n6764 & n6765;
  assign n6767 = n12972 & n6766;
  assign n6768 = n12972 | n6766;
  assign n6769 = ~n6767 & n6768;
  assign n6770 = x61 & x94;
  assign n6771 = n6769 & n6770;
  assign n6772 = n6769 | n6770;
  assign n6773 = ~n6771 & n6772;
  assign n6774 = n12970 & n6773;
  assign n6775 = n12970 | n6773;
  assign n6776 = ~n6774 & n6775;
  assign n6777 = x60 & x95;
  assign n6778 = n6776 & n6777;
  assign n6779 = n6776 | n6777;
  assign n6780 = ~n6778 & n6779;
  assign n6781 = n12968 & n6780;
  assign n6782 = n12968 | n6780;
  assign n6783 = ~n6781 & n6782;
  assign n6784 = x59 & x96;
  assign n6785 = n6783 & n6784;
  assign n6786 = n6783 | n6784;
  assign n6787 = ~n6785 & n6786;
  assign n6788 = n12966 & n6787;
  assign n6789 = n12966 | n6787;
  assign n6790 = ~n6788 & n6789;
  assign n6791 = x58 & x97;
  assign n6792 = n6790 & n6791;
  assign n6793 = n6790 | n6791;
  assign n6794 = ~n6792 & n6793;
  assign n6795 = n12964 & n6794;
  assign n6796 = n12964 | n6794;
  assign n6797 = ~n6795 & n6796;
  assign n6798 = x57 & x98;
  assign n6799 = n6797 & n6798;
  assign n6800 = n6797 | n6798;
  assign n6801 = ~n6799 & n6800;
  assign n6802 = n12962 & n6801;
  assign n6803 = n12962 | n6801;
  assign n6804 = ~n6802 & n6803;
  assign n6805 = x56 & x99;
  assign n6806 = n6804 & n6805;
  assign n6807 = n6804 | n6805;
  assign n6808 = ~n6806 & n6807;
  assign n6809 = n12960 & n6808;
  assign n6810 = n12960 | n6808;
  assign n6811 = ~n6809 & n6810;
  assign n6812 = x55 & x100;
  assign n6813 = n6811 & n6812;
  assign n6814 = n6811 | n6812;
  assign n6815 = ~n6813 & n6814;
  assign n6816 = n6658 & n6815;
  assign n6817 = n6658 | n6815;
  assign n6818 = ~n6816 & n6817;
  assign n6819 = x54 & x101;
  assign n6820 = n6818 & n6819;
  assign n6821 = n6818 | n6819;
  assign n6822 = ~n6820 & n6821;
  assign n6823 = n16184 & n6822;
  assign n6824 = n16184 | n6822;
  assign n6825 = ~n6823 & n6824;
  assign n6826 = x53 & x102;
  assign n6827 = n6825 & n6826;
  assign n6828 = n6825 | n6826;
  assign n6829 = ~n6827 & n6828;
  assign n6830 = n12958 & n6829;
  assign n6831 = n12958 | n6829;
  assign n6832 = ~n6830 & n6831;
  assign n6833 = x52 & x103;
  assign n6834 = n6832 & n6833;
  assign n6835 = n6832 | n6833;
  assign n6836 = ~n6834 & n6835;
  assign n6837 = n12956 & n6836;
  assign n6838 = n12956 | n6836;
  assign n6839 = ~n6837 & n6838;
  assign n6840 = x51 & x104;
  assign n6841 = n6839 & n6840;
  assign n6842 = n6839 | n6840;
  assign n6843 = ~n6841 & n6842;
  assign n6844 = n12954 & n6843;
  assign n6845 = n12954 | n6843;
  assign n6846 = ~n6844 & n6845;
  assign n6847 = x50 & x105;
  assign n6848 = n6846 & n6847;
  assign n6849 = n6846 | n6847;
  assign n6850 = ~n6848 & n6849;
  assign n6851 = n12952 & n6850;
  assign n6852 = n12952 | n6850;
  assign n6853 = ~n6851 & n6852;
  assign n6854 = x49 & x106;
  assign n6855 = n6853 & n6854;
  assign n6856 = n6853 | n6854;
  assign n6857 = ~n6855 & n6856;
  assign n6858 = n6650 & n6857;
  assign n6859 = n6650 | n6857;
  assign n6860 = ~n6858 & n6859;
  assign n6861 = x48 & x107;
  assign n6862 = n6860 & n6861;
  assign n6863 = n6860 | n6861;
  assign n6864 = ~n6862 & n6863;
  assign n49909 = n6649 | n6854;
  assign n49910 = (n6648 & n6854) | (n6648 & n49909) | (n6854 & n49909);
  assign n16229 = (n6650 & n6853) | (n6650 & n49910) | (n6853 & n49910);
  assign n13036 = (n6855 & n6857) | (n6855 & n16229) | (n6857 & n16229);
  assign n13037 = n6848 | n12952;
  assign n13038 = (n6848 & n6850) | (n6848 & n13037) | (n6850 & n13037);
  assign n13039 = n6841 | n12954;
  assign n13040 = (n6841 & n6843) | (n6841 & n13039) | (n6843 & n13039);
  assign n13041 = n6834 | n12956;
  assign n13042 = (n6834 & n6836) | (n6834 & n13041) | (n6836 & n13041);
  assign n13043 = n6827 | n12958;
  assign n13044 = (n6827 & n6829) | (n6827 & n13043) | (n6829 & n13043);
  assign n16230 = n6820 | n16184;
  assign n16231 = (n6820 & n6822) | (n6820 & n16230) | (n6822 & n16230);
  assign n13045 = n6813 | n6815;
  assign n13046 = (n6658 & n6813) | (n6658 & n13045) | (n6813 & n13045);
  assign n13047 = n6806 | n6808;
  assign n13048 = (n6806 & n12960) | (n6806 & n13047) | (n12960 & n13047);
  assign n13049 = n6799 | n6801;
  assign n13050 = (n6799 & n12962) | (n6799 & n13049) | (n12962 & n13049);
  assign n13051 = n6792 | n6794;
  assign n13052 = (n6792 & n12964) | (n6792 & n13051) | (n12964 & n13051);
  assign n13053 = n6785 | n6787;
  assign n13054 = (n6785 & n12966) | (n6785 & n13053) | (n12966 & n13053);
  assign n13055 = n6778 | n6780;
  assign n13056 = (n6778 & n12968) | (n6778 & n13055) | (n12968 & n13055);
  assign n13057 = n6771 | n6773;
  assign n13058 = (n6771 & n12970) | (n6771 & n13057) | (n12970 & n13057);
  assign n12974 = (n6552 & n12892) | (n6552 & n12973) | (n12892 & n12973);
  assign n12976 = (n6545 & n12894) | (n6545 & n12975) | (n12894 & n12975);
  assign n13066 = n6736 | n6738;
  assign n16232 = n6531 | n6736;
  assign n16233 = (n6736 & n6738) | (n6736 & n16232) | (n6738 & n16232);
  assign n16234 = (n12946 & n13066) | (n12946 & n16233) | (n13066 & n16233);
  assign n16235 = (n12945 & n13066) | (n12945 & n16233) | (n13066 & n16233);
  assign n16236 = (n16079 & n16234) | (n16079 & n16235) | (n16234 & n16235);
  assign n13071 = n6715 | n6717;
  assign n16237 = n6510 | n6715;
  assign n16238 = (n6715 & n6717) | (n6715 & n16237) | (n6717 & n16237);
  assign n16239 = (n12936 & n13071) | (n12936 & n16238) | (n13071 & n16238);
  assign n16240 = (n12935 & n13071) | (n12935 & n16238) | (n13071 & n16238);
  assign n16241 = (n16084 & n16239) | (n16084 & n16240) | (n16239 & n16240);
  assign n16242 = n6503 | n6708;
  assign n16243 = (n6708 & n6710) | (n6708 & n16242) | (n6710 & n16242);
  assign n13074 = n6708 | n13009;
  assign n13075 = (n16143 & n16243) | (n16143 & n13074) | (n16243 & n13074);
  assign n6891 = x76 & x80;
  assign n6892 = x75 & x81;
  assign n6893 = n6891 & n6892;
  assign n6894 = n6891 | n6892;
  assign n6895 = ~n6893 & n6894;
  assign n16244 = n6680 | n6682;
  assign n16246 = n6895 & n16244;
  assign n16247 = n6680 & n6895;
  assign n16248 = (n16201 & n16246) | (n16201 & n16247) | (n16246 & n16247);
  assign n16249 = (n6680 & n16203) | (n6680 & n16244) | (n16203 & n16244);
  assign n13087 = n6895 & n16249;
  assign n13088 = (n16089 & n16248) | (n16089 & n13087) | (n16248 & n13087);
  assign n16250 = n6895 | n16244;
  assign n16251 = n6680 | n6895;
  assign n16252 = (n16201 & n16250) | (n16201 & n16251) | (n16250 & n16251);
  assign n13090 = n6895 | n16249;
  assign n13091 = (n16089 & n16252) | (n16089 & n13090) | (n16252 & n13090);
  assign n6898 = ~n13088 & n13091;
  assign n6899 = x74 & x82;
  assign n6900 = n6898 & n6899;
  assign n6901 = n6898 | n6899;
  assign n6902 = ~n6900 & n6901;
  assign n16253 = n6687 | n6689;
  assign n16254 = (n6687 & n12992) | (n6687 & n16253) | (n12992 & n16253);
  assign n13092 = n6902 & n16254;
  assign n16255 = n6482 | n6687;
  assign n16256 = (n6687 & n6689) | (n6687 & n16255) | (n6689 & n16255);
  assign n13093 = n6902 & n16256;
  assign n13094 = (n16148 & n13092) | (n16148 & n13093) | (n13092 & n13093);
  assign n13095 = n6902 | n16254;
  assign n13096 = n6902 | n16256;
  assign n13097 = (n16148 & n13095) | (n16148 & n13096) | (n13095 & n13096);
  assign n6905 = ~n13094 & n13097;
  assign n6906 = x73 & x83;
  assign n6907 = n6905 & n6906;
  assign n6908 = n6905 | n6906;
  assign n6909 = ~n6907 & n6908;
  assign n13078 = n6694 | n6696;
  assign n13098 = n6909 & n13078;
  assign n13099 = n6694 & n6909;
  assign n13100 = (n16199 & n13098) | (n16199 & n13099) | (n13098 & n13099);
  assign n13101 = n6909 | n13078;
  assign n13102 = n6694 | n6909;
  assign n13103 = (n16199 & n13101) | (n16199 & n13102) | (n13101 & n13102);
  assign n6912 = ~n13100 & n13103;
  assign n6913 = x72 & x84;
  assign n6914 = n6912 & n6913;
  assign n6915 = n6912 | n6913;
  assign n6916 = ~n6914 & n6915;
  assign n13076 = n6701 | n6703;
  assign n13104 = n6916 & n13076;
  assign n13105 = n6701 & n6916;
  assign n13106 = (n16196 & n13104) | (n16196 & n13105) | (n13104 & n13105);
  assign n13107 = n6916 | n13076;
  assign n13108 = n6701 | n6916;
  assign n13109 = (n16196 & n13107) | (n16196 & n13108) | (n13107 & n13108);
  assign n6919 = ~n13106 & n13109;
  assign n6920 = x71 & x85;
  assign n6921 = n6919 & n6920;
  assign n6922 = n6919 | n6920;
  assign n6923 = ~n6921 & n6922;
  assign n6924 = n13075 & n6923;
  assign n6925 = n13075 | n6923;
  assign n6926 = ~n6924 & n6925;
  assign n6927 = x70 & x86;
  assign n6928 = n6926 & n6927;
  assign n6929 = n6926 | n6927;
  assign n6930 = ~n6928 & n6929;
  assign n6931 = n16241 & n6930;
  assign n6932 = n16241 | n6930;
  assign n6933 = ~n6931 & n6932;
  assign n6934 = x69 & x87;
  assign n6935 = n6933 & n6934;
  assign n6936 = n6933 | n6934;
  assign n6937 = ~n6935 & n6936;
  assign n13068 = n6722 | n6724;
  assign n13110 = n6937 & n13068;
  assign n13111 = n6722 & n6937;
  assign n13112 = (n16189 & n13110) | (n16189 & n13111) | (n13110 & n13111);
  assign n13113 = n6937 | n13068;
  assign n13114 = n6722 | n6937;
  assign n13115 = (n16189 & n13113) | (n16189 & n13114) | (n13113 & n13114);
  assign n6940 = ~n13112 & n13115;
  assign n6941 = x68 & x88;
  assign n6942 = n6940 & n6941;
  assign n6943 = n6940 | n6941;
  assign n6944 = ~n6942 & n6943;
  assign n13116 = n6729 & n6944;
  assign n16257 = (n6944 & n13020) | (n6944 & n13116) | (n13020 & n13116);
  assign n16258 = (n6944 & n13019) | (n6944 & n13116) | (n13019 & n13116);
  assign n16259 = (n16138 & n16257) | (n16138 & n16258) | (n16257 & n16258);
  assign n13118 = n6729 | n6944;
  assign n16260 = n13020 | n13118;
  assign n16261 = n13019 | n13118;
  assign n16262 = (n16138 & n16260) | (n16138 & n16261) | (n16260 & n16261);
  assign n6947 = ~n16259 & n16262;
  assign n6948 = x67 & x89;
  assign n6949 = n6947 & n6948;
  assign n6950 = n6947 | n6948;
  assign n6951 = ~n6949 & n6950;
  assign n6952 = n16236 & n6951;
  assign n6953 = n16236 | n6951;
  assign n6954 = ~n6952 & n6953;
  assign n6955 = x66 & x90;
  assign n6956 = n6954 & n6955;
  assign n6957 = n6954 | n6955;
  assign n6958 = ~n6956 & n6957;
  assign n13120 = n6743 & n6958;
  assign n16263 = (n6958 & n13029) | (n6958 & n13120) | (n13029 & n13120);
  assign n16264 = (n6958 & n13030) | (n6958 & n13120) | (n13030 & n13120);
  assign n16265 = (n12896 & n16263) | (n12896 & n16264) | (n16263 & n16264);
  assign n13122 = n6743 | n6958;
  assign n16266 = n13029 | n13122;
  assign n16267 = n13030 | n13122;
  assign n16268 = (n12896 & n16266) | (n12896 & n16267) | (n16266 & n16267);
  assign n6961 = ~n16265 & n16268;
  assign n6962 = x65 & x91;
  assign n6963 = n6961 & n6962;
  assign n6964 = n6961 | n6962;
  assign n6965 = ~n6963 & n6964;
  assign n13063 = n6750 | n6752;
  assign n13124 = n6965 & n13063;
  assign n13125 = n6750 & n6965;
  assign n13126 = (n12976 & n13124) | (n12976 & n13125) | (n13124 & n13125);
  assign n13127 = n6965 | n13063;
  assign n13128 = n6750 | n6965;
  assign n13129 = (n12976 & n13127) | (n12976 & n13128) | (n13127 & n13128);
  assign n6968 = ~n13126 & n13129;
  assign n6969 = x64 & x92;
  assign n6970 = n6968 & n6969;
  assign n6971 = n6968 | n6969;
  assign n6972 = ~n6970 & n6971;
  assign n13061 = n6757 | n6759;
  assign n16269 = n6972 & n13061;
  assign n16270 = n6757 & n6972;
  assign n16271 = (n12974 & n16269) | (n12974 & n16270) | (n16269 & n16270);
  assign n16272 = n6972 | n13061;
  assign n16273 = n6757 | n6972;
  assign n16274 = (n12974 & n16272) | (n12974 & n16273) | (n16272 & n16273);
  assign n6975 = ~n16271 & n16274;
  assign n6976 = x63 & x93;
  assign n6977 = n6975 & n6976;
  assign n6978 = n6975 | n6976;
  assign n6979 = ~n6977 & n6978;
  assign n13059 = n6764 | n6766;
  assign n16275 = n6979 & n13059;
  assign n16276 = n6764 & n6979;
  assign n16277 = (n12972 & n16275) | (n12972 & n16276) | (n16275 & n16276);
  assign n16278 = n6979 | n13059;
  assign n16279 = n6764 | n6979;
  assign n16280 = (n12972 & n16278) | (n12972 & n16279) | (n16278 & n16279);
  assign n6982 = ~n16277 & n16280;
  assign n6983 = x62 & x94;
  assign n6984 = n6982 & n6983;
  assign n6985 = n6982 | n6983;
  assign n6986 = ~n6984 & n6985;
  assign n6987 = n13058 & n6986;
  assign n6988 = n13058 | n6986;
  assign n6989 = ~n6987 & n6988;
  assign n6990 = x61 & x95;
  assign n6991 = n6989 & n6990;
  assign n6992 = n6989 | n6990;
  assign n6993 = ~n6991 & n6992;
  assign n6994 = n13056 & n6993;
  assign n6995 = n13056 | n6993;
  assign n6996 = ~n6994 & n6995;
  assign n6997 = x60 & x96;
  assign n6998 = n6996 & n6997;
  assign n6999 = n6996 | n6997;
  assign n7000 = ~n6998 & n6999;
  assign n7001 = n13054 & n7000;
  assign n7002 = n13054 | n7000;
  assign n7003 = ~n7001 & n7002;
  assign n7004 = x59 & x97;
  assign n7005 = n7003 & n7004;
  assign n7006 = n7003 | n7004;
  assign n7007 = ~n7005 & n7006;
  assign n7008 = n13052 & n7007;
  assign n7009 = n13052 | n7007;
  assign n7010 = ~n7008 & n7009;
  assign n7011 = x58 & x98;
  assign n7012 = n7010 & n7011;
  assign n7013 = n7010 | n7011;
  assign n7014 = ~n7012 & n7013;
  assign n7015 = n13050 & n7014;
  assign n7016 = n13050 | n7014;
  assign n7017 = ~n7015 & n7016;
  assign n7018 = x57 & x99;
  assign n7019 = n7017 & n7018;
  assign n7020 = n7017 | n7018;
  assign n7021 = ~n7019 & n7020;
  assign n7022 = n13048 & n7021;
  assign n7023 = n13048 | n7021;
  assign n7024 = ~n7022 & n7023;
  assign n7025 = x56 & x100;
  assign n7026 = n7024 & n7025;
  assign n7027 = n7024 | n7025;
  assign n7028 = ~n7026 & n7027;
  assign n7029 = n13046 & n7028;
  assign n7030 = n13046 | n7028;
  assign n7031 = ~n7029 & n7030;
  assign n7032 = x55 & x101;
  assign n7033 = n7031 & n7032;
  assign n7034 = n7031 | n7032;
  assign n7035 = ~n7033 & n7034;
  assign n7036 = n16231 & n7035;
  assign n7037 = n16231 | n7035;
  assign n7038 = ~n7036 & n7037;
  assign n7039 = x54 & x102;
  assign n7040 = n7038 & n7039;
  assign n7041 = n7038 | n7039;
  assign n7042 = ~n7040 & n7041;
  assign n7043 = n13044 & n7042;
  assign n7044 = n13044 | n7042;
  assign n7045 = ~n7043 & n7044;
  assign n7046 = x53 & x103;
  assign n7047 = n7045 & n7046;
  assign n7048 = n7045 | n7046;
  assign n7049 = ~n7047 & n7048;
  assign n7050 = n13042 & n7049;
  assign n7051 = n13042 | n7049;
  assign n7052 = ~n7050 & n7051;
  assign n7053 = x52 & x104;
  assign n7054 = n7052 & n7053;
  assign n7055 = n7052 | n7053;
  assign n7056 = ~n7054 & n7055;
  assign n7057 = n13040 & n7056;
  assign n7058 = n13040 | n7056;
  assign n7059 = ~n7057 & n7058;
  assign n7060 = x51 & x105;
  assign n7061 = n7059 & n7060;
  assign n7062 = n7059 | n7060;
  assign n7063 = ~n7061 & n7062;
  assign n7064 = n13038 & n7063;
  assign n7065 = n13038 | n7063;
  assign n7066 = ~n7064 & n7065;
  assign n7067 = x50 & x106;
  assign n7068 = n7066 & n7067;
  assign n7069 = n7066 | n7067;
  assign n7070 = ~n7068 & n7069;
  assign n7071 = n13036 & n7070;
  assign n7072 = n13036 | n7070;
  assign n7073 = ~n7071 & n7072;
  assign n7074 = x49 & x107;
  assign n7075 = n7073 & n7074;
  assign n7076 = n7073 | n7074;
  assign n7077 = ~n7075 & n7076;
  assign n7078 = n6862 & n7077;
  assign n7079 = n6862 | n7077;
  assign n7080 = ~n7078 & n7079;
  assign n7081 = x48 & x108;
  assign n7082 = n7080 & n7081;
  assign n7083 = n7080 | n7081;
  assign n7084 = ~n7082 & n7083;
  assign n13130 = n6862 | n7075;
  assign n13131 = (n7075 & n7077) | (n7075 & n13130) | (n7077 & n13130);
  assign n13132 = n7068 | n13036;
  assign n13133 = (n7068 & n7070) | (n7068 & n13132) | (n7070 & n13132);
  assign n13134 = n7061 | n13038;
  assign n13135 = (n7061 & n7063) | (n7061 & n13134) | (n7063 & n13134);
  assign n13136 = n7054 | n13040;
  assign n13137 = (n7054 & n7056) | (n7054 & n13136) | (n7056 & n13136);
  assign n13138 = n7047 | n13042;
  assign n13139 = (n7047 & n7049) | (n7047 & n13138) | (n7049 & n13138);
  assign n13140 = n7040 | n13044;
  assign n13141 = (n7040 & n7042) | (n7040 & n13140) | (n7042 & n13140);
  assign n13142 = n7033 | n7035;
  assign n13143 = (n16231 & n7033) | (n16231 & n13142) | (n7033 & n13142);
  assign n13144 = n7026 | n7028;
  assign n13145 = (n7026 & n13046) | (n7026 & n13144) | (n13046 & n13144);
  assign n13146 = n7019 | n7021;
  assign n13147 = (n7019 & n13048) | (n7019 & n13146) | (n13048 & n13146);
  assign n13148 = n7012 | n7014;
  assign n13149 = (n7012 & n13050) | (n7012 & n13148) | (n13050 & n13148);
  assign n13150 = n7005 | n7007;
  assign n13151 = (n7005 & n13052) | (n7005 & n13150) | (n13052 & n13150);
  assign n13152 = n6998 | n7000;
  assign n13153 = (n6998 & n13054) | (n6998 & n13152) | (n13054 & n13152);
  assign n13154 = n6991 | n6993;
  assign n13155 = (n6991 & n13056) | (n6991 & n13154) | (n13056 & n13154);
  assign n13060 = (n6764 & n12972) | (n6764 & n13059) | (n12972 & n13059);
  assign n13062 = (n6757 & n12974) | (n6757 & n13061) | (n12974 & n13061);
  assign n13165 = n6942 | n6944;
  assign n16281 = n6729 | n6942;
  assign n16282 = (n6942 & n6944) | (n6942 & n16281) | (n6944 & n16281);
  assign n16283 = (n13020 & n13165) | (n13020 & n16282) | (n13165 & n16282);
  assign n16284 = (n13019 & n13165) | (n13019 & n16282) | (n13165 & n16282);
  assign n16285 = (n16138 & n16283) | (n16138 & n16284) | (n16283 & n16284);
  assign n7112 = x77 & x80;
  assign n7113 = x76 & x81;
  assign n7114 = n7112 & n7113;
  assign n7115 = n7112 | n7113;
  assign n7116 = ~n7114 & n7115;
  assign n16293 = n6893 & n7116;
  assign n16294 = (n7116 & n16248) | (n7116 & n16293) | (n16248 & n16293);
  assign n16295 = n6893 | n6895;
  assign n16297 = n7116 & n16295;
  assign n16298 = (n16249 & n16293) | (n16249 & n16297) | (n16293 & n16297);
  assign n13185 = (n16089 & n16294) | (n16089 & n16298) | (n16294 & n16298);
  assign n16299 = n6893 | n7116;
  assign n16300 = n16248 | n16299;
  assign n16301 = n7116 | n16295;
  assign n16302 = (n16249 & n16299) | (n16249 & n16301) | (n16299 & n16301);
  assign n13188 = (n16089 & n16300) | (n16089 & n16302) | (n16300 & n16302);
  assign n7119 = ~n13185 & n13188;
  assign n7120 = x75 & x82;
  assign n7121 = n7119 & n7120;
  assign n7122 = n7119 | n7120;
  assign n7123 = ~n7121 & n7122;
  assign n16290 = n6900 | n6902;
  assign n49911 = n7123 & n16290;
  assign n49912 = n6900 & n7123;
  assign n49913 = (n16254 & n49911) | (n16254 & n49912) | (n49911 & n49912);
  assign n16292 = (n6900 & n16256) | (n6900 & n16290) | (n16256 & n16290);
  assign n16304 = n7123 & n16292;
  assign n16305 = (n16148 & n49913) | (n16148 & n16304) | (n49913 & n16304);
  assign n49914 = n7123 | n16290;
  assign n49915 = n6900 | n7123;
  assign n49916 = (n16254 & n49914) | (n16254 & n49915) | (n49914 & n49915);
  assign n16307 = n7123 | n16292;
  assign n16308 = (n16148 & n49916) | (n16148 & n16307) | (n49916 & n16307);
  assign n7126 = ~n16305 & n16308;
  assign n7127 = x74 & x83;
  assign n7128 = n7126 & n7127;
  assign n7129 = n7126 | n7127;
  assign n7130 = ~n7128 & n7129;
  assign n16309 = n6907 | n6909;
  assign n16310 = (n6907 & n13078) | (n6907 & n16309) | (n13078 & n16309);
  assign n13189 = n7130 & n16310;
  assign n16311 = n6694 | n6907;
  assign n16312 = (n6907 & n6909) | (n6907 & n16311) | (n6909 & n16311);
  assign n13190 = n7130 & n16312;
  assign n13191 = (n16199 & n13189) | (n16199 & n13190) | (n13189 & n13190);
  assign n13192 = n7130 | n16310;
  assign n13193 = n7130 | n16312;
  assign n13194 = (n16199 & n13192) | (n16199 & n13193) | (n13192 & n13193);
  assign n7133 = ~n13191 & n13194;
  assign n7134 = x73 & x84;
  assign n7135 = n7133 & n7134;
  assign n7136 = n7133 | n7134;
  assign n7137 = ~n7135 & n7136;
  assign n16286 = n6914 | n6916;
  assign n16287 = (n6914 & n13076) | (n6914 & n16286) | (n13076 & n16286);
  assign n16313 = n7137 & n16287;
  assign n16288 = n6701 | n6914;
  assign n16289 = (n6914 & n6916) | (n6914 & n16288) | (n6916 & n16288);
  assign n16314 = n7137 & n16289;
  assign n16315 = (n16196 & n16313) | (n16196 & n16314) | (n16313 & n16314);
  assign n16316 = n7137 | n16287;
  assign n16317 = n7137 | n16289;
  assign n16318 = (n16196 & n16316) | (n16196 & n16317) | (n16316 & n16317);
  assign n7140 = ~n16315 & n16318;
  assign n7141 = x72 & x85;
  assign n7142 = n7140 & n7141;
  assign n7143 = n7140 | n7141;
  assign n7144 = ~n7142 & n7143;
  assign n13169 = n6921 | n6923;
  assign n13195 = n7144 & n13169;
  assign n13196 = n6921 & n7144;
  assign n13197 = (n13075 & n13195) | (n13075 & n13196) | (n13195 & n13196);
  assign n13198 = n7144 | n13169;
  assign n13199 = n6921 | n7144;
  assign n13200 = (n13075 & n13198) | (n13075 & n13199) | (n13198 & n13199);
  assign n7147 = ~n13197 & n13200;
  assign n7148 = x71 & x86;
  assign n7149 = n7147 & n7148;
  assign n7150 = n7147 | n7148;
  assign n7151 = ~n7149 & n7150;
  assign n13167 = n6928 | n6930;
  assign n13201 = n7151 & n13167;
  assign n13202 = n6928 & n7151;
  assign n13203 = (n16241 & n13201) | (n16241 & n13202) | (n13201 & n13202);
  assign n13204 = n7151 | n13167;
  assign n13205 = n6928 | n7151;
  assign n13206 = (n16241 & n13204) | (n16241 & n13205) | (n13204 & n13205);
  assign n7154 = ~n13203 & n13206;
  assign n7155 = x70 & x87;
  assign n7156 = n7154 & n7155;
  assign n7157 = n7154 | n7155;
  assign n7158 = ~n7156 & n7157;
  assign n13207 = n6935 & n7158;
  assign n16319 = (n7158 & n13111) | (n7158 & n13207) | (n13111 & n13207);
  assign n16320 = (n7158 & n13110) | (n7158 & n13207) | (n13110 & n13207);
  assign n16321 = (n16189 & n16319) | (n16189 & n16320) | (n16319 & n16320);
  assign n13209 = n6935 | n7158;
  assign n16322 = n13111 | n13209;
  assign n16323 = n13110 | n13209;
  assign n16324 = (n16189 & n16322) | (n16189 & n16323) | (n16322 & n16323);
  assign n7161 = ~n16321 & n16324;
  assign n7162 = x69 & x88;
  assign n7163 = n7161 & n7162;
  assign n7164 = n7161 | n7162;
  assign n7165 = ~n7163 & n7164;
  assign n7166 = n16285 & n7165;
  assign n7167 = n16285 | n7165;
  assign n7168 = ~n7166 & n7167;
  assign n7169 = x68 & x89;
  assign n7170 = n7168 & n7169;
  assign n7171 = n7168 | n7169;
  assign n7172 = ~n7170 & n7171;
  assign n13162 = n6949 | n6951;
  assign n13211 = n7172 & n13162;
  assign n13212 = n6949 & n7172;
  assign n13213 = (n16236 & n13211) | (n16236 & n13212) | (n13211 & n13212);
  assign n13214 = n7172 | n13162;
  assign n13215 = n6949 | n7172;
  assign n13216 = (n16236 & n13214) | (n16236 & n13215) | (n13214 & n13215);
  assign n7175 = ~n13213 & n13216;
  assign n7176 = x67 & x90;
  assign n7177 = n7175 & n7176;
  assign n7178 = n7175 | n7176;
  assign n7179 = ~n7177 & n7178;
  assign n13217 = n6956 & n7179;
  assign n13218 = (n7179 & n16265) | (n7179 & n13217) | (n16265 & n13217);
  assign n13219 = n6956 | n7179;
  assign n13220 = n16265 | n13219;
  assign n7182 = ~n13218 & n13220;
  assign n7183 = x66 & x91;
  assign n7184 = n7182 & n7183;
  assign n7185 = n7182 | n7183;
  assign n7186 = ~n7184 & n7185;
  assign n13221 = n6963 & n7186;
  assign n13222 = (n7186 & n13126) | (n7186 & n13221) | (n13126 & n13221);
  assign n13223 = n6963 | n7186;
  assign n13224 = n13126 | n13223;
  assign n7189 = ~n13222 & n13224;
  assign n7190 = x65 & x92;
  assign n7191 = n7189 & n7190;
  assign n7192 = n7189 | n7190;
  assign n7193 = ~n7191 & n7192;
  assign n13160 = n6970 | n6972;
  assign n13225 = n7193 & n13160;
  assign n13226 = n6970 & n7193;
  assign n13227 = (n13062 & n13225) | (n13062 & n13226) | (n13225 & n13226);
  assign n13228 = n7193 | n13160;
  assign n13229 = n6970 | n7193;
  assign n13230 = (n13062 & n13228) | (n13062 & n13229) | (n13228 & n13229);
  assign n7196 = ~n13227 & n13230;
  assign n7197 = x64 & x93;
  assign n7198 = n7196 & n7197;
  assign n7199 = n7196 | n7197;
  assign n7200 = ~n7198 & n7199;
  assign n13158 = n6977 | n6979;
  assign n16325 = n7200 & n13158;
  assign n16326 = n6977 & n7200;
  assign n16327 = (n13060 & n16325) | (n13060 & n16326) | (n16325 & n16326);
  assign n16328 = n7200 | n13158;
  assign n16329 = n6977 | n7200;
  assign n16330 = (n13060 & n16328) | (n13060 & n16329) | (n16328 & n16329);
  assign n7203 = ~n16327 & n16330;
  assign n7204 = x63 & x94;
  assign n7205 = n7203 & n7204;
  assign n7206 = n7203 | n7204;
  assign n7207 = ~n7205 & n7206;
  assign n13156 = n6984 | n6986;
  assign n16331 = n7207 & n13156;
  assign n16332 = n6984 & n7207;
  assign n16333 = (n13058 & n16331) | (n13058 & n16332) | (n16331 & n16332);
  assign n16334 = n7207 | n13156;
  assign n16335 = n6984 | n7207;
  assign n16336 = (n13058 & n16334) | (n13058 & n16335) | (n16334 & n16335);
  assign n7210 = ~n16333 & n16336;
  assign n7211 = x62 & x95;
  assign n7212 = n7210 & n7211;
  assign n7213 = n7210 | n7211;
  assign n7214 = ~n7212 & n7213;
  assign n7215 = n13155 & n7214;
  assign n7216 = n13155 | n7214;
  assign n7217 = ~n7215 & n7216;
  assign n7218 = x61 & x96;
  assign n7219 = n7217 & n7218;
  assign n7220 = n7217 | n7218;
  assign n7221 = ~n7219 & n7220;
  assign n7222 = n13153 & n7221;
  assign n7223 = n13153 | n7221;
  assign n7224 = ~n7222 & n7223;
  assign n7225 = x60 & x97;
  assign n7226 = n7224 & n7225;
  assign n7227 = n7224 | n7225;
  assign n7228 = ~n7226 & n7227;
  assign n7229 = n13151 & n7228;
  assign n7230 = n13151 | n7228;
  assign n7231 = ~n7229 & n7230;
  assign n7232 = x59 & x98;
  assign n7233 = n7231 & n7232;
  assign n7234 = n7231 | n7232;
  assign n7235 = ~n7233 & n7234;
  assign n7236 = n13149 & n7235;
  assign n7237 = n13149 | n7235;
  assign n7238 = ~n7236 & n7237;
  assign n7239 = x58 & x99;
  assign n7240 = n7238 & n7239;
  assign n7241 = n7238 | n7239;
  assign n7242 = ~n7240 & n7241;
  assign n7243 = n13147 & n7242;
  assign n7244 = n13147 | n7242;
  assign n7245 = ~n7243 & n7244;
  assign n7246 = x57 & x100;
  assign n7247 = n7245 & n7246;
  assign n7248 = n7245 | n7246;
  assign n7249 = ~n7247 & n7248;
  assign n7250 = n13145 & n7249;
  assign n7251 = n13145 | n7249;
  assign n7252 = ~n7250 & n7251;
  assign n7253 = x56 & x101;
  assign n7254 = n7252 & n7253;
  assign n7255 = n7252 | n7253;
  assign n7256 = ~n7254 & n7255;
  assign n7257 = n13143 & n7256;
  assign n7258 = n13143 | n7256;
  assign n7259 = ~n7257 & n7258;
  assign n7260 = x55 & x102;
  assign n7261 = n7259 & n7260;
  assign n7262 = n7259 | n7260;
  assign n7263 = ~n7261 & n7262;
  assign n7264 = n13141 & n7263;
  assign n7265 = n13141 | n7263;
  assign n7266 = ~n7264 & n7265;
  assign n7267 = x54 & x103;
  assign n7268 = n7266 & n7267;
  assign n7269 = n7266 | n7267;
  assign n7270 = ~n7268 & n7269;
  assign n7271 = n13139 & n7270;
  assign n7272 = n13139 | n7270;
  assign n7273 = ~n7271 & n7272;
  assign n7274 = x53 & x104;
  assign n7275 = n7273 & n7274;
  assign n7276 = n7273 | n7274;
  assign n7277 = ~n7275 & n7276;
  assign n7278 = n13137 & n7277;
  assign n7279 = n13137 | n7277;
  assign n7280 = ~n7278 & n7279;
  assign n7281 = x52 & x105;
  assign n7282 = n7280 & n7281;
  assign n7283 = n7280 | n7281;
  assign n7284 = ~n7282 & n7283;
  assign n7285 = n13135 & n7284;
  assign n7286 = n13135 | n7284;
  assign n7287 = ~n7285 & n7286;
  assign n7288 = x51 & x106;
  assign n7289 = n7287 & n7288;
  assign n7290 = n7287 | n7288;
  assign n7291 = ~n7289 & n7290;
  assign n7292 = n13133 & n7291;
  assign n7293 = n13133 | n7291;
  assign n7294 = ~n7292 & n7293;
  assign n7295 = x50 & x107;
  assign n7296 = n7294 & n7295;
  assign n7297 = n7294 | n7295;
  assign n7298 = ~n7296 & n7297;
  assign n7299 = n13131 & n7298;
  assign n7300 = n13131 | n7298;
  assign n7301 = ~n7299 & n7300;
  assign n7302 = x49 & x108;
  assign n7303 = n7301 & n7302;
  assign n7304 = n7301 | n7302;
  assign n7305 = ~n7303 & n7304;
  assign n7306 = n7082 & n7305;
  assign n7307 = n7082 | n7305;
  assign n7308 = ~n7306 & n7307;
  assign n7309 = x48 & x109;
  assign n7310 = n7308 & n7309;
  assign n7311 = n7308 | n7309;
  assign n7312 = ~n7310 & n7311;
  assign n49917 = n7081 | n7302;
  assign n49918 = (n7080 & n7302) | (n7080 & n49917) | (n7302 & n49917);
  assign n16338 = (n7082 & n7301) | (n7082 & n49918) | (n7301 & n49918);
  assign n13232 = (n7303 & n7305) | (n7303 & n16338) | (n7305 & n16338);
  assign n16339 = n7296 | n13131;
  assign n16340 = (n7296 & n7298) | (n7296 & n16339) | (n7298 & n16339);
  assign n7315 = n7289 | n7292;
  assign n7316 = n7282 | n7285;
  assign n7317 = n7275 | n7278;
  assign n7318 = n7268 | n7271;
  assign n7319 = n7261 | n7264;
  assign n13233 = n7254 | n7256;
  assign n13234 = (n7254 & n13143) | (n7254 & n13233) | (n13143 & n13233);
  assign n13235 = n7247 | n7249;
  assign n13236 = (n7247 & n13145) | (n7247 & n13235) | (n13145 & n13235);
  assign n13237 = n7240 | n7242;
  assign n13238 = (n7240 & n13147) | (n7240 & n13237) | (n13147 & n13237);
  assign n13239 = n7233 | n7235;
  assign n13240 = (n7233 & n13149) | (n7233 & n13239) | (n13149 & n13239);
  assign n13241 = n7226 | n7228;
  assign n13242 = (n7226 & n13151) | (n7226 & n13241) | (n13151 & n13241);
  assign n13243 = n7219 | n7221;
  assign n13244 = (n7219 & n13153) | (n7219 & n13243) | (n13153 & n13243);
  assign n13157 = (n6984 & n13058) | (n6984 & n13156) | (n13058 & n13156);
  assign n13159 = (n6977 & n13060) | (n6977 & n13158) | (n13060 & n13158);
  assign n13257 = n7156 | n7158;
  assign n16343 = n6935 | n7156;
  assign n16344 = (n7156 & n7158) | (n7156 & n16343) | (n7158 & n16343);
  assign n16345 = (n13111 & n13257) | (n13111 & n16344) | (n13257 & n16344);
  assign n16346 = (n13110 & n13257) | (n13110 & n16344) | (n13257 & n16344);
  assign n16347 = (n16189 & n16345) | (n16189 & n16346) | (n16345 & n16346);
  assign n7341 = x78 & x80;
  assign n7342 = x77 & x81;
  assign n7343 = n7341 & n7342;
  assign n7344 = n7341 | n7342;
  assign n7345 = ~n7343 & n7344;
  assign n49919 = n7114 & n7345;
  assign n49920 = (n7345 & n16298) | (n7345 & n49919) | (n16298 & n49919);
  assign n16353 = n7114 | n7116;
  assign n49923 = n7345 & n16353;
  assign n49921 = n6893 | n7114;
  assign n49922 = (n7114 & n7116) | (n7114 & n49921) | (n7116 & n49921);
  assign n49924 = n7345 & n49922;
  assign n49925 = (n16248 & n49923) | (n16248 & n49924) | (n49923 & n49924);
  assign n16357 = (n16089 & n49920) | (n16089 & n49925) | (n49920 & n49925);
  assign n49926 = n7114 | n7345;
  assign n49927 = n16298 | n49926;
  assign n49928 = n7345 | n16353;
  assign n49929 = n7345 | n49922;
  assign n49930 = (n16248 & n49928) | (n16248 & n49929) | (n49928 & n49929);
  assign n16360 = (n16089 & n49927) | (n16089 & n49930) | (n49927 & n49930);
  assign n7348 = ~n16357 & n16360;
  assign n7349 = x76 & x82;
  assign n7350 = n7348 & n7349;
  assign n7351 = n7348 | n7349;
  assign n7352 = ~n7350 & n7351;
  assign n13264 = n7121 | n7123;
  assign n13269 = n7352 & n13264;
  assign n13270 = n7121 & n7352;
  assign n16291 = (n6900 & n16254) | (n6900 & n16290) | (n16254 & n16290);
  assign n16361 = (n13269 & n13270) | (n13269 & n16291) | (n13270 & n16291);
  assign n16362 = (n13269 & n13270) | (n13269 & n16292) | (n13270 & n16292);
  assign n16363 = (n16148 & n16361) | (n16148 & n16362) | (n16361 & n16362);
  assign n13272 = n7352 | n13264;
  assign n13273 = n7121 | n7352;
  assign n16364 = (n13272 & n13273) | (n13272 & n16291) | (n13273 & n16291);
  assign n16365 = (n13272 & n13273) | (n13272 & n16292) | (n13273 & n16292);
  assign n16366 = (n16148 & n16364) | (n16148 & n16365) | (n16364 & n16365);
  assign n7355 = ~n16363 & n16366;
  assign n7356 = x75 & x83;
  assign n7357 = n7355 & n7356;
  assign n7358 = n7355 | n7356;
  assign n7359 = ~n7357 & n7358;
  assign n13275 = n7128 & n7359;
  assign n49931 = (n7130 & n7359) | (n7130 & n13275) | (n7359 & n13275);
  assign n49932 = n7359 & n13275;
  assign n49933 = (n16310 & n49931) | (n16310 & n49932) | (n49931 & n49932);
  assign n16368 = (n7359 & n13190) | (n7359 & n13275) | (n13190 & n13275);
  assign n16369 = (n16199 & n49933) | (n16199 & n16368) | (n49933 & n16368);
  assign n13277 = n7128 | n7359;
  assign n49934 = n7130 | n13277;
  assign n49935 = (n13277 & n16310) | (n13277 & n49934) | (n16310 & n49934);
  assign n16371 = n13190 | n13277;
  assign n16372 = (n16199 & n49935) | (n16199 & n16371) | (n49935 & n16371);
  assign n7362 = ~n16369 & n16372;
  assign n7363 = x74 & x84;
  assign n7364 = n7362 & n7363;
  assign n7365 = n7362 | n7363;
  assign n7366 = ~n7364 & n7365;
  assign n13262 = n7135 | n7137;
  assign n13279 = n7366 & n13262;
  assign n13280 = n7135 & n7366;
  assign n16373 = (n13279 & n13280) | (n13279 & n16287) | (n13280 & n16287);
  assign n16374 = (n13279 & n13280) | (n13279 & n16289) | (n13280 & n16289);
  assign n16375 = (n16196 & n16373) | (n16196 & n16374) | (n16373 & n16374);
  assign n13282 = n7366 | n13262;
  assign n13283 = n7135 | n7366;
  assign n16376 = (n13282 & n13283) | (n13282 & n16287) | (n13283 & n16287);
  assign n16377 = (n13282 & n13283) | (n13282 & n16289) | (n13283 & n16289);
  assign n16378 = (n16196 & n16376) | (n16196 & n16377) | (n16376 & n16377);
  assign n7369 = ~n16375 & n16378;
  assign n7370 = x73 & x85;
  assign n7371 = n7369 & n7370;
  assign n7372 = n7369 | n7370;
  assign n7373 = ~n7371 & n7372;
  assign n16350 = n7142 | n7144;
  assign n16351 = (n7142 & n13169) | (n7142 & n16350) | (n13169 & n16350);
  assign n16379 = n7373 & n16351;
  assign n16348 = n6921 | n7142;
  assign n16349 = (n7142 & n7144) | (n7142 & n16348) | (n7144 & n16348);
  assign n16380 = n7373 & n16349;
  assign n16381 = (n13075 & n16379) | (n13075 & n16380) | (n16379 & n16380);
  assign n16382 = n7373 | n16351;
  assign n16383 = n7373 | n16349;
  assign n16384 = (n13075 & n16382) | (n13075 & n16383) | (n16382 & n16383);
  assign n7376 = ~n16381 & n16384;
  assign n7377 = x72 & x86;
  assign n7378 = n7376 & n7377;
  assign n7379 = n7376 | n7377;
  assign n7380 = ~n7378 & n7379;
  assign n13285 = n7149 & n7380;
  assign n13286 = (n7380 & n13203) | (n7380 & n13285) | (n13203 & n13285);
  assign n13287 = n7149 | n7380;
  assign n13288 = n13203 | n13287;
  assign n7383 = ~n13286 & n13288;
  assign n7384 = x71 & x87;
  assign n7385 = n7383 & n7384;
  assign n7386 = n7383 | n7384;
  assign n7387 = ~n7385 & n7386;
  assign n7388 = n16347 & n7387;
  assign n7389 = n16347 | n7387;
  assign n7390 = ~n7388 & n7389;
  assign n7391 = x70 & x88;
  assign n7392 = n7390 & n7391;
  assign n7393 = n7390 | n7391;
  assign n7394 = ~n7392 & n7393;
  assign n13254 = n7163 | n7165;
  assign n13289 = n7394 & n13254;
  assign n13290 = n7163 & n7394;
  assign n13291 = (n16285 & n13289) | (n16285 & n13290) | (n13289 & n13290);
  assign n13292 = n7394 | n13254;
  assign n13293 = n7163 | n7394;
  assign n13294 = (n16285 & n13292) | (n16285 & n13293) | (n13292 & n13293);
  assign n7397 = ~n13291 & n13294;
  assign n7398 = x69 & x89;
  assign n7399 = n7397 & n7398;
  assign n7400 = n7397 | n7398;
  assign n7401 = ~n7399 & n7400;
  assign n13295 = n7170 & n7401;
  assign n16385 = (n7401 & n13212) | (n7401 & n13295) | (n13212 & n13295);
  assign n16386 = (n7401 & n13211) | (n7401 & n13295) | (n13211 & n13295);
  assign n16387 = (n16236 & n16385) | (n16236 & n16386) | (n16385 & n16386);
  assign n13297 = n7170 | n7401;
  assign n16388 = n13212 | n13297;
  assign n16389 = n13211 | n13297;
  assign n16390 = (n16236 & n16388) | (n16236 & n16389) | (n16388 & n16389);
  assign n7404 = ~n16387 & n16390;
  assign n7405 = x68 & x90;
  assign n7406 = n7404 & n7405;
  assign n7407 = n7404 | n7405;
  assign n7408 = ~n7406 & n7407;
  assign n13252 = n7177 | n7179;
  assign n16391 = n7408 & n13252;
  assign n16341 = n6956 | n7177;
  assign n16342 = (n7177 & n7179) | (n7177 & n16341) | (n7179 & n16341);
  assign n16392 = n7408 & n16342;
  assign n16393 = (n16265 & n16391) | (n16265 & n16392) | (n16391 & n16392);
  assign n16394 = n7408 | n13252;
  assign n16395 = n7408 | n16342;
  assign n16396 = (n16265 & n16394) | (n16265 & n16395) | (n16394 & n16395);
  assign n7411 = ~n16393 & n16396;
  assign n7412 = x67 & x91;
  assign n7413 = n7411 & n7412;
  assign n7414 = n7411 | n7412;
  assign n7415 = ~n7413 & n7414;
  assign n13299 = n7184 & n7415;
  assign n16397 = (n7415 & n13221) | (n7415 & n13299) | (n13221 & n13299);
  assign n16398 = (n7186 & n7415) | (n7186 & n13299) | (n7415 & n13299);
  assign n16399 = (n13126 & n16397) | (n13126 & n16398) | (n16397 & n16398);
  assign n13301 = n7184 | n7415;
  assign n16400 = n13221 | n13301;
  assign n16401 = n7186 | n13301;
  assign n16402 = (n13126 & n16400) | (n13126 & n16401) | (n16400 & n16401);
  assign n7418 = ~n16399 & n16402;
  assign n7419 = x66 & x92;
  assign n7420 = n7418 & n7419;
  assign n7421 = n7418 | n7419;
  assign n7422 = ~n7420 & n7421;
  assign n13303 = n7191 & n7422;
  assign n13304 = (n7422 & n13227) | (n7422 & n13303) | (n13227 & n13303);
  assign n13305 = n7191 | n7422;
  assign n13306 = n13227 | n13305;
  assign n7425 = ~n13304 & n13306;
  assign n7426 = x65 & x93;
  assign n7427 = n7425 & n7426;
  assign n7428 = n7425 | n7426;
  assign n7429 = ~n7427 & n7428;
  assign n13249 = n7198 | n7200;
  assign n13307 = n7429 & n13249;
  assign n13308 = n7198 & n7429;
  assign n13309 = (n13159 & n13307) | (n13159 & n13308) | (n13307 & n13308);
  assign n13310 = n7429 | n13249;
  assign n13311 = n7198 | n7429;
  assign n13312 = (n13159 & n13310) | (n13159 & n13311) | (n13310 & n13311);
  assign n7432 = ~n13309 & n13312;
  assign n7433 = x64 & x94;
  assign n7434 = n7432 & n7433;
  assign n7435 = n7432 | n7433;
  assign n7436 = ~n7434 & n7435;
  assign n13247 = n7205 | n7207;
  assign n16403 = n7436 & n13247;
  assign n16404 = n7205 & n7436;
  assign n16405 = (n13157 & n16403) | (n13157 & n16404) | (n16403 & n16404);
  assign n16406 = n7436 | n13247;
  assign n16407 = n7205 | n7436;
  assign n16408 = (n13157 & n16406) | (n13157 & n16407) | (n16406 & n16407);
  assign n7439 = ~n16405 & n16408;
  assign n7440 = x63 & x95;
  assign n7441 = n7439 & n7440;
  assign n7442 = n7439 | n7440;
  assign n7443 = ~n7441 & n7442;
  assign n13245 = n7212 | n7214;
  assign n16409 = n7443 & n13245;
  assign n16410 = n7212 & n7443;
  assign n16411 = (n13155 & n16409) | (n13155 & n16410) | (n16409 & n16410);
  assign n16412 = n7443 | n13245;
  assign n16413 = n7212 | n7443;
  assign n16414 = (n13155 & n16412) | (n13155 & n16413) | (n16412 & n16413);
  assign n7446 = ~n16411 & n16414;
  assign n7447 = x62 & x96;
  assign n7448 = n7446 & n7447;
  assign n7449 = n7446 | n7447;
  assign n7450 = ~n7448 & n7449;
  assign n7451 = n13244 & n7450;
  assign n7452 = n13244 | n7450;
  assign n7453 = ~n7451 & n7452;
  assign n7454 = x61 & x97;
  assign n7455 = n7453 & n7454;
  assign n7456 = n7453 | n7454;
  assign n7457 = ~n7455 & n7456;
  assign n7458 = n13242 & n7457;
  assign n7459 = n13242 | n7457;
  assign n7460 = ~n7458 & n7459;
  assign n7461 = x60 & x98;
  assign n7462 = n7460 & n7461;
  assign n7463 = n7460 | n7461;
  assign n7464 = ~n7462 & n7463;
  assign n7465 = n13240 & n7464;
  assign n7466 = n13240 | n7464;
  assign n7467 = ~n7465 & n7466;
  assign n7468 = x59 & x99;
  assign n7469 = n7467 & n7468;
  assign n7470 = n7467 | n7468;
  assign n7471 = ~n7469 & n7470;
  assign n7472 = n13238 & n7471;
  assign n7473 = n13238 | n7471;
  assign n7474 = ~n7472 & n7473;
  assign n7475 = x58 & x100;
  assign n7476 = n7474 & n7475;
  assign n7477 = n7474 | n7475;
  assign n7478 = ~n7476 & n7477;
  assign n7479 = n13236 & n7478;
  assign n7480 = n13236 | n7478;
  assign n7481 = ~n7479 & n7480;
  assign n7482 = x57 & x101;
  assign n7483 = n7481 & n7482;
  assign n7484 = n7481 | n7482;
  assign n7485 = ~n7483 & n7484;
  assign n7486 = n13234 & n7485;
  assign n7487 = n13234 | n7485;
  assign n7488 = ~n7486 & n7487;
  assign n7489 = x56 & x102;
  assign n7490 = n7488 & n7489;
  assign n7491 = n7488 | n7489;
  assign n7492 = ~n7490 & n7491;
  assign n7493 = n7319 & n7492;
  assign n7494 = n7319 | n7492;
  assign n7495 = ~n7493 & n7494;
  assign n7496 = x55 & x103;
  assign n7497 = n7495 & n7496;
  assign n7498 = n7495 | n7496;
  assign n7499 = ~n7497 & n7498;
  assign n7500 = n7318 & n7499;
  assign n7501 = n7318 | n7499;
  assign n7502 = ~n7500 & n7501;
  assign n7503 = x54 & x104;
  assign n7504 = n7502 & n7503;
  assign n7505 = n7502 | n7503;
  assign n7506 = ~n7504 & n7505;
  assign n7507 = n7317 & n7506;
  assign n7508 = n7317 | n7506;
  assign n7509 = ~n7507 & n7508;
  assign n7510 = x53 & x105;
  assign n7511 = n7509 & n7510;
  assign n7512 = n7509 | n7510;
  assign n7513 = ~n7511 & n7512;
  assign n7514 = n7316 & n7513;
  assign n7515 = n7316 | n7513;
  assign n7516 = ~n7514 & n7515;
  assign n7517 = x52 & x106;
  assign n7518 = n7516 & n7517;
  assign n7519 = n7516 | n7517;
  assign n7520 = ~n7518 & n7519;
  assign n7521 = n7315 & n7520;
  assign n7522 = n7315 | n7520;
  assign n7523 = ~n7521 & n7522;
  assign n7524 = x51 & x107;
  assign n7525 = n7523 & n7524;
  assign n7526 = n7523 | n7524;
  assign n7527 = ~n7525 & n7526;
  assign n7528 = n16340 & n7527;
  assign n7529 = n16340 | n7527;
  assign n7530 = ~n7528 & n7529;
  assign n7531 = x50 & x108;
  assign n7532 = n7530 & n7531;
  assign n7533 = n7530 | n7531;
  assign n7534 = ~n7532 & n7533;
  assign n7535 = n13232 & n7534;
  assign n7536 = n13232 | n7534;
  assign n7537 = ~n7535 & n7536;
  assign n7538 = x49 & x109;
  assign n7539 = n7537 & n7538;
  assign n7540 = n7537 | n7538;
  assign n7541 = ~n7539 & n7540;
  assign n7542 = n7310 & n7541;
  assign n7543 = n7310 | n7541;
  assign n7544 = ~n7542 & n7543;
  assign n7545 = x48 & x110;
  assign n7546 = n7544 & n7545;
  assign n7547 = n7544 | n7545;
  assign n7548 = ~n7546 & n7547;
  assign n49936 = n7309 | n7538;
  assign n49937 = (n7308 & n7538) | (n7308 & n49936) | (n7538 & n49936);
  assign n16416 = (n7310 & n7537) | (n7310 & n49937) | (n7537 & n49937);
  assign n13314 = (n7539 & n7541) | (n7539 & n16416) | (n7541 & n16416);
  assign n13315 = n7532 | n13232;
  assign n13316 = (n7532 & n7534) | (n7532 & n13315) | (n7534 & n13315);
  assign n16417 = n7525 | n16340;
  assign n16418 = (n7525 & n7527) | (n7525 & n16417) | (n7527 & n16417);
  assign n7552 = n7518 | n7521;
  assign n7553 = n7511 | n7514;
  assign n7554 = n7504 | n7507;
  assign n7555 = n7497 | n7500;
  assign n13317 = n7490 | n7492;
  assign n13318 = (n7319 & n7490) | (n7319 & n13317) | (n7490 & n13317);
  assign n13319 = n7483 | n7485;
  assign n13320 = (n7483 & n13234) | (n7483 & n13319) | (n13234 & n13319);
  assign n13321 = n7476 | n7478;
  assign n13322 = (n7476 & n13236) | (n7476 & n13321) | (n13236 & n13321);
  assign n13323 = n7469 | n7471;
  assign n13324 = (n7469 & n13238) | (n7469 & n13323) | (n13238 & n13323);
  assign n13325 = n7462 | n7464;
  assign n13326 = (n7462 & n13240) | (n7462 & n13325) | (n13240 & n13325);
  assign n13327 = n7455 | n7457;
  assign n13328 = (n7455 & n13242) | (n7455 & n13327) | (n13242 & n13327);
  assign n13246 = (n7212 & n13155) | (n7212 & n13245) | (n13155 & n13245);
  assign n13248 = (n7205 & n13157) | (n7205 & n13247) | (n13157 & n13247);
  assign n13338 = n7399 | n7401;
  assign n16419 = n7170 | n7399;
  assign n16420 = (n7399 & n7401) | (n7399 & n16419) | (n7401 & n16419);
  assign n16421 = (n13212 & n13338) | (n13212 & n16420) | (n13338 & n16420);
  assign n16422 = (n13211 & n13338) | (n13211 & n16420) | (n13338 & n16420);
  assign n16423 = (n16236 & n16421) | (n16236 & n16422) | (n16421 & n16422);
  assign n13173 = (n16196 & n16287) | (n16196 & n16289) | (n16287 & n16289);
  assign n7578 = x79 & x80;
  assign n7579 = x78 & x81;
  assign n7580 = n7578 & n7579;
  assign n7581 = n7578 | n7579;
  assign n7582 = ~n7580 & n7581;
  assign n13356 = n7343 | n7345;
  assign n13358 = n7582 & n13356;
  assign n13359 = n7343 & n7582;
  assign n49938 = (n7114 & n13358) | (n7114 & n13359) | (n13358 & n13359);
  assign n49939 = n13358 | n13359;
  assign n49940 = (n16298 & n49938) | (n16298 & n49939) | (n49938 & n49939);
  assign n49941 = (n13358 & n13359) | (n13358 & n16353) | (n13359 & n16353);
  assign n49942 = (n13358 & n13359) | (n13358 & n49922) | (n13359 & n49922);
  assign n49943 = (n16248 & n49941) | (n16248 & n49942) | (n49941 & n49942);
  assign n16428 = (n16089 & n49940) | (n16089 & n49943) | (n49940 & n49943);
  assign n13361 = n7582 | n13356;
  assign n13362 = n7343 | n7582;
  assign n49944 = (n7114 & n13361) | (n7114 & n13362) | (n13361 & n13362);
  assign n49945 = n13361 | n13362;
  assign n49946 = (n16298 & n49944) | (n16298 & n49945) | (n49944 & n49945);
  assign n49947 = (n13361 & n13362) | (n13361 & n16353) | (n13362 & n16353);
  assign n49948 = (n13361 & n13362) | (n13361 & n49922) | (n13362 & n49922);
  assign n49949 = (n16248 & n49947) | (n16248 & n49948) | (n49947 & n49948);
  assign n16431 = (n16089 & n49946) | (n16089 & n49949) | (n49946 & n49949);
  assign n7585 = ~n16428 & n16431;
  assign n7586 = x77 & x82;
  assign n7587 = n7585 & n7586;
  assign n7588 = n7585 | n7586;
  assign n7589 = ~n7587 & n7588;
  assign n16432 = n7350 | n7352;
  assign n16433 = (n7350 & n13264) | (n7350 & n16432) | (n13264 & n16432);
  assign n13364 = n7589 & n16433;
  assign n16434 = n7121 | n7350;
  assign n16435 = (n7350 & n7352) | (n7350 & n16434) | (n7352 & n16434);
  assign n13365 = n7589 & n16435;
  assign n16436 = (n13364 & n13365) | (n13364 & n16291) | (n13365 & n16291);
  assign n16437 = (n13364 & n13365) | (n13364 & n16292) | (n13365 & n16292);
  assign n16438 = (n16148 & n16436) | (n16148 & n16437) | (n16436 & n16437);
  assign n13367 = n7589 | n16433;
  assign n13368 = n7589 | n16435;
  assign n16439 = (n13367 & n13368) | (n13367 & n16291) | (n13368 & n16291);
  assign n16440 = (n13367 & n13368) | (n13367 & n16292) | (n13368 & n16292);
  assign n16441 = (n16148 & n16439) | (n16148 & n16440) | (n16439 & n16440);
  assign n7592 = ~n16438 & n16441;
  assign n7593 = x76 & x83;
  assign n7594 = n7592 & n7593;
  assign n7595 = n7592 | n7593;
  assign n7596 = ~n7594 & n7595;
  assign n16442 = n7128 | n7357;
  assign n16443 = (n7357 & n7359) | (n7357 & n16442) | (n7359 & n16442);
  assign n13370 = n7596 & n16443;
  assign n13351 = n7357 | n7359;
  assign n13371 = n7596 & n13351;
  assign n16444 = (n13189 & n13370) | (n13189 & n13371) | (n13370 & n13371);
  assign n16445 = (n13190 & n13370) | (n13190 & n13371) | (n13370 & n13371);
  assign n16446 = (n16199 & n16444) | (n16199 & n16445) | (n16444 & n16445);
  assign n13373 = n7596 | n16443;
  assign n13374 = n7596 | n13351;
  assign n16447 = (n13189 & n13373) | (n13189 & n13374) | (n13373 & n13374);
  assign n16448 = (n13190 & n13373) | (n13190 & n13374) | (n13373 & n13374);
  assign n16449 = (n16199 & n16447) | (n16199 & n16448) | (n16447 & n16448);
  assign n7599 = ~n16446 & n16449;
  assign n7600 = x75 & x84;
  assign n7601 = n7599 & n7600;
  assign n7602 = n7599 | n7600;
  assign n7603 = ~n7601 & n7602;
  assign n16450 = n7364 | n7366;
  assign n16451 = (n7364 & n13262) | (n7364 & n16450) | (n13262 & n16450);
  assign n13376 = n7603 & n16451;
  assign n16452 = n7135 | n7364;
  assign n16453 = (n7364 & n7366) | (n7364 & n16452) | (n7366 & n16452);
  assign n13377 = n7603 & n16453;
  assign n13378 = (n13173 & n13376) | (n13173 & n13377) | (n13376 & n13377);
  assign n13379 = n7603 | n16451;
  assign n13380 = n7603 | n16453;
  assign n13381 = (n13173 & n13379) | (n13173 & n13380) | (n13379 & n13380);
  assign n7606 = ~n13378 & n13381;
  assign n7607 = x74 & x85;
  assign n7608 = n7606 & n7607;
  assign n7609 = n7606 | n7607;
  assign n7610 = ~n7608 & n7609;
  assign n13345 = n7371 | n7373;
  assign n13382 = n7610 & n13345;
  assign n13383 = n7371 & n7610;
  assign n16454 = (n13382 & n13383) | (n13382 & n16351) | (n13383 & n16351);
  assign n16455 = (n13382 & n13383) | (n13382 & n16349) | (n13383 & n16349);
  assign n16456 = (n13075 & n16454) | (n13075 & n16455) | (n16454 & n16455);
  assign n13385 = n7610 | n13345;
  assign n13386 = n7371 | n7610;
  assign n16457 = (n13385 & n13386) | (n13385 & n16351) | (n13386 & n16351);
  assign n16458 = (n13385 & n13386) | (n13385 & n16349) | (n13386 & n16349);
  assign n16459 = (n13075 & n16457) | (n13075 & n16458) | (n16457 & n16458);
  assign n7613 = ~n16456 & n16459;
  assign n7614 = x73 & x86;
  assign n7615 = n7613 & n7614;
  assign n7616 = n7613 | n7614;
  assign n7617 = ~n7615 & n7616;
  assign n13343 = n7378 | n7380;
  assign n16460 = n7617 & n13343;
  assign n16424 = n7149 | n7378;
  assign n16425 = (n7378 & n7380) | (n7378 & n16424) | (n7380 & n16424);
  assign n16461 = n7617 & n16425;
  assign n16462 = (n13203 & n16460) | (n13203 & n16461) | (n16460 & n16461);
  assign n16463 = n7617 | n13343;
  assign n16464 = n7617 | n16425;
  assign n16465 = (n13203 & n16463) | (n13203 & n16464) | (n16463 & n16464);
  assign n7620 = ~n16462 & n16465;
  assign n7621 = x72 & x87;
  assign n7622 = n7620 & n7621;
  assign n7623 = n7620 | n7621;
  assign n7624 = ~n7622 & n7623;
  assign n13340 = n7385 | n7387;
  assign n13388 = n7624 & n13340;
  assign n13389 = n7385 & n7624;
  assign n13390 = (n16347 & n13388) | (n16347 & n13389) | (n13388 & n13389);
  assign n13391 = n7624 | n13340;
  assign n13392 = n7385 | n7624;
  assign n13393 = (n16347 & n13391) | (n16347 & n13392) | (n13391 & n13392);
  assign n7627 = ~n13390 & n13393;
  assign n7628 = x71 & x88;
  assign n7629 = n7627 & n7628;
  assign n7630 = n7627 | n7628;
  assign n7631 = ~n7629 & n7630;
  assign n13394 = n7392 & n7631;
  assign n16466 = (n7631 & n13290) | (n7631 & n13394) | (n13290 & n13394);
  assign n16467 = (n7631 & n13289) | (n7631 & n13394) | (n13289 & n13394);
  assign n16468 = (n16285 & n16466) | (n16285 & n16467) | (n16466 & n16467);
  assign n13396 = n7392 | n7631;
  assign n16469 = n13290 | n13396;
  assign n16470 = n13289 | n13396;
  assign n16471 = (n16285 & n16469) | (n16285 & n16470) | (n16469 & n16470);
  assign n7634 = ~n16468 & n16471;
  assign n7635 = x70 & x89;
  assign n7636 = n7634 & n7635;
  assign n7637 = n7634 | n7635;
  assign n7638 = ~n7636 & n7637;
  assign n7639 = n16423 & n7638;
  assign n7640 = n16423 | n7638;
  assign n7641 = ~n7639 & n7640;
  assign n7642 = x69 & x90;
  assign n7643 = n7641 & n7642;
  assign n7644 = n7641 | n7642;
  assign n7645 = ~n7643 & n7644;
  assign n13335 = n7406 | n7408;
  assign n13398 = n7645 & n13335;
  assign n13399 = n7406 & n7645;
  assign n16472 = (n13252 & n13398) | (n13252 & n13399) | (n13398 & n13399);
  assign n16473 = (n13398 & n13399) | (n13398 & n16342) | (n13399 & n16342);
  assign n16474 = (n16265 & n16472) | (n16265 & n16473) | (n16472 & n16473);
  assign n13401 = n7645 | n13335;
  assign n13402 = n7406 | n7645;
  assign n16475 = (n13252 & n13401) | (n13252 & n13402) | (n13401 & n13402);
  assign n16476 = (n13401 & n13402) | (n13401 & n16342) | (n13402 & n16342);
  assign n16477 = (n16265 & n16475) | (n16265 & n16476) | (n16475 & n16476);
  assign n7648 = ~n16474 & n16477;
  assign n7649 = x68 & x91;
  assign n7650 = n7648 & n7649;
  assign n7651 = n7648 | n7649;
  assign n7652 = ~n7650 & n7651;
  assign n13404 = n7413 & n7652;
  assign n13405 = (n7652 & n16399) | (n7652 & n13404) | (n16399 & n13404);
  assign n13406 = n7413 | n7652;
  assign n13407 = n16399 | n13406;
  assign n7655 = ~n13405 & n13407;
  assign n7656 = x67 & x92;
  assign n7657 = n7655 & n7656;
  assign n7658 = n7655 | n7656;
  assign n7659 = ~n7657 & n7658;
  assign n13408 = n7420 & n7659;
  assign n13409 = (n7659 & n13304) | (n7659 & n13408) | (n13304 & n13408);
  assign n13410 = n7420 | n7659;
  assign n13411 = n13304 | n13410;
  assign n7662 = ~n13409 & n13411;
  assign n7663 = x66 & x93;
  assign n7664 = n7662 & n7663;
  assign n7665 = n7662 | n7663;
  assign n7666 = ~n7664 & n7665;
  assign n13412 = n7427 & n7666;
  assign n13413 = (n7666 & n13309) | (n7666 & n13412) | (n13309 & n13412);
  assign n13414 = n7427 | n7666;
  assign n13415 = n13309 | n13414;
  assign n7669 = ~n13413 & n13415;
  assign n7670 = x65 & x94;
  assign n7671 = n7669 & n7670;
  assign n7672 = n7669 | n7670;
  assign n7673 = ~n7671 & n7672;
  assign n13333 = n7434 | n7436;
  assign n13416 = n7673 & n13333;
  assign n13417 = n7434 & n7673;
  assign n13418 = (n13248 & n13416) | (n13248 & n13417) | (n13416 & n13417);
  assign n13419 = n7673 | n13333;
  assign n13420 = n7434 | n7673;
  assign n13421 = (n13248 & n13419) | (n13248 & n13420) | (n13419 & n13420);
  assign n7676 = ~n13418 & n13421;
  assign n7677 = x64 & x95;
  assign n7678 = n7676 & n7677;
  assign n7679 = n7676 | n7677;
  assign n7680 = ~n7678 & n7679;
  assign n13331 = n7441 | n7443;
  assign n16478 = n7680 & n13331;
  assign n16479 = n7441 & n7680;
  assign n16480 = (n13246 & n16478) | (n13246 & n16479) | (n16478 & n16479);
  assign n16481 = n7680 | n13331;
  assign n16482 = n7441 | n7680;
  assign n16483 = (n13246 & n16481) | (n13246 & n16482) | (n16481 & n16482);
  assign n7683 = ~n16480 & n16483;
  assign n7684 = x63 & x96;
  assign n7685 = n7683 & n7684;
  assign n7686 = n7683 | n7684;
  assign n7687 = ~n7685 & n7686;
  assign n13329 = n7448 | n7450;
  assign n16484 = n7687 & n13329;
  assign n16485 = n7448 & n7687;
  assign n16486 = (n13244 & n16484) | (n13244 & n16485) | (n16484 & n16485);
  assign n16487 = n7687 | n13329;
  assign n16488 = n7448 | n7687;
  assign n16489 = (n13244 & n16487) | (n13244 & n16488) | (n16487 & n16488);
  assign n7690 = ~n16486 & n16489;
  assign n7691 = x62 & x97;
  assign n7692 = n7690 & n7691;
  assign n7693 = n7690 | n7691;
  assign n7694 = ~n7692 & n7693;
  assign n7695 = n13328 & n7694;
  assign n7696 = n13328 | n7694;
  assign n7697 = ~n7695 & n7696;
  assign n7698 = x61 & x98;
  assign n7699 = n7697 & n7698;
  assign n7700 = n7697 | n7698;
  assign n7701 = ~n7699 & n7700;
  assign n7702 = n13326 & n7701;
  assign n7703 = n13326 | n7701;
  assign n7704 = ~n7702 & n7703;
  assign n7705 = x60 & x99;
  assign n7706 = n7704 & n7705;
  assign n7707 = n7704 | n7705;
  assign n7708 = ~n7706 & n7707;
  assign n7709 = n13324 & n7708;
  assign n7710 = n13324 | n7708;
  assign n7711 = ~n7709 & n7710;
  assign n7712 = x59 & x100;
  assign n7713 = n7711 & n7712;
  assign n7714 = n7711 | n7712;
  assign n7715 = ~n7713 & n7714;
  assign n7716 = n13322 & n7715;
  assign n7717 = n13322 | n7715;
  assign n7718 = ~n7716 & n7717;
  assign n7719 = x58 & x101;
  assign n7720 = n7718 & n7719;
  assign n7721 = n7718 | n7719;
  assign n7722 = ~n7720 & n7721;
  assign n7723 = n13320 & n7722;
  assign n7724 = n13320 | n7722;
  assign n7725 = ~n7723 & n7724;
  assign n7726 = x57 & x102;
  assign n7727 = n7725 & n7726;
  assign n7728 = n7725 | n7726;
  assign n7729 = ~n7727 & n7728;
  assign n7730 = n13318 & n7729;
  assign n7731 = n13318 | n7729;
  assign n7732 = ~n7730 & n7731;
  assign n7733 = x56 & x103;
  assign n7734 = n7732 & n7733;
  assign n7735 = n7732 | n7733;
  assign n7736 = ~n7734 & n7735;
  assign n7737 = n7555 & n7736;
  assign n7738 = n7555 | n7736;
  assign n7739 = ~n7737 & n7738;
  assign n7740 = x55 & x104;
  assign n7741 = n7739 & n7740;
  assign n7742 = n7739 | n7740;
  assign n7743 = ~n7741 & n7742;
  assign n7744 = n7554 & n7743;
  assign n7745 = n7554 | n7743;
  assign n7746 = ~n7744 & n7745;
  assign n7747 = x54 & x105;
  assign n7748 = n7746 & n7747;
  assign n7749 = n7746 | n7747;
  assign n7750 = ~n7748 & n7749;
  assign n7751 = n7553 & n7750;
  assign n7752 = n7553 | n7750;
  assign n7753 = ~n7751 & n7752;
  assign n7754 = x53 & x106;
  assign n7755 = n7753 & n7754;
  assign n7756 = n7753 | n7754;
  assign n7757 = ~n7755 & n7756;
  assign n7758 = n7552 & n7757;
  assign n7759 = n7552 | n7757;
  assign n7760 = ~n7758 & n7759;
  assign n7761 = x52 & x107;
  assign n7762 = n7760 & n7761;
  assign n7763 = n7760 | n7761;
  assign n7764 = ~n7762 & n7763;
  assign n7765 = n16418 & n7764;
  assign n7766 = n16418 | n7764;
  assign n7767 = ~n7765 & n7766;
  assign n7768 = x51 & x108;
  assign n7769 = n7767 & n7768;
  assign n7770 = n7767 | n7768;
  assign n7771 = ~n7769 & n7770;
  assign n7772 = n13316 & n7771;
  assign n7773 = n13316 | n7771;
  assign n7774 = ~n7772 & n7773;
  assign n7775 = x50 & x109;
  assign n7776 = n7774 & n7775;
  assign n7777 = n7774 | n7775;
  assign n7778 = ~n7776 & n7777;
  assign n7779 = n13314 & n7778;
  assign n7780 = n13314 | n7778;
  assign n7781 = ~n7779 & n7780;
  assign n7782 = x49 & x110;
  assign n7783 = n7781 & n7782;
  assign n7784 = n7781 | n7782;
  assign n7785 = ~n7783 & n7784;
  assign n7786 = n7546 & n7785;
  assign n7787 = n7546 | n7785;
  assign n7788 = ~n7786 & n7787;
  assign n7789 = x48 & x111;
  assign n7790 = n7788 & n7789;
  assign n7791 = n7788 | n7789;
  assign n7792 = ~n7790 & n7791;
  assign n49950 = n7545 | n7782;
  assign n49951 = (n7544 & n7782) | (n7544 & n49950) | (n7782 & n49950);
  assign n16491 = (n7546 & n7781) | (n7546 & n49951) | (n7781 & n49951);
  assign n13423 = (n7783 & n7785) | (n7783 & n16491) | (n7785 & n16491);
  assign n13424 = n7776 | n13314;
  assign n13425 = (n7776 & n7778) | (n7776 & n13424) | (n7778 & n13424);
  assign n13426 = n7769 | n13316;
  assign n13427 = (n7769 & n7771) | (n7769 & n13426) | (n7771 & n13426);
  assign n16492 = n7762 | n16418;
  assign n16493 = (n7762 & n7764) | (n7762 & n16492) | (n7764 & n16492);
  assign n7797 = n7755 | n7758;
  assign n7798 = n7748 | n7751;
  assign n7799 = n7741 | n7744;
  assign n13428 = n7734 | n7736;
  assign n13429 = (n7555 & n7734) | (n7555 & n13428) | (n7734 & n13428);
  assign n13430 = n7727 | n7729;
  assign n13431 = (n7727 & n13318) | (n7727 & n13430) | (n13318 & n13430);
  assign n13432 = n7720 | n7722;
  assign n13433 = (n7720 & n13320) | (n7720 & n13432) | (n13320 & n13432);
  assign n13434 = n7713 | n7715;
  assign n13435 = (n7713 & n13322) | (n7713 & n13434) | (n13322 & n13434);
  assign n13436 = n7706 | n7708;
  assign n13437 = (n7706 & n13324) | (n7706 & n13436) | (n13324 & n13436);
  assign n13438 = n7699 | n7701;
  assign n13439 = (n7699 & n13326) | (n7699 & n13438) | (n13326 & n13438);
  assign n13330 = (n7448 & n13244) | (n7448 & n13329) | (n13244 & n13329);
  assign n13332 = (n7441 & n13246) | (n7441 & n13331) | (n13246 & n13331);
  assign n13452 = n7629 | n7631;
  assign n16496 = n7392 | n7629;
  assign n16497 = (n7629 & n7631) | (n7629 & n16496) | (n7631 & n16496);
  assign n16498 = (n13290 & n13452) | (n13290 & n16497) | (n13452 & n16497);
  assign n16499 = (n13289 & n13452) | (n13289 & n16497) | (n13452 & n16497);
  assign n16500 = (n16285 & n16498) | (n16285 & n16499) | (n16498 & n16499);
  assign n13261 = (n13075 & n16349) | (n13075 & n16351) | (n16349 & n16351);
  assign n16503 = n7594 | n7596;
  assign n16504 = (n7594 & n16443) | (n7594 & n16503) | (n16443 & n16503);
  assign n16505 = (n7594 & n13351) | (n7594 & n16503) | (n13351 & n16503);
  assign n16506 = (n13189 & n16504) | (n13189 & n16505) | (n16504 & n16505);
  assign n16507 = (n13190 & n16504) | (n13190 & n16505) | (n16504 & n16505);
  assign n16508 = (n16199 & n16506) | (n16199 & n16507) | (n16506 & n16507);
  assign n13267 = n7114 | n16298;
  assign n7823 = x79 & x81;
  assign n16509 = n7580 | n7582;
  assign n16510 = (n7580 & n13356) | (n7580 & n16509) | (n13356 & n16509);
  assign n13468 = n7823 & n16510;
  assign n16511 = n7343 | n7580;
  assign n16512 = (n7580 & n7582) | (n7580 & n16511) | (n7582 & n16511);
  assign n13469 = n7823 & n16512;
  assign n16513 = (n13267 & n13468) | (n13267 & n13469) | (n13468 & n13469);
  assign n16354 = (n16248 & n49922) | (n16248 & n16353) | (n49922 & n16353);
  assign n16514 = (n13468 & n13469) | (n13468 & n16354) | (n13469 & n16354);
  assign n16515 = (n16089 & n16513) | (n16089 & n16514) | (n16513 & n16514);
  assign n13471 = n7823 | n16510;
  assign n13472 = n7823 | n16512;
  assign n16516 = (n13267 & n13471) | (n13267 & n13472) | (n13471 & n13472);
  assign n16517 = (n13471 & n13472) | (n13471 & n16354) | (n13472 & n16354);
  assign n16518 = (n16089 & n16516) | (n16089 & n16517) | (n16516 & n16517);
  assign n7826 = ~n16515 & n16518;
  assign n7827 = x78 & x82;
  assign n7828 = n7826 & n7827;
  assign n7829 = n7826 | n7827;
  assign n7830 = ~n7828 & n7829;
  assign n16519 = n7587 | n7589;
  assign n16524 = (n7587 & n16435) | (n7587 & n16519) | (n16435 & n16519);
  assign n13475 = n7830 & n16524;
  assign n16521 = n7830 & n16519;
  assign n16522 = n7587 & n7830;
  assign n16523 = (n16433 & n16521) | (n16433 & n16522) | (n16521 & n16522);
  assign n16525 = (n13475 & n16291) | (n13475 & n16523) | (n16291 & n16523);
  assign n16526 = (n13475 & n16292) | (n13475 & n16523) | (n16292 & n16523);
  assign n16527 = (n16148 & n16525) | (n16148 & n16526) | (n16525 & n16526);
  assign n13478 = n7830 | n16524;
  assign n16528 = n7830 | n16519;
  assign n16529 = n7587 | n7830;
  assign n16530 = (n16433 & n16528) | (n16433 & n16529) | (n16528 & n16529);
  assign n16531 = (n13478 & n16291) | (n13478 & n16530) | (n16291 & n16530);
  assign n16532 = (n13478 & n16292) | (n13478 & n16530) | (n16292 & n16530);
  assign n16533 = (n16148 & n16531) | (n16148 & n16532) | (n16531 & n16532);
  assign n7833 = ~n16527 & n16533;
  assign n7834 = x77 & x83;
  assign n7835 = n7833 & n7834;
  assign n7836 = n7833 | n7834;
  assign n7837 = ~n7835 & n7836;
  assign n7838 = n16508 & n7837;
  assign n7839 = n16508 | n7837;
  assign n7840 = ~n7838 & n7839;
  assign n7841 = x76 & x84;
  assign n7842 = n7840 & n7841;
  assign n7843 = n7840 | n7841;
  assign n7844 = ~n7842 & n7843;
  assign n13480 = n7601 & n7844;
  assign n16534 = (n7844 & n13376) | (n7844 & n13480) | (n13376 & n13480);
  assign n16535 = (n7844 & n13377) | (n7844 & n13480) | (n13377 & n13480);
  assign n16536 = (n13173 & n16534) | (n13173 & n16535) | (n16534 & n16535);
  assign n13482 = n7601 | n7844;
  assign n16537 = n13376 | n13482;
  assign n16538 = n13377 | n13482;
  assign n16539 = (n13173 & n16537) | (n13173 & n16538) | (n16537 & n16538);
  assign n7847 = ~n16536 & n16539;
  assign n7848 = x75 & x85;
  assign n7849 = n7847 & n7848;
  assign n7850 = n7847 | n7848;
  assign n7851 = ~n7849 & n7850;
  assign n49952 = n7608 & n7851;
  assign n49953 = (n7851 & n13382) | (n7851 & n49952) | (n13382 & n49952);
  assign n16501 = n7371 | n7608;
  assign n16502 = (n7608 & n7610) | (n7608 & n16501) | (n7610 & n16501);
  assign n16541 = n7851 & n16502;
  assign n16542 = (n13261 & n49953) | (n13261 & n16541) | (n49953 & n16541);
  assign n49954 = n7608 | n7851;
  assign n49955 = n13382 | n49954;
  assign n16544 = n7851 | n16502;
  assign n16545 = (n13261 & n49955) | (n13261 & n16544) | (n49955 & n16544);
  assign n7854 = ~n16542 & n16545;
  assign n7855 = x74 & x86;
  assign n7856 = n7854 & n7855;
  assign n7857 = n7854 | n7855;
  assign n7858 = ~n7856 & n7857;
  assign n13454 = n7615 | n7617;
  assign n13484 = n7858 & n13454;
  assign n13485 = n7615 & n7858;
  assign n16546 = (n13343 & n13484) | (n13343 & n13485) | (n13484 & n13485);
  assign n16547 = (n13484 & n13485) | (n13484 & n16425) | (n13485 & n16425);
  assign n16548 = (n13203 & n16546) | (n13203 & n16547) | (n16546 & n16547);
  assign n13487 = n7858 | n13454;
  assign n13488 = n7615 | n7858;
  assign n16549 = (n13343 & n13487) | (n13343 & n13488) | (n13487 & n13488);
  assign n16550 = (n13487 & n13488) | (n13487 & n16425) | (n13488 & n16425);
  assign n16551 = (n13203 & n16549) | (n13203 & n16550) | (n16549 & n16550);
  assign n7861 = ~n16548 & n16551;
  assign n7862 = x73 & x87;
  assign n7863 = n7861 & n7862;
  assign n7864 = n7861 | n7862;
  assign n7865 = ~n7863 & n7864;
  assign n13490 = n7622 & n7865;
  assign n13491 = (n7865 & n13390) | (n7865 & n13490) | (n13390 & n13490);
  assign n13492 = n7622 | n7865;
  assign n13493 = n13390 | n13492;
  assign n7868 = ~n13491 & n13493;
  assign n7869 = x72 & x88;
  assign n7870 = n7868 & n7869;
  assign n7871 = n7868 | n7869;
  assign n7872 = ~n7870 & n7871;
  assign n7873 = n16500 & n7872;
  assign n7874 = n16500 | n7872;
  assign n7875 = ~n7873 & n7874;
  assign n7876 = x71 & x89;
  assign n7877 = n7875 & n7876;
  assign n7878 = n7875 | n7876;
  assign n7879 = ~n7877 & n7878;
  assign n13449 = n7636 | n7638;
  assign n13494 = n7879 & n13449;
  assign n13495 = n7636 & n7879;
  assign n13496 = (n16423 & n13494) | (n16423 & n13495) | (n13494 & n13495);
  assign n13497 = n7879 | n13449;
  assign n13498 = n7636 | n7879;
  assign n13499 = (n16423 & n13497) | (n16423 & n13498) | (n13497 & n13498);
  assign n7882 = ~n13496 & n13499;
  assign n7883 = x70 & x90;
  assign n7884 = n7882 & n7883;
  assign n7885 = n7882 | n7883;
  assign n7886 = ~n7884 & n7885;
  assign n13500 = n7643 & n7886;
  assign n13501 = (n7886 & n16474) | (n7886 & n13500) | (n16474 & n13500);
  assign n13502 = n7643 | n7886;
  assign n13503 = n16474 | n13502;
  assign n7889 = ~n13501 & n13503;
  assign n7890 = x69 & x91;
  assign n7891 = n7889 & n7890;
  assign n7892 = n7889 | n7890;
  assign n7893 = ~n7891 & n7892;
  assign n13447 = n7650 | n7652;
  assign n16552 = n7893 & n13447;
  assign n16494 = n7413 | n7650;
  assign n16495 = (n7650 & n7652) | (n7650 & n16494) | (n7652 & n16494);
  assign n16553 = n7893 & n16495;
  assign n16554 = (n16399 & n16552) | (n16399 & n16553) | (n16552 & n16553);
  assign n16555 = n7893 | n13447;
  assign n16556 = n7893 | n16495;
  assign n16557 = (n16399 & n16555) | (n16399 & n16556) | (n16555 & n16556);
  assign n7896 = ~n16554 & n16557;
  assign n7897 = x68 & x92;
  assign n7898 = n7896 & n7897;
  assign n7899 = n7896 | n7897;
  assign n7900 = ~n7898 & n7899;
  assign n13504 = n7657 & n7900;
  assign n16558 = (n7900 & n13408) | (n7900 & n13504) | (n13408 & n13504);
  assign n16559 = (n7659 & n7900) | (n7659 & n13504) | (n7900 & n13504);
  assign n16560 = (n13304 & n16558) | (n13304 & n16559) | (n16558 & n16559);
  assign n13506 = n7657 | n7900;
  assign n16561 = n13408 | n13506;
  assign n16562 = n7659 | n13506;
  assign n16563 = (n13304 & n16561) | (n13304 & n16562) | (n16561 & n16562);
  assign n7903 = ~n16560 & n16563;
  assign n7904 = x67 & x93;
  assign n7905 = n7903 & n7904;
  assign n7906 = n7903 | n7904;
  assign n7907 = ~n7905 & n7906;
  assign n13508 = n7664 & n7907;
  assign n13509 = (n7907 & n13413) | (n7907 & n13508) | (n13413 & n13508);
  assign n13510 = n7664 | n7907;
  assign n13511 = n13413 | n13510;
  assign n7910 = ~n13509 & n13511;
  assign n7911 = x66 & x94;
  assign n7912 = n7910 & n7911;
  assign n7913 = n7910 | n7911;
  assign n7914 = ~n7912 & n7913;
  assign n13512 = n7671 & n7914;
  assign n13513 = (n7914 & n13418) | (n7914 & n13512) | (n13418 & n13512);
  assign n13514 = n7671 | n7914;
  assign n13515 = n13418 | n13514;
  assign n7917 = ~n13513 & n13515;
  assign n7918 = x65 & x95;
  assign n7919 = n7917 & n7918;
  assign n7920 = n7917 | n7918;
  assign n7921 = ~n7919 & n7920;
  assign n13444 = n7678 | n7680;
  assign n13516 = n7921 & n13444;
  assign n13517 = n7678 & n7921;
  assign n13518 = (n13332 & n13516) | (n13332 & n13517) | (n13516 & n13517);
  assign n13519 = n7921 | n13444;
  assign n13520 = n7678 | n7921;
  assign n13521 = (n13332 & n13519) | (n13332 & n13520) | (n13519 & n13520);
  assign n7924 = ~n13518 & n13521;
  assign n7925 = x64 & x96;
  assign n7926 = n7924 & n7925;
  assign n7927 = n7924 | n7925;
  assign n7928 = ~n7926 & n7927;
  assign n13442 = n7685 | n7687;
  assign n16564 = n7928 & n13442;
  assign n16565 = n7685 & n7928;
  assign n16566 = (n13330 & n16564) | (n13330 & n16565) | (n16564 & n16565);
  assign n16567 = n7928 | n13442;
  assign n16568 = n7685 | n7928;
  assign n16569 = (n13330 & n16567) | (n13330 & n16568) | (n16567 & n16568);
  assign n7931 = ~n16566 & n16569;
  assign n7932 = x63 & x97;
  assign n7933 = n7931 & n7932;
  assign n7934 = n7931 | n7932;
  assign n7935 = ~n7933 & n7934;
  assign n13440 = n7692 | n7694;
  assign n16570 = n7935 & n13440;
  assign n16571 = n7692 & n7935;
  assign n16572 = (n13328 & n16570) | (n13328 & n16571) | (n16570 & n16571);
  assign n16573 = n7935 | n13440;
  assign n16574 = n7692 | n7935;
  assign n16575 = (n13328 & n16573) | (n13328 & n16574) | (n16573 & n16574);
  assign n7938 = ~n16572 & n16575;
  assign n7939 = x62 & x98;
  assign n7940 = n7938 & n7939;
  assign n7941 = n7938 | n7939;
  assign n7942 = ~n7940 & n7941;
  assign n7943 = n13439 & n7942;
  assign n7944 = n13439 | n7942;
  assign n7945 = ~n7943 & n7944;
  assign n7946 = x61 & x99;
  assign n7947 = n7945 & n7946;
  assign n7948 = n7945 | n7946;
  assign n7949 = ~n7947 & n7948;
  assign n7950 = n13437 & n7949;
  assign n7951 = n13437 | n7949;
  assign n7952 = ~n7950 & n7951;
  assign n7953 = x60 & x100;
  assign n7954 = n7952 & n7953;
  assign n7955 = n7952 | n7953;
  assign n7956 = ~n7954 & n7955;
  assign n7957 = n13435 & n7956;
  assign n7958 = n13435 | n7956;
  assign n7959 = ~n7957 & n7958;
  assign n7960 = x59 & x101;
  assign n7961 = n7959 & n7960;
  assign n7962 = n7959 | n7960;
  assign n7963 = ~n7961 & n7962;
  assign n7964 = n13433 & n7963;
  assign n7965 = n13433 | n7963;
  assign n7966 = ~n7964 & n7965;
  assign n7967 = x58 & x102;
  assign n7968 = n7966 & n7967;
  assign n7969 = n7966 | n7967;
  assign n7970 = ~n7968 & n7969;
  assign n7971 = n13431 & n7970;
  assign n7972 = n13431 | n7970;
  assign n7973 = ~n7971 & n7972;
  assign n7974 = x57 & x103;
  assign n7975 = n7973 & n7974;
  assign n7976 = n7973 | n7974;
  assign n7977 = ~n7975 & n7976;
  assign n7978 = n13429 & n7977;
  assign n7979 = n13429 | n7977;
  assign n7980 = ~n7978 & n7979;
  assign n7981 = x56 & x104;
  assign n7982 = n7980 & n7981;
  assign n7983 = n7980 | n7981;
  assign n7984 = ~n7982 & n7983;
  assign n7985 = n7799 & n7984;
  assign n7986 = n7799 | n7984;
  assign n7987 = ~n7985 & n7986;
  assign n7988 = x55 & x105;
  assign n7989 = n7987 & n7988;
  assign n7990 = n7987 | n7988;
  assign n7991 = ~n7989 & n7990;
  assign n7992 = n7798 & n7991;
  assign n7993 = n7798 | n7991;
  assign n7994 = ~n7992 & n7993;
  assign n7995 = x54 & x106;
  assign n7996 = n7994 & n7995;
  assign n7997 = n7994 | n7995;
  assign n7998 = ~n7996 & n7997;
  assign n7999 = n7797 & n7998;
  assign n8000 = n7797 | n7998;
  assign n8001 = ~n7999 & n8000;
  assign n8002 = x53 & x107;
  assign n8003 = n8001 & n8002;
  assign n8004 = n8001 | n8002;
  assign n8005 = ~n8003 & n8004;
  assign n8006 = n16493 & n8005;
  assign n8007 = n16493 | n8005;
  assign n8008 = ~n8006 & n8007;
  assign n8009 = x52 & x108;
  assign n8010 = n8008 & n8009;
  assign n8011 = n8008 | n8009;
  assign n8012 = ~n8010 & n8011;
  assign n8013 = n13427 & n8012;
  assign n8014 = n13427 | n8012;
  assign n8015 = ~n8013 & n8014;
  assign n8016 = x51 & x109;
  assign n8017 = n8015 & n8016;
  assign n8018 = n8015 | n8016;
  assign n8019 = ~n8017 & n8018;
  assign n8020 = n13425 & n8019;
  assign n8021 = n13425 | n8019;
  assign n8022 = ~n8020 & n8021;
  assign n8023 = x50 & x110;
  assign n8024 = n8022 & n8023;
  assign n8025 = n8022 | n8023;
  assign n8026 = ~n8024 & n8025;
  assign n8027 = n13423 & n8026;
  assign n8028 = n13423 | n8026;
  assign n8029 = ~n8027 & n8028;
  assign n8030 = x49 & x111;
  assign n8031 = n8029 & n8030;
  assign n8032 = n8029 | n8030;
  assign n8033 = ~n8031 & n8032;
  assign n8034 = n7790 & n8033;
  assign n8035 = n7790 | n8033;
  assign n8036 = ~n8034 & n8035;
  assign n49956 = n7789 | n8030;
  assign n49957 = (n7788 & n8030) | (n7788 & n49956) | (n8030 & n49956);
  assign n16577 = (n7790 & n8029) | (n7790 & n49957) | (n8029 & n49957);
  assign n13523 = (n8031 & n8033) | (n8031 & n16577) | (n8033 & n16577);
  assign n13524 = n8024 | n13423;
  assign n13525 = (n8024 & n8026) | (n8024 & n13524) | (n8026 & n13524);
  assign n13526 = n8017 | n13425;
  assign n13527 = (n8017 & n8019) | (n8017 & n13526) | (n8019 & n13526);
  assign n13528 = n8010 | n13427;
  assign n13529 = (n8010 & n8012) | (n8010 & n13528) | (n8012 & n13528);
  assign n16578 = n8003 | n16493;
  assign n16579 = (n8003 & n8005) | (n8003 & n16578) | (n8005 & n16578);
  assign n8042 = n7996 | n7999;
  assign n8043 = n7989 | n7992;
  assign n13530 = n7982 | n7984;
  assign n13531 = (n7799 & n7982) | (n7799 & n13530) | (n7982 & n13530);
  assign n13532 = n7975 | n7977;
  assign n13533 = (n7975 & n13429) | (n7975 & n13532) | (n13429 & n13532);
  assign n13534 = n7968 | n7970;
  assign n13535 = (n7968 & n13431) | (n7968 & n13534) | (n13431 & n13534);
  assign n13536 = n7961 | n7963;
  assign n13537 = (n7961 & n13433) | (n7961 & n13536) | (n13433 & n13536);
  assign n13538 = n7954 | n7956;
  assign n13539 = (n7954 & n13435) | (n7954 & n13538) | (n13435 & n13538);
  assign n13540 = n7947 | n7949;
  assign n13541 = (n7947 & n13437) | (n7947 & n13540) | (n13437 & n13540);
  assign n13441 = (n7692 & n13328) | (n7692 & n13440) | (n13328 & n13440);
  assign n13443 = (n7685 & n13330) | (n7685 & n13442) | (n13330 & n13442);
  assign n13448 = (n16399 & n16495) | (n16399 & n13447) | (n16495 & n13447);
  assign n13344 = (n13203 & n16425) | (n13203 & n13343) | (n16425 & n13343);
  assign n13456 = n7608 | n13382;
  assign n8067 = x79 & x82;
  assign n16586 = n7823 & n8067;
  assign n16587 = n16510 & n16586;
  assign n16588 = n16512 & n16586;
  assign n16589 = (n13267 & n16587) | (n13267 & n16588) | (n16587 & n16588);
  assign n16590 = (n16354 & n16587) | (n16354 & n16588) | (n16587 & n16588);
  assign n16591 = (n16089 & n16589) | (n16089 & n16590) | (n16589 & n16590);
  assign n16592 = n7823 | n8067;
  assign n16593 = (n8067 & n16510) | (n8067 & n16592) | (n16510 & n16592);
  assign n16594 = (n8067 & n16512) | (n8067 & n16592) | (n16512 & n16592);
  assign n16595 = (n13267 & n16593) | (n13267 & n16594) | (n16593 & n16594);
  assign n16596 = (n16354 & n16593) | (n16354 & n16594) | (n16593 & n16594);
  assign n16597 = (n16089 & n16595) | (n16089 & n16596) | (n16595 & n16596);
  assign n8070 = ~n16591 & n16597;
  assign n13574 = n7828 & n8070;
  assign n13575 = (n8070 & n16527) | (n8070 & n13574) | (n16527 & n13574);
  assign n13576 = n7828 | n8070;
  assign n13577 = n16527 | n13576;
  assign n8073 = ~n13575 & n13577;
  assign n8074 = x78 & x83;
  assign n8075 = n8073 & n8074;
  assign n8076 = n8073 | n8074;
  assign n8077 = ~n8075 & n8076;
  assign n13566 = n7835 | n7837;
  assign n13578 = n8077 & n13566;
  assign n13579 = n7835 & n8077;
  assign n13580 = (n16508 & n13578) | (n16508 & n13579) | (n13578 & n13579);
  assign n13581 = n8077 | n13566;
  assign n13582 = n7835 | n8077;
  assign n13583 = (n16508 & n13581) | (n16508 & n13582) | (n13581 & n13582);
  assign n8080 = ~n13580 & n13583;
  assign n8081 = x77 & x84;
  assign n8082 = n8080 & n8081;
  assign n8083 = n8080 | n8081;
  assign n8084 = ~n8082 & n8083;
  assign n16598 = n7601 | n7842;
  assign n16599 = (n7842 & n7844) | (n7842 & n16598) | (n7844 & n16598);
  assign n13584 = n8084 & n16599;
  assign n13564 = n7842 | n7844;
  assign n13585 = n8084 & n13564;
  assign n16600 = (n13376 & n13584) | (n13376 & n13585) | (n13584 & n13585);
  assign n16601 = (n13377 & n13584) | (n13377 & n13585) | (n13584 & n13585);
  assign n16602 = (n13173 & n16600) | (n13173 & n16601) | (n16600 & n16601);
  assign n13587 = n8084 | n16599;
  assign n13588 = n8084 | n13564;
  assign n16603 = (n13376 & n13587) | (n13376 & n13588) | (n13587 & n13588);
  assign n16604 = (n13377 & n13587) | (n13377 & n13588) | (n13587 & n13588);
  assign n16605 = (n13173 & n16603) | (n13173 & n16604) | (n16603 & n16604);
  assign n8087 = ~n16602 & n16605;
  assign n8088 = x76 & x85;
  assign n8089 = n8087 & n8088;
  assign n8090 = n8087 | n8088;
  assign n8091 = ~n8089 & n8090;
  assign n13561 = n7849 | n7851;
  assign n13590 = n8091 & n13561;
  assign n13591 = n7849 & n8091;
  assign n16606 = (n13456 & n13590) | (n13456 & n13591) | (n13590 & n13591);
  assign n16607 = (n13590 & n13591) | (n13590 & n16502) | (n13591 & n16502);
  assign n16608 = (n13261 & n16606) | (n13261 & n16607) | (n16606 & n16607);
  assign n13593 = n8091 | n13561;
  assign n13594 = n7849 | n8091;
  assign n16609 = (n13456 & n13593) | (n13456 & n13594) | (n13593 & n13594);
  assign n16610 = (n13593 & n13594) | (n13593 & n16502) | (n13594 & n16502);
  assign n16611 = (n13261 & n16609) | (n13261 & n16610) | (n16609 & n16610);
  assign n8094 = ~n16608 & n16611;
  assign n8095 = x75 & x86;
  assign n8096 = n8094 & n8095;
  assign n8097 = n8094 | n8095;
  assign n8098 = ~n8096 & n8097;
  assign n49958 = n7856 & n8098;
  assign n49959 = (n8098 & n13484) | (n8098 & n49958) | (n13484 & n49958);
  assign n16584 = n7615 | n7856;
  assign n16585 = (n7856 & n7858) | (n7856 & n16584) | (n7858 & n16584);
  assign n16613 = n8098 & n16585;
  assign n16614 = (n13344 & n49959) | (n13344 & n16613) | (n49959 & n16613);
  assign n49960 = n7856 | n8098;
  assign n49961 = n13484 | n49960;
  assign n16616 = n8098 | n16585;
  assign n16617 = (n13344 & n49961) | (n13344 & n16616) | (n49961 & n16616);
  assign n8101 = ~n16614 & n16617;
  assign n8102 = x74 & x87;
  assign n8103 = n8101 & n8102;
  assign n8104 = n8101 | n8102;
  assign n8105 = ~n8103 & n8104;
  assign n13556 = n7863 | n7865;
  assign n16618 = n8105 & n13556;
  assign n16582 = n7622 | n7863;
  assign n16583 = (n7863 & n7865) | (n7863 & n16582) | (n7865 & n16582);
  assign n16619 = n8105 & n16583;
  assign n16620 = (n13390 & n16618) | (n13390 & n16619) | (n16618 & n16619);
  assign n16621 = n8105 | n13556;
  assign n16622 = n8105 | n16583;
  assign n16623 = (n13390 & n16621) | (n13390 & n16622) | (n16621 & n16622);
  assign n8108 = ~n16620 & n16623;
  assign n8109 = x73 & x88;
  assign n8110 = n8108 & n8109;
  assign n8111 = n8108 | n8109;
  assign n8112 = ~n8110 & n8111;
  assign n13553 = n7870 | n7872;
  assign n13596 = n8112 & n13553;
  assign n13597 = n7870 & n8112;
  assign n13598 = (n16500 & n13596) | (n16500 & n13597) | (n13596 & n13597);
  assign n13599 = n8112 | n13553;
  assign n13600 = n7870 | n8112;
  assign n13601 = (n16500 & n13599) | (n16500 & n13600) | (n13599 & n13600);
  assign n8115 = ~n13598 & n13601;
  assign n8116 = x72 & x89;
  assign n8117 = n8115 & n8116;
  assign n8118 = n8115 | n8116;
  assign n8119 = ~n8117 & n8118;
  assign n13602 = n7877 & n8119;
  assign n16624 = (n8119 & n13495) | (n8119 & n13602) | (n13495 & n13602);
  assign n16625 = (n8119 & n13494) | (n8119 & n13602) | (n13494 & n13602);
  assign n16626 = (n16423 & n16624) | (n16423 & n16625) | (n16624 & n16625);
  assign n13604 = n7877 | n8119;
  assign n16627 = n13495 | n13604;
  assign n16628 = n13494 | n13604;
  assign n16629 = (n16423 & n16627) | (n16423 & n16628) | (n16627 & n16628);
  assign n8122 = ~n16626 & n16629;
  assign n8123 = x71 & x90;
  assign n8124 = n8122 & n8123;
  assign n8125 = n8122 | n8123;
  assign n8126 = ~n8124 & n8125;
  assign n13551 = n7884 | n7886;
  assign n16630 = n8126 & n13551;
  assign n16580 = n7643 | n7884;
  assign n16581 = (n7884 & n7886) | (n7884 & n16580) | (n7886 & n16580);
  assign n16631 = n8126 & n16581;
  assign n16632 = (n16474 & n16630) | (n16474 & n16631) | (n16630 & n16631);
  assign n16633 = n8126 | n13551;
  assign n16634 = n8126 | n16581;
  assign n16635 = (n16474 & n16633) | (n16474 & n16634) | (n16633 & n16634);
  assign n8129 = ~n16632 & n16635;
  assign n8130 = x70 & x91;
  assign n8131 = n8129 & n8130;
  assign n8132 = n8129 | n8130;
  assign n8133 = ~n8131 & n8132;
  assign n13548 = n7891 | n7893;
  assign n13606 = n8133 & n13548;
  assign n13607 = n7891 & n8133;
  assign n13608 = (n13448 & n13606) | (n13448 & n13607) | (n13606 & n13607);
  assign n13609 = n8133 | n13548;
  assign n13610 = n7891 | n8133;
  assign n13611 = (n13448 & n13609) | (n13448 & n13610) | (n13609 & n13610);
  assign n8136 = ~n13608 & n13611;
  assign n8137 = x69 & x92;
  assign n8138 = n8136 & n8137;
  assign n8139 = n8136 | n8137;
  assign n8140 = ~n8138 & n8139;
  assign n13612 = n7898 & n8140;
  assign n13613 = (n8140 & n16560) | (n8140 & n13612) | (n16560 & n13612);
  assign n13614 = n7898 | n8140;
  assign n13615 = n16560 | n13614;
  assign n8143 = ~n13613 & n13615;
  assign n8144 = x68 & x93;
  assign n8145 = n8143 & n8144;
  assign n8146 = n8143 | n8144;
  assign n8147 = ~n8145 & n8146;
  assign n13616 = n7905 & n8147;
  assign n13617 = (n8147 & n13509) | (n8147 & n13616) | (n13509 & n13616);
  assign n13618 = n7905 | n8147;
  assign n13619 = n13509 | n13618;
  assign n8150 = ~n13617 & n13619;
  assign n8151 = x67 & x94;
  assign n8152 = n8150 & n8151;
  assign n8153 = n8150 | n8151;
  assign n8154 = ~n8152 & n8153;
  assign n13620 = n7912 & n8154;
  assign n13621 = (n8154 & n13513) | (n8154 & n13620) | (n13513 & n13620);
  assign n13622 = n7912 | n8154;
  assign n13623 = n13513 | n13622;
  assign n8157 = ~n13621 & n13623;
  assign n8158 = x66 & x95;
  assign n8159 = n8157 & n8158;
  assign n8160 = n8157 | n8158;
  assign n8161 = ~n8159 & n8160;
  assign n13624 = n7919 & n8161;
  assign n13625 = (n8161 & n13518) | (n8161 & n13624) | (n13518 & n13624);
  assign n13626 = n7919 | n8161;
  assign n13627 = n13518 | n13626;
  assign n8164 = ~n13625 & n13627;
  assign n8165 = x65 & x96;
  assign n8166 = n8164 & n8165;
  assign n8167 = n8164 | n8165;
  assign n8168 = ~n8166 & n8167;
  assign n13546 = n7926 | n7928;
  assign n13628 = n8168 & n13546;
  assign n13629 = n7926 & n8168;
  assign n13630 = (n13443 & n13628) | (n13443 & n13629) | (n13628 & n13629);
  assign n13631 = n8168 | n13546;
  assign n13632 = n7926 | n8168;
  assign n13633 = (n13443 & n13631) | (n13443 & n13632) | (n13631 & n13632);
  assign n8171 = ~n13630 & n13633;
  assign n8172 = x64 & x97;
  assign n8173 = n8171 & n8172;
  assign n8174 = n8171 | n8172;
  assign n8175 = ~n8173 & n8174;
  assign n13544 = n7933 | n7935;
  assign n16636 = n8175 & n13544;
  assign n16637 = n7933 & n8175;
  assign n16638 = (n13441 & n16636) | (n13441 & n16637) | (n16636 & n16637);
  assign n16639 = n8175 | n13544;
  assign n16640 = n7933 | n8175;
  assign n16641 = (n13441 & n16639) | (n13441 & n16640) | (n16639 & n16640);
  assign n8178 = ~n16638 & n16641;
  assign n8179 = x63 & x98;
  assign n8180 = n8178 & n8179;
  assign n8181 = n8178 | n8179;
  assign n8182 = ~n8180 & n8181;
  assign n13542 = n7940 | n7942;
  assign n16642 = n8182 & n13542;
  assign n16643 = n7940 & n8182;
  assign n16644 = (n13439 & n16642) | (n13439 & n16643) | (n16642 & n16643);
  assign n16645 = n8182 | n13542;
  assign n16646 = n7940 | n8182;
  assign n16647 = (n13439 & n16645) | (n13439 & n16646) | (n16645 & n16646);
  assign n8185 = ~n16644 & n16647;
  assign n8186 = x62 & x99;
  assign n8187 = n8185 & n8186;
  assign n8188 = n8185 | n8186;
  assign n8189 = ~n8187 & n8188;
  assign n8190 = n13541 & n8189;
  assign n8191 = n13541 | n8189;
  assign n8192 = ~n8190 & n8191;
  assign n8193 = x61 & x100;
  assign n8194 = n8192 & n8193;
  assign n8195 = n8192 | n8193;
  assign n8196 = ~n8194 & n8195;
  assign n8197 = n13539 & n8196;
  assign n8198 = n13539 | n8196;
  assign n8199 = ~n8197 & n8198;
  assign n8200 = x60 & x101;
  assign n8201 = n8199 & n8200;
  assign n8202 = n8199 | n8200;
  assign n8203 = ~n8201 & n8202;
  assign n8204 = n13537 & n8203;
  assign n8205 = n13537 | n8203;
  assign n8206 = ~n8204 & n8205;
  assign n8207 = x59 & x102;
  assign n8208 = n8206 & n8207;
  assign n8209 = n8206 | n8207;
  assign n8210 = ~n8208 & n8209;
  assign n8211 = n13535 & n8210;
  assign n8212 = n13535 | n8210;
  assign n8213 = ~n8211 & n8212;
  assign n8214 = x58 & x103;
  assign n8215 = n8213 & n8214;
  assign n8216 = n8213 | n8214;
  assign n8217 = ~n8215 & n8216;
  assign n8218 = n13533 & n8217;
  assign n8219 = n13533 | n8217;
  assign n8220 = ~n8218 & n8219;
  assign n8221 = x57 & x104;
  assign n8222 = n8220 & n8221;
  assign n8223 = n8220 | n8221;
  assign n8224 = ~n8222 & n8223;
  assign n8225 = n13531 & n8224;
  assign n8226 = n13531 | n8224;
  assign n8227 = ~n8225 & n8226;
  assign n8228 = x56 & x105;
  assign n8229 = n8227 & n8228;
  assign n8230 = n8227 | n8228;
  assign n8231 = ~n8229 & n8230;
  assign n8232 = n8043 & n8231;
  assign n8233 = n8043 | n8231;
  assign n8234 = ~n8232 & n8233;
  assign n8235 = x55 & x106;
  assign n8236 = n8234 & n8235;
  assign n8237 = n8234 | n8235;
  assign n8238 = ~n8236 & n8237;
  assign n8239 = n8042 & n8238;
  assign n8240 = n8042 | n8238;
  assign n8241 = ~n8239 & n8240;
  assign n8242 = x54 & x107;
  assign n8243 = n8241 & n8242;
  assign n8244 = n8241 | n8242;
  assign n8245 = ~n8243 & n8244;
  assign n8246 = n16579 & n8245;
  assign n8247 = n16579 | n8245;
  assign n8248 = ~n8246 & n8247;
  assign n8249 = x53 & x108;
  assign n8250 = n8248 & n8249;
  assign n8251 = n8248 | n8249;
  assign n8252 = ~n8250 & n8251;
  assign n8253 = n13529 & n8252;
  assign n8254 = n13529 | n8252;
  assign n8255 = ~n8253 & n8254;
  assign n8256 = x52 & x109;
  assign n8257 = n8255 & n8256;
  assign n8258 = n8255 | n8256;
  assign n8259 = ~n8257 & n8258;
  assign n8260 = n13527 & n8259;
  assign n8261 = n13527 | n8259;
  assign n8262 = ~n8260 & n8261;
  assign n8263 = x51 & x110;
  assign n8264 = n8262 & n8263;
  assign n8265 = n8262 | n8263;
  assign n8266 = ~n8264 & n8265;
  assign n8267 = n13525 & n8266;
  assign n8268 = n13525 | n8266;
  assign n8269 = ~n8267 & n8268;
  assign n8270 = x50 & x111;
  assign n8271 = n8269 & n8270;
  assign n8272 = n8269 | n8270;
  assign n8273 = ~n8271 & n8272;
  assign n8274 = n13523 & n8273;
  assign n8275 = n13523 | n8273;
  assign n8276 = ~n8274 & n8275;
  assign n13634 = n8271 | n13523;
  assign n13635 = (n8271 & n8273) | (n8271 & n13634) | (n8273 & n13634);
  assign n13636 = n8264 | n13525;
  assign n13637 = (n8264 & n8266) | (n8264 & n13636) | (n8266 & n13636);
  assign n13638 = n8257 | n13527;
  assign n13639 = (n8257 & n8259) | (n8257 & n13638) | (n8259 & n13638);
  assign n13640 = n8250 | n13529;
  assign n13641 = (n8250 & n8252) | (n8250 & n13640) | (n8252 & n13640);
  assign n16648 = n8243 | n16579;
  assign n16649 = (n8243 & n8245) | (n8243 & n16648) | (n8245 & n16648);
  assign n8282 = n8236 | n8239;
  assign n13642 = n8229 | n8231;
  assign n13643 = (n8043 & n8229) | (n8043 & n13642) | (n8229 & n13642);
  assign n13644 = n8222 | n8224;
  assign n13645 = (n8222 & n13531) | (n8222 & n13644) | (n13531 & n13644);
  assign n13646 = n8215 | n8217;
  assign n13647 = (n8215 & n13533) | (n8215 & n13646) | (n13533 & n13646);
  assign n13648 = n8208 | n8210;
  assign n13649 = (n8208 & n13535) | (n8208 & n13648) | (n13535 & n13648);
  assign n13650 = n8201 | n8203;
  assign n13651 = (n8201 & n13537) | (n8201 & n13650) | (n13537 & n13650);
  assign n13652 = n8194 | n8196;
  assign n13653 = (n8194 & n13539) | (n8194 & n13652) | (n13539 & n13652);
  assign n13543 = (n7940 & n13439) | (n7940 & n13542) | (n13439 & n13542);
  assign n13545 = (n7933 & n13441) | (n7933 & n13544) | (n13441 & n13544);
  assign n13666 = n8117 | n8119;
  assign n16652 = n7877 | n8117;
  assign n16653 = (n8117 & n8119) | (n8117 & n16652) | (n8119 & n16652);
  assign n16654 = (n13495 & n13666) | (n13495 & n16653) | (n13666 & n16653);
  assign n16655 = (n13494 & n13666) | (n13494 & n16653) | (n13666 & n16653);
  assign n16656 = (n16423 & n16654) | (n16423 & n16655) | (n16654 & n16655);
  assign n13557 = (n13390 & n16583) | (n13390 & n13556) | (n16583 & n13556);
  assign n13559 = n7856 | n13484;
  assign n16657 = n8089 | n8091;
  assign n16658 = (n8089 & n13561) | (n8089 & n16657) | (n13561 & n16657);
  assign n16659 = n7849 | n8089;
  assign n16660 = (n8089 & n8091) | (n8089 & n16659) | (n8091 & n16659);
  assign n16661 = (n13456 & n16658) | (n13456 & n16660) | (n16658 & n16660);
  assign n16662 = (n16502 & n16658) | (n16502 & n16660) | (n16658 & n16660);
  assign n16663 = (n13261 & n16661) | (n13261 & n16662) | (n16661 & n16662);
  assign n8307 = x79 & x83;
  assign n16664 = n8070 | n16591;
  assign n16665 = (n7828 & n16591) | (n7828 & n16664) | (n16591 & n16664);
  assign n13681 = n8307 & n16665;
  assign n66363 = n8307 & n16587;
  assign n66364 = n8307 & n16588;
  assign n66365 = (n16354 & n66363) | (n16354 & n66364) | (n66363 & n66364);
  assign n66366 = (n13267 & n66363) | (n13267 & n66364) | (n66363 & n66364);
  assign n49964 = (n16089 & n66365) | (n16089 & n66366) | (n66365 & n66366);
  assign n16667 = (n8070 & n8307) | (n8070 & n49964) | (n8307 & n49964);
  assign n13683 = (n16527 & n13681) | (n16527 & n16667) | (n13681 & n16667);
  assign n13684 = n8307 | n16665;
  assign n66367 = n8307 | n16587;
  assign n66368 = n8307 | n16588;
  assign n66369 = (n16354 & n66367) | (n16354 & n66368) | (n66367 & n66368);
  assign n66370 = (n13267 & n66367) | (n13267 & n66368) | (n66367 & n66368);
  assign n49967 = (n16089 & n66369) | (n16089 & n66370) | (n66369 & n66370);
  assign n16669 = n8070 | n49967;
  assign n13686 = (n16527 & n13684) | (n16527 & n16669) | (n13684 & n16669);
  assign n8310 = ~n13683 & n13686;
  assign n16670 = n8075 & n8310;
  assign n16671 = (n8310 & n13578) | (n8310 & n16670) | (n13578 & n16670);
  assign n16672 = n7835 | n8075;
  assign n16673 = (n8075 & n8077) | (n8075 & n16672) | (n8077 & n16672);
  assign n13688 = n8310 & n16673;
  assign n13689 = (n16508 & n16671) | (n16508 & n13688) | (n16671 & n13688);
  assign n16674 = n8075 | n8310;
  assign n16675 = n13578 | n16674;
  assign n13691 = n8310 | n16673;
  assign n13692 = (n16508 & n16675) | (n16508 & n13691) | (n16675 & n13691);
  assign n8313 = ~n13689 & n13692;
  assign n8314 = x78 & x84;
  assign n8315 = n8313 & n8314;
  assign n8316 = n8313 | n8314;
  assign n8317 = ~n8315 & n8316;
  assign n13693 = n8082 & n8317;
  assign n13694 = (n8317 & n16602) | (n8317 & n13693) | (n16602 & n13693);
  assign n13695 = n8082 | n8317;
  assign n13696 = n16602 | n13695;
  assign n8320 = ~n13694 & n13696;
  assign n8321 = x77 & x85;
  assign n8322 = n8320 & n8321;
  assign n8323 = n8320 | n8321;
  assign n8324 = ~n8322 & n8323;
  assign n8325 = n16663 & n8324;
  assign n8326 = n16663 | n8324;
  assign n8327 = ~n8325 & n8326;
  assign n8328 = x76 & x86;
  assign n8329 = n8327 & n8328;
  assign n8330 = n8327 | n8328;
  assign n8331 = ~n8329 & n8330;
  assign n13670 = n8096 | n8098;
  assign n13697 = n8331 & n13670;
  assign n13698 = n8096 & n8331;
  assign n16676 = (n13559 & n13697) | (n13559 & n13698) | (n13697 & n13698);
  assign n16677 = (n13697 & n13698) | (n13697 & n16585) | (n13698 & n16585);
  assign n16678 = (n13344 & n16676) | (n13344 & n16677) | (n16676 & n16677);
  assign n13700 = n8331 | n13670;
  assign n13701 = n8096 | n8331;
  assign n16679 = (n13559 & n13700) | (n13559 & n13701) | (n13700 & n13701);
  assign n16680 = (n13700 & n13701) | (n13700 & n16585) | (n13701 & n16585);
  assign n16681 = (n13344 & n16679) | (n13344 & n16680) | (n16679 & n16680);
  assign n8334 = ~n16678 & n16681;
  assign n8335 = x75 & x87;
  assign n8336 = n8334 & n8335;
  assign n8337 = n8334 | n8335;
  assign n8338 = ~n8336 & n8337;
  assign n13668 = n8103 | n8105;
  assign n13703 = n8338 & n13668;
  assign n13704 = n8103 & n8338;
  assign n13705 = (n13557 & n13703) | (n13557 & n13704) | (n13703 & n13704);
  assign n13706 = n8338 | n13668;
  assign n13707 = n8103 | n8338;
  assign n13708 = (n13557 & n13706) | (n13557 & n13707) | (n13706 & n13707);
  assign n8341 = ~n13705 & n13708;
  assign n8342 = x74 & x88;
  assign n8343 = n8341 & n8342;
  assign n8344 = n8341 | n8342;
  assign n8345 = ~n8343 & n8344;
  assign n13709 = n8110 & n8345;
  assign n13710 = (n8345 & n13598) | (n8345 & n13709) | (n13598 & n13709);
  assign n13711 = n8110 | n8345;
  assign n13712 = n13598 | n13711;
  assign n8348 = ~n13710 & n13712;
  assign n8349 = x73 & x89;
  assign n8350 = n8348 & n8349;
  assign n8351 = n8348 | n8349;
  assign n8352 = ~n8350 & n8351;
  assign n8353 = n16656 & n8352;
  assign n8354 = n16656 | n8352;
  assign n8355 = ~n8353 & n8354;
  assign n8356 = x72 & x90;
  assign n8357 = n8355 & n8356;
  assign n8358 = n8355 | n8356;
  assign n8359 = ~n8357 & n8358;
  assign n13663 = n8124 | n8126;
  assign n13713 = n8359 & n13663;
  assign n13714 = n8124 & n8359;
  assign n16682 = (n13551 & n13713) | (n13551 & n13714) | (n13713 & n13714);
  assign n16683 = (n13713 & n13714) | (n13713 & n16581) | (n13714 & n16581);
  assign n16684 = (n16474 & n16682) | (n16474 & n16683) | (n16682 & n16683);
  assign n13716 = n8359 | n13663;
  assign n13717 = n8124 | n8359;
  assign n16685 = (n13551 & n13716) | (n13551 & n13717) | (n13716 & n13717);
  assign n16686 = (n13716 & n13717) | (n13716 & n16581) | (n13717 & n16581);
  assign n16687 = (n16474 & n16685) | (n16474 & n16686) | (n16685 & n16686);
  assign n8362 = ~n16684 & n16687;
  assign n8363 = x71 & x91;
  assign n8364 = n8362 & n8363;
  assign n8365 = n8362 | n8363;
  assign n8366 = ~n8364 & n8365;
  assign n13719 = n8131 & n8366;
  assign n16688 = (n8366 & n13606) | (n8366 & n13719) | (n13606 & n13719);
  assign n16689 = (n8366 & n13607) | (n8366 & n13719) | (n13607 & n13719);
  assign n16690 = (n13448 & n16688) | (n13448 & n16689) | (n16688 & n16689);
  assign n13721 = n8131 | n8366;
  assign n16691 = n13606 | n13721;
  assign n16692 = n13607 | n13721;
  assign n16693 = (n13448 & n16691) | (n13448 & n16692) | (n16691 & n16692);
  assign n8369 = ~n16690 & n16693;
  assign n8370 = x70 & x92;
  assign n8371 = n8369 & n8370;
  assign n8372 = n8369 | n8370;
  assign n8373 = ~n8371 & n8372;
  assign n13661 = n8138 | n8140;
  assign n16694 = n8373 & n13661;
  assign n16650 = n7898 | n8138;
  assign n16651 = (n8138 & n8140) | (n8138 & n16650) | (n8140 & n16650);
  assign n16695 = n8373 & n16651;
  assign n16696 = (n16560 & n16694) | (n16560 & n16695) | (n16694 & n16695);
  assign n16697 = n8373 | n13661;
  assign n16698 = n8373 | n16651;
  assign n16699 = (n16560 & n16697) | (n16560 & n16698) | (n16697 & n16698);
  assign n8376 = ~n16696 & n16699;
  assign n8377 = x69 & x93;
  assign n8378 = n8376 & n8377;
  assign n8379 = n8376 | n8377;
  assign n8380 = ~n8378 & n8379;
  assign n13723 = n8145 & n8380;
  assign n16700 = (n8380 & n13616) | (n8380 & n13723) | (n13616 & n13723);
  assign n16701 = (n8147 & n8380) | (n8147 & n13723) | (n8380 & n13723);
  assign n16702 = (n13509 & n16700) | (n13509 & n16701) | (n16700 & n16701);
  assign n13725 = n8145 | n8380;
  assign n16703 = n13616 | n13725;
  assign n16704 = n8147 | n13725;
  assign n16705 = (n13509 & n16703) | (n13509 & n16704) | (n16703 & n16704);
  assign n8383 = ~n16702 & n16705;
  assign n8384 = x68 & x94;
  assign n8385 = n8383 & n8384;
  assign n8386 = n8383 | n8384;
  assign n8387 = ~n8385 & n8386;
  assign n13727 = n8152 & n8387;
  assign n13728 = (n8387 & n13621) | (n8387 & n13727) | (n13621 & n13727);
  assign n13729 = n8152 | n8387;
  assign n13730 = n13621 | n13729;
  assign n8390 = ~n13728 & n13730;
  assign n8391 = x67 & x95;
  assign n8392 = n8390 & n8391;
  assign n8393 = n8390 | n8391;
  assign n8394 = ~n8392 & n8393;
  assign n13731 = n8159 & n8394;
  assign n13732 = (n8394 & n13625) | (n8394 & n13731) | (n13625 & n13731);
  assign n13733 = n8159 | n8394;
  assign n13734 = n13625 | n13733;
  assign n8397 = ~n13732 & n13734;
  assign n8398 = x66 & x96;
  assign n8399 = n8397 & n8398;
  assign n8400 = n8397 | n8398;
  assign n8401 = ~n8399 & n8400;
  assign n13735 = n8166 & n8401;
  assign n13736 = (n8401 & n13630) | (n8401 & n13735) | (n13630 & n13735);
  assign n13737 = n8166 | n8401;
  assign n13738 = n13630 | n13737;
  assign n8404 = ~n13736 & n13738;
  assign n8405 = x65 & x97;
  assign n8406 = n8404 & n8405;
  assign n8407 = n8404 | n8405;
  assign n8408 = ~n8406 & n8407;
  assign n13658 = n8173 | n8175;
  assign n13739 = n8408 & n13658;
  assign n13740 = n8173 & n8408;
  assign n13741 = (n13545 & n13739) | (n13545 & n13740) | (n13739 & n13740);
  assign n13742 = n8408 | n13658;
  assign n13743 = n8173 | n8408;
  assign n13744 = (n13545 & n13742) | (n13545 & n13743) | (n13742 & n13743);
  assign n8411 = ~n13741 & n13744;
  assign n8412 = x64 & x98;
  assign n8413 = n8411 & n8412;
  assign n8414 = n8411 | n8412;
  assign n8415 = ~n8413 & n8414;
  assign n13656 = n8180 | n8182;
  assign n16706 = n8415 & n13656;
  assign n16707 = n8180 & n8415;
  assign n16708 = (n13543 & n16706) | (n13543 & n16707) | (n16706 & n16707);
  assign n16709 = n8415 | n13656;
  assign n16710 = n8180 | n8415;
  assign n16711 = (n13543 & n16709) | (n13543 & n16710) | (n16709 & n16710);
  assign n8418 = ~n16708 & n16711;
  assign n8419 = x63 & x99;
  assign n8420 = n8418 & n8419;
  assign n8421 = n8418 | n8419;
  assign n8422 = ~n8420 & n8421;
  assign n13654 = n8187 | n8189;
  assign n16712 = n8422 & n13654;
  assign n16713 = n8187 & n8422;
  assign n16714 = (n13541 & n16712) | (n13541 & n16713) | (n16712 & n16713);
  assign n16715 = n8422 | n13654;
  assign n16716 = n8187 | n8422;
  assign n16717 = (n13541 & n16715) | (n13541 & n16716) | (n16715 & n16716);
  assign n8425 = ~n16714 & n16717;
  assign n8426 = x62 & x100;
  assign n8427 = n8425 & n8426;
  assign n8428 = n8425 | n8426;
  assign n8429 = ~n8427 & n8428;
  assign n8430 = n13653 & n8429;
  assign n8431 = n13653 | n8429;
  assign n8432 = ~n8430 & n8431;
  assign n8433 = x61 & x101;
  assign n8434 = n8432 & n8433;
  assign n8435 = n8432 | n8433;
  assign n8436 = ~n8434 & n8435;
  assign n8437 = n13651 & n8436;
  assign n8438 = n13651 | n8436;
  assign n8439 = ~n8437 & n8438;
  assign n8440 = x60 & x102;
  assign n8441 = n8439 & n8440;
  assign n8442 = n8439 | n8440;
  assign n8443 = ~n8441 & n8442;
  assign n8444 = n13649 & n8443;
  assign n8445 = n13649 | n8443;
  assign n8446 = ~n8444 & n8445;
  assign n8447 = x59 & x103;
  assign n8448 = n8446 & n8447;
  assign n8449 = n8446 | n8447;
  assign n8450 = ~n8448 & n8449;
  assign n8451 = n13647 & n8450;
  assign n8452 = n13647 | n8450;
  assign n8453 = ~n8451 & n8452;
  assign n8454 = x58 & x104;
  assign n8455 = n8453 & n8454;
  assign n8456 = n8453 | n8454;
  assign n8457 = ~n8455 & n8456;
  assign n8458 = n13645 & n8457;
  assign n8459 = n13645 | n8457;
  assign n8460 = ~n8458 & n8459;
  assign n8461 = x57 & x105;
  assign n8462 = n8460 & n8461;
  assign n8463 = n8460 | n8461;
  assign n8464 = ~n8462 & n8463;
  assign n8465 = n13643 & n8464;
  assign n8466 = n13643 | n8464;
  assign n8467 = ~n8465 & n8466;
  assign n8468 = x56 & x106;
  assign n8469 = n8467 & n8468;
  assign n8470 = n8467 | n8468;
  assign n8471 = ~n8469 & n8470;
  assign n8472 = n8282 & n8471;
  assign n8473 = n8282 | n8471;
  assign n8474 = ~n8472 & n8473;
  assign n8475 = x55 & x107;
  assign n8476 = n8474 & n8475;
  assign n8477 = n8474 | n8475;
  assign n8478 = ~n8476 & n8477;
  assign n8479 = n16649 & n8478;
  assign n8480 = n16649 | n8478;
  assign n8481 = ~n8479 & n8480;
  assign n8482 = x54 & x108;
  assign n8483 = n8481 & n8482;
  assign n8484 = n8481 | n8482;
  assign n8485 = ~n8483 & n8484;
  assign n8486 = n13641 & n8485;
  assign n8487 = n13641 | n8485;
  assign n8488 = ~n8486 & n8487;
  assign n8489 = x53 & x109;
  assign n8490 = n8488 & n8489;
  assign n8491 = n8488 | n8489;
  assign n8492 = ~n8490 & n8491;
  assign n8493 = n13639 & n8492;
  assign n8494 = n13639 | n8492;
  assign n8495 = ~n8493 & n8494;
  assign n8496 = x52 & x110;
  assign n8497 = n8495 & n8496;
  assign n8498 = n8495 | n8496;
  assign n8499 = ~n8497 & n8498;
  assign n8500 = n13637 & n8499;
  assign n8501 = n13637 | n8499;
  assign n8502 = ~n8500 & n8501;
  assign n8503 = x51 & x111;
  assign n8504 = n8502 & n8503;
  assign n8505 = n8502 | n8503;
  assign n8506 = ~n8504 & n8505;
  assign n8507 = n13635 & n8506;
  assign n8508 = n13635 | n8506;
  assign n8509 = ~n8507 & n8508;
  assign n13745 = n8504 | n13635;
  assign n13746 = (n8504 & n8506) | (n8504 & n13745) | (n8506 & n13745);
  assign n13747 = n8497 | n13637;
  assign n13748 = (n8497 & n8499) | (n8497 & n13747) | (n8499 & n13747);
  assign n13749 = n8490 | n13639;
  assign n13750 = (n8490 & n8492) | (n8490 & n13749) | (n8492 & n13749);
  assign n13751 = n8483 | n13641;
  assign n13752 = (n8483 & n8485) | (n8483 & n13751) | (n8485 & n13751);
  assign n16718 = n8476 | n16649;
  assign n16719 = (n8476 & n8478) | (n8476 & n16718) | (n8478 & n16718);
  assign n13753 = n8469 | n8471;
  assign n13754 = (n8282 & n8469) | (n8282 & n13753) | (n8469 & n13753);
  assign n13755 = n8462 | n8464;
  assign n13756 = (n8462 & n13643) | (n8462 & n13755) | (n13643 & n13755);
  assign n13757 = n8455 | n8457;
  assign n13758 = (n8455 & n13645) | (n8455 & n13757) | (n13645 & n13757);
  assign n13759 = n8448 | n8450;
  assign n13760 = (n8448 & n13647) | (n8448 & n13759) | (n13647 & n13759);
  assign n13761 = n8441 | n8443;
  assign n13762 = (n8441 & n13649) | (n8441 & n13761) | (n13649 & n13761);
  assign n13763 = n8434 | n8436;
  assign n13764 = (n8434 & n13651) | (n8434 & n13763) | (n13651 & n13763);
  assign n13655 = (n8187 & n13541) | (n8187 & n13654) | (n13541 & n13654);
  assign n13657 = (n8180 & n13543) | (n8180 & n13656) | (n13543 & n13656);
  assign n13662 = (n16560 & n16651) | (n16560 & n13661) | (n16651 & n13661);
  assign n13774 = n8364 | n8366;
  assign n16720 = n8131 | n8364;
  assign n16721 = (n8364 & n8366) | (n8364 & n16720) | (n8366 & n16720);
  assign n16722 = (n13606 & n13774) | (n13606 & n16721) | (n13774 & n16721);
  assign n16723 = (n13607 & n13774) | (n13607 & n16721) | (n13774 & n16721);
  assign n16724 = (n13448 & n16722) | (n13448 & n16723) | (n16722 & n16723);
  assign n13560 = (n13344 & n16585) | (n13344 & n13559) | (n16585 & n13559);
  assign n8539 = x79 & x84;
  assign n16729 = n8310 | n13683;
  assign n49968 = (n8075 & n13683) | (n8075 & n16729) | (n13683 & n16729);
  assign n49969 = n8539 & n49968;
  assign n66372 = n8539 & n13681;
  assign n66373 = n8539 & n16667;
  assign n66374 = (n16527 & n66372) | (n16527 & n66373) | (n66372 & n66373);
  assign n66371 = (n8310 & n8539) | (n8310 & n66374) | (n8539 & n66374);
  assign n49971 = (n13578 & n49969) | (n13578 & n66371) | (n49969 & n66371);
  assign n49973 = (n16673 & n66371) | (n16673 & n66374) | (n66371 & n66374);
  assign n16735 = (n16508 & n49971) | (n16508 & n49973) | (n49971 & n49973);
  assign n49974 = n8539 | n49968;
  assign n66376 = n8539 | n13681;
  assign n66377 = n8539 | n16667;
  assign n66378 = (n16527 & n66376) | (n16527 & n66377) | (n66376 & n66377);
  assign n66375 = n8310 | n66378;
  assign n49976 = (n13578 & n49974) | (n13578 & n66375) | (n49974 & n66375);
  assign n49978 = (n16673 & n66375) | (n16673 & n66378) | (n66375 & n66378);
  assign n16738 = (n16508 & n49976) | (n16508 & n49978) | (n49976 & n49978);
  assign n8542 = ~n16735 & n16738;
  assign n16739 = n8082 | n8315;
  assign n16740 = (n8315 & n8317) | (n8315 & n16739) | (n8317 & n16739);
  assign n13792 = n8542 & n16740;
  assign n16741 = n8315 & n8542;
  assign n16742 = (n8317 & n8542) | (n8317 & n16741) | (n8542 & n16741);
  assign n13794 = (n16602 & n13792) | (n16602 & n16742) | (n13792 & n16742);
  assign n13795 = n8542 | n16740;
  assign n16743 = n8315 | n8542;
  assign n16744 = n8317 | n16743;
  assign n13797 = (n16602 & n13795) | (n16602 & n16744) | (n13795 & n16744);
  assign n8545 = ~n13794 & n13797;
  assign n8546 = x78 & x85;
  assign n8547 = n8545 & n8546;
  assign n8548 = n8545 | n8546;
  assign n8549 = ~n8547 & n8548;
  assign n13784 = n8322 | n8324;
  assign n13798 = n8549 & n13784;
  assign n13799 = n8322 & n8549;
  assign n13800 = (n16663 & n13798) | (n16663 & n13799) | (n13798 & n13799);
  assign n13801 = n8549 | n13784;
  assign n13802 = n8322 | n8549;
  assign n13803 = (n16663 & n13801) | (n16663 & n13802) | (n13801 & n13802);
  assign n8552 = ~n13800 & n13803;
  assign n8553 = x77 & x86;
  assign n8554 = n8552 & n8553;
  assign n8555 = n8552 | n8553;
  assign n8556 = ~n8554 & n8555;
  assign n49979 = n8329 & n8556;
  assign n49980 = (n8556 & n13697) | (n8556 & n49979) | (n13697 & n49979);
  assign n16727 = n8096 | n8329;
  assign n16728 = (n8329 & n8331) | (n8329 & n16727) | (n8331 & n16727);
  assign n16746 = n8556 & n16728;
  assign n16747 = (n13560 & n49980) | (n13560 & n16746) | (n49980 & n16746);
  assign n49981 = n8329 | n8556;
  assign n49982 = n13697 | n49981;
  assign n16749 = n8556 | n16728;
  assign n16750 = (n13560 & n49982) | (n13560 & n16749) | (n49982 & n16749);
  assign n8559 = ~n16747 & n16750;
  assign n8560 = x76 & x87;
  assign n8561 = n8559 & n8560;
  assign n8562 = n8559 | n8560;
  assign n8563 = ~n8561 & n8562;
  assign n13804 = n8336 & n8563;
  assign n16751 = (n8563 & n13703) | (n8563 & n13804) | (n13703 & n13804);
  assign n16752 = (n8563 & n13704) | (n8563 & n13804) | (n13704 & n13804);
  assign n16753 = (n13557 & n16751) | (n13557 & n16752) | (n16751 & n16752);
  assign n13806 = n8336 | n8563;
  assign n16754 = n13703 | n13806;
  assign n16755 = n13704 | n13806;
  assign n16756 = (n13557 & n16754) | (n13557 & n16755) | (n16754 & n16755);
  assign n8566 = ~n16753 & n16756;
  assign n8567 = x75 & x88;
  assign n8568 = n8566 & n8567;
  assign n8569 = n8566 | n8567;
  assign n8570 = ~n8568 & n8569;
  assign n13779 = n8343 | n8345;
  assign n16757 = n8570 & n13779;
  assign n16725 = n8110 | n8343;
  assign n16726 = (n8343 & n8345) | (n8343 & n16725) | (n8345 & n16725);
  assign n16758 = n8570 & n16726;
  assign n16759 = (n13598 & n16757) | (n13598 & n16758) | (n16757 & n16758);
  assign n16760 = n8570 | n13779;
  assign n16761 = n8570 | n16726;
  assign n16762 = (n13598 & n16760) | (n13598 & n16761) | (n16760 & n16761);
  assign n8573 = ~n16759 & n16762;
  assign n8574 = x74 & x89;
  assign n8575 = n8573 & n8574;
  assign n8576 = n8573 | n8574;
  assign n8577 = ~n8575 & n8576;
  assign n13776 = n8350 | n8352;
  assign n13808 = n8577 & n13776;
  assign n13809 = n8350 & n8577;
  assign n13810 = (n16656 & n13808) | (n16656 & n13809) | (n13808 & n13809);
  assign n13811 = n8577 | n13776;
  assign n13812 = n8350 | n8577;
  assign n13813 = (n16656 & n13811) | (n16656 & n13812) | (n13811 & n13812);
  assign n8580 = ~n13810 & n13813;
  assign n8581 = x73 & x90;
  assign n8582 = n8580 & n8581;
  assign n8583 = n8580 | n8581;
  assign n8584 = ~n8582 & n8583;
  assign n13814 = n8357 & n8584;
  assign n13815 = (n8584 & n16684) | (n8584 & n13814) | (n16684 & n13814);
  assign n13816 = n8357 | n8584;
  assign n13817 = n16684 | n13816;
  assign n8587 = ~n13815 & n13817;
  assign n8588 = x72 & x91;
  assign n8589 = n8587 & n8588;
  assign n8590 = n8587 | n8588;
  assign n8591 = ~n8589 & n8590;
  assign n8592 = n16724 & n8591;
  assign n8593 = n16724 | n8591;
  assign n8594 = ~n8592 & n8593;
  assign n8595 = x71 & x92;
  assign n8596 = n8594 & n8595;
  assign n8597 = n8594 | n8595;
  assign n8598 = ~n8596 & n8597;
  assign n13771 = n8371 | n8373;
  assign n13818 = n8598 & n13771;
  assign n13819 = n8371 & n8598;
  assign n13820 = (n13662 & n13818) | (n13662 & n13819) | (n13818 & n13819);
  assign n13821 = n8598 | n13771;
  assign n13822 = n8371 | n8598;
  assign n13823 = (n13662 & n13821) | (n13662 & n13822) | (n13821 & n13822);
  assign n8601 = ~n13820 & n13823;
  assign n8602 = x70 & x93;
  assign n8603 = n8601 & n8602;
  assign n8604 = n8601 | n8602;
  assign n8605 = ~n8603 & n8604;
  assign n13824 = n8378 & n8605;
  assign n13825 = (n8605 & n16702) | (n8605 & n13824) | (n16702 & n13824);
  assign n13826 = n8378 | n8605;
  assign n13827 = n16702 | n13826;
  assign n8608 = ~n13825 & n13827;
  assign n8609 = x69 & x94;
  assign n8610 = n8608 & n8609;
  assign n8611 = n8608 | n8609;
  assign n8612 = ~n8610 & n8611;
  assign n13828 = n8385 & n8612;
  assign n13829 = (n8612 & n13728) | (n8612 & n13828) | (n13728 & n13828);
  assign n13830 = n8385 | n8612;
  assign n13831 = n13728 | n13830;
  assign n8615 = ~n13829 & n13831;
  assign n8616 = x68 & x95;
  assign n8617 = n8615 & n8616;
  assign n8618 = n8615 | n8616;
  assign n8619 = ~n8617 & n8618;
  assign n13832 = n8392 & n8619;
  assign n13833 = (n8619 & n13732) | (n8619 & n13832) | (n13732 & n13832);
  assign n13834 = n8392 | n8619;
  assign n13835 = n13732 | n13834;
  assign n8622 = ~n13833 & n13835;
  assign n8623 = x67 & x96;
  assign n8624 = n8622 & n8623;
  assign n8625 = n8622 | n8623;
  assign n8626 = ~n8624 & n8625;
  assign n13836 = n8399 & n8626;
  assign n13837 = (n8626 & n13736) | (n8626 & n13836) | (n13736 & n13836);
  assign n13838 = n8399 | n8626;
  assign n13839 = n13736 | n13838;
  assign n8629 = ~n13837 & n13839;
  assign n8630 = x66 & x97;
  assign n8631 = n8629 & n8630;
  assign n8632 = n8629 | n8630;
  assign n8633 = ~n8631 & n8632;
  assign n13840 = n8406 & n8633;
  assign n13841 = (n8633 & n13741) | (n8633 & n13840) | (n13741 & n13840);
  assign n13842 = n8406 | n8633;
  assign n13843 = n13741 | n13842;
  assign n8636 = ~n13841 & n13843;
  assign n8637 = x65 & x98;
  assign n8638 = n8636 & n8637;
  assign n8639 = n8636 | n8637;
  assign n8640 = ~n8638 & n8639;
  assign n13769 = n8413 | n8415;
  assign n13844 = n8640 & n13769;
  assign n13845 = n8413 & n8640;
  assign n13846 = (n13657 & n13844) | (n13657 & n13845) | (n13844 & n13845);
  assign n13847 = n8640 | n13769;
  assign n13848 = n8413 | n8640;
  assign n13849 = (n13657 & n13847) | (n13657 & n13848) | (n13847 & n13848);
  assign n8643 = ~n13846 & n13849;
  assign n8644 = x64 & x99;
  assign n8645 = n8643 & n8644;
  assign n8646 = n8643 | n8644;
  assign n8647 = ~n8645 & n8646;
  assign n13767 = n8420 | n8422;
  assign n16763 = n8647 & n13767;
  assign n16764 = n8420 & n8647;
  assign n16765 = (n13655 & n16763) | (n13655 & n16764) | (n16763 & n16764);
  assign n16766 = n8647 | n13767;
  assign n16767 = n8420 | n8647;
  assign n16768 = (n13655 & n16766) | (n13655 & n16767) | (n16766 & n16767);
  assign n8650 = ~n16765 & n16768;
  assign n8651 = x63 & x100;
  assign n8652 = n8650 & n8651;
  assign n8653 = n8650 | n8651;
  assign n8654 = ~n8652 & n8653;
  assign n13765 = n8427 | n8429;
  assign n16769 = n8654 & n13765;
  assign n16770 = n8427 & n8654;
  assign n16771 = (n13653 & n16769) | (n13653 & n16770) | (n16769 & n16770);
  assign n16772 = n8654 | n13765;
  assign n16773 = n8427 | n8654;
  assign n16774 = (n13653 & n16772) | (n13653 & n16773) | (n16772 & n16773);
  assign n8657 = ~n16771 & n16774;
  assign n8658 = x62 & x101;
  assign n8659 = n8657 & n8658;
  assign n8660 = n8657 | n8658;
  assign n8661 = ~n8659 & n8660;
  assign n8662 = n13764 & n8661;
  assign n8663 = n13764 | n8661;
  assign n8664 = ~n8662 & n8663;
  assign n8665 = x61 & x102;
  assign n8666 = n8664 & n8665;
  assign n8667 = n8664 | n8665;
  assign n8668 = ~n8666 & n8667;
  assign n8669 = n13762 & n8668;
  assign n8670 = n13762 | n8668;
  assign n8671 = ~n8669 & n8670;
  assign n8672 = x60 & x103;
  assign n8673 = n8671 & n8672;
  assign n8674 = n8671 | n8672;
  assign n8675 = ~n8673 & n8674;
  assign n8676 = n13760 & n8675;
  assign n8677 = n13760 | n8675;
  assign n8678 = ~n8676 & n8677;
  assign n8679 = x59 & x104;
  assign n8680 = n8678 & n8679;
  assign n8681 = n8678 | n8679;
  assign n8682 = ~n8680 & n8681;
  assign n8683 = n13758 & n8682;
  assign n8684 = n13758 | n8682;
  assign n8685 = ~n8683 & n8684;
  assign n8686 = x58 & x105;
  assign n8687 = n8685 & n8686;
  assign n8688 = n8685 | n8686;
  assign n8689 = ~n8687 & n8688;
  assign n8690 = n13756 & n8689;
  assign n8691 = n13756 | n8689;
  assign n8692 = ~n8690 & n8691;
  assign n8693 = x57 & x106;
  assign n8694 = n8692 & n8693;
  assign n8695 = n8692 | n8693;
  assign n8696 = ~n8694 & n8695;
  assign n8697 = n13754 & n8696;
  assign n8698 = n13754 | n8696;
  assign n8699 = ~n8697 & n8698;
  assign n8700 = x56 & x107;
  assign n8701 = n8699 & n8700;
  assign n8702 = n8699 | n8700;
  assign n8703 = ~n8701 & n8702;
  assign n8704 = n16719 & n8703;
  assign n8705 = n16719 | n8703;
  assign n8706 = ~n8704 & n8705;
  assign n8707 = x55 & x108;
  assign n8708 = n8706 & n8707;
  assign n8709 = n8706 | n8707;
  assign n8710 = ~n8708 & n8709;
  assign n8711 = n13752 & n8710;
  assign n8712 = n13752 | n8710;
  assign n8713 = ~n8711 & n8712;
  assign n8714 = x54 & x109;
  assign n8715 = n8713 & n8714;
  assign n8716 = n8713 | n8714;
  assign n8717 = ~n8715 & n8716;
  assign n8718 = n13750 & n8717;
  assign n8719 = n13750 | n8717;
  assign n8720 = ~n8718 & n8719;
  assign n8721 = x53 & x110;
  assign n8722 = n8720 & n8721;
  assign n8723 = n8720 | n8721;
  assign n8724 = ~n8722 & n8723;
  assign n8725 = n13748 & n8724;
  assign n8726 = n13748 | n8724;
  assign n8727 = ~n8725 & n8726;
  assign n8728 = x52 & x111;
  assign n8729 = n8727 & n8728;
  assign n8730 = n8727 | n8728;
  assign n8731 = ~n8729 & n8730;
  assign n8732 = n13746 & n8731;
  assign n8733 = n13746 | n8731;
  assign n8734 = ~n8732 & n8733;
  assign n13850 = n8729 | n13746;
  assign n13851 = (n8729 & n8731) | (n8729 & n13850) | (n8731 & n13850);
  assign n13852 = n8722 | n13748;
  assign n13853 = (n8722 & n8724) | (n8722 & n13852) | (n8724 & n13852);
  assign n13854 = n8715 | n13750;
  assign n13855 = (n8715 & n8717) | (n8715 & n13854) | (n8717 & n13854);
  assign n13856 = n8708 | n13752;
  assign n13857 = (n8708 & n8710) | (n8708 & n13856) | (n8710 & n13856);
  assign n13858 = n8701 | n8703;
  assign n13859 = (n16719 & n8701) | (n16719 & n13858) | (n8701 & n13858);
  assign n13860 = n8694 | n8696;
  assign n13861 = (n8694 & n13754) | (n8694 & n13860) | (n13754 & n13860);
  assign n13862 = n8687 | n8689;
  assign n13863 = (n8687 & n13756) | (n8687 & n13862) | (n13756 & n13862);
  assign n13864 = n8680 | n8682;
  assign n13865 = (n8680 & n13758) | (n8680 & n13864) | (n13758 & n13864);
  assign n13866 = n8673 | n8675;
  assign n13867 = (n8673 & n13760) | (n8673 & n13866) | (n13760 & n13866);
  assign n13868 = n8666 | n8668;
  assign n13869 = (n8666 & n13762) | (n8666 & n13868) | (n13762 & n13868);
  assign n13766 = (n8427 & n13653) | (n8427 & n13765) | (n13653 & n13765);
  assign n13768 = (n8420 & n13655) | (n8420 & n13767) | (n13655 & n13767);
  assign n13780 = (n13598 & n16726) | (n13598 & n13779) | (n16726 & n13779);
  assign n13887 = n8561 | n8563;
  assign n16779 = n8336 | n8561;
  assign n16780 = (n8561 & n8563) | (n8561 & n16779) | (n8563 & n16779);
  assign n16781 = (n13703 & n13887) | (n13703 & n16780) | (n13887 & n16780);
  assign n16782 = (n13704 & n13887) | (n13704 & n16780) | (n13887 & n16780);
  assign n16783 = (n13557 & n16781) | (n13557 & n16782) | (n16781 & n16782);
  assign n13782 = n8329 | n13697;
  assign n8763 = x79 & x85;
  assign n66379 = n8763 & n49973;
  assign n66380 = n8763 & n49971;
  assign n66381 = (n16508 & n66379) | (n16508 & n66380) | (n66379 & n66380);
  assign n49984 = (n8763 & n16742) | (n8763 & n66381) | (n16742 & n66381);
  assign n49983 = n8763 & n16735;
  assign n66382 = (n8542 & n8763) | (n8542 & n49983) | (n8763 & n49983);
  assign n49986 = (n16740 & n66381) | (n16740 & n66382) | (n66381 & n66382);
  assign n16792 = (n16602 & n49984) | (n16602 & n49986) | (n49984 & n49986);
  assign n66383 = n8763 | n49973;
  assign n66384 = n8763 | n49971;
  assign n66385 = (n16508 & n66383) | (n16508 & n66384) | (n66383 & n66384);
  assign n49988 = n16742 | n66385;
  assign n49987 = n8763 | n16735;
  assign n66386 = n8542 | n49987;
  assign n49990 = (n16740 & n66385) | (n16740 & n66386) | (n66385 & n66386);
  assign n16795 = (n16602 & n49988) | (n16602 & n49990) | (n49988 & n49990);
  assign n8766 = ~n16792 & n16795;
  assign n16784 = n8547 | n8549;
  assign n16785 = (n8547 & n13784) | (n8547 & n16784) | (n13784 & n16784);
  assign n16796 = n8766 & n16785;
  assign n16786 = n8322 | n8547;
  assign n16787 = (n8547 & n8549) | (n8547 & n16786) | (n8549 & n16786);
  assign n16797 = n8766 & n16787;
  assign n16798 = (n16663 & n16796) | (n16663 & n16797) | (n16796 & n16797);
  assign n16799 = n8766 | n16785;
  assign n16800 = n8766 | n16787;
  assign n16801 = (n16663 & n16799) | (n16663 & n16800) | (n16799 & n16800);
  assign n8769 = ~n16798 & n16801;
  assign n8770 = x78 & x86;
  assign n8771 = n8769 & n8770;
  assign n8772 = n8769 | n8770;
  assign n8773 = ~n8771 & n8772;
  assign n13889 = n8554 | n8556;
  assign n13897 = n8773 & n13889;
  assign n13898 = n8554 & n8773;
  assign n16802 = (n13782 & n13897) | (n13782 & n13898) | (n13897 & n13898);
  assign n16803 = (n13897 & n13898) | (n13897 & n16728) | (n13898 & n16728);
  assign n16804 = (n13560 & n16802) | (n13560 & n16803) | (n16802 & n16803);
  assign n13900 = n8773 | n13889;
  assign n13901 = n8554 | n8773;
  assign n16805 = (n13782 & n13900) | (n13782 & n13901) | (n13900 & n13901);
  assign n16806 = (n13900 & n13901) | (n13900 & n16728) | (n13901 & n16728);
  assign n16807 = (n13560 & n16805) | (n13560 & n16806) | (n16805 & n16806);
  assign n8776 = ~n16804 & n16807;
  assign n8777 = x77 & x87;
  assign n8778 = n8776 & n8777;
  assign n8779 = n8776 | n8777;
  assign n8780 = ~n8778 & n8779;
  assign n8781 = n16783 & n8780;
  assign n8782 = n16783 | n8780;
  assign n8783 = ~n8781 & n8782;
  assign n8784 = x76 & x88;
  assign n8785 = n8783 & n8784;
  assign n8786 = n8783 | n8784;
  assign n8787 = ~n8785 & n8786;
  assign n13884 = n8568 | n8570;
  assign n13903 = n8787 & n13884;
  assign n13904 = n8568 & n8787;
  assign n13905 = (n13780 & n13903) | (n13780 & n13904) | (n13903 & n13904);
  assign n13906 = n8787 | n13884;
  assign n13907 = n8568 | n8787;
  assign n13908 = (n13780 & n13906) | (n13780 & n13907) | (n13906 & n13907);
  assign n8790 = ~n13905 & n13908;
  assign n8791 = x75 & x89;
  assign n8792 = n8790 & n8791;
  assign n8793 = n8790 | n8791;
  assign n8794 = ~n8792 & n8793;
  assign n13909 = n8575 & n8794;
  assign n13910 = (n8794 & n13810) | (n8794 & n13909) | (n13810 & n13909);
  assign n13911 = n8575 | n8794;
  assign n13912 = n13810 | n13911;
  assign n8797 = ~n13910 & n13912;
  assign n8798 = x74 & x90;
  assign n8799 = n8797 & n8798;
  assign n8800 = n8797 | n8798;
  assign n8801 = ~n8799 & n8800;
  assign n13882 = n8582 | n8584;
  assign n16808 = n8801 & n13882;
  assign n16777 = n8357 | n8582;
  assign n16778 = (n8582 & n8584) | (n8582 & n16777) | (n8584 & n16777);
  assign n16809 = n8801 & n16778;
  assign n16810 = (n16684 & n16808) | (n16684 & n16809) | (n16808 & n16809);
  assign n16811 = n8801 | n13882;
  assign n16812 = n8801 | n16778;
  assign n16813 = (n16684 & n16811) | (n16684 & n16812) | (n16811 & n16812);
  assign n8804 = ~n16810 & n16813;
  assign n8805 = x73 & x91;
  assign n8806 = n8804 & n8805;
  assign n8807 = n8804 | n8805;
  assign n8808 = ~n8806 & n8807;
  assign n13879 = n8589 | n8591;
  assign n13913 = n8808 & n13879;
  assign n13914 = n8589 & n8808;
  assign n13915 = (n16724 & n13913) | (n16724 & n13914) | (n13913 & n13914);
  assign n13916 = n8808 | n13879;
  assign n13917 = n8589 | n8808;
  assign n13918 = (n16724 & n13916) | (n16724 & n13917) | (n13916 & n13917);
  assign n8811 = ~n13915 & n13918;
  assign n8812 = x72 & x92;
  assign n8813 = n8811 & n8812;
  assign n8814 = n8811 | n8812;
  assign n8815 = ~n8813 & n8814;
  assign n13919 = n8596 & n8815;
  assign n16814 = (n8815 & n13819) | (n8815 & n13919) | (n13819 & n13919);
  assign n16815 = (n8815 & n13818) | (n8815 & n13919) | (n13818 & n13919);
  assign n16816 = (n13662 & n16814) | (n13662 & n16815) | (n16814 & n16815);
  assign n13921 = n8596 | n8815;
  assign n16817 = n13819 | n13921;
  assign n16818 = n13818 | n13921;
  assign n16819 = (n13662 & n16817) | (n13662 & n16818) | (n16817 & n16818);
  assign n8818 = ~n16816 & n16819;
  assign n8819 = x71 & x93;
  assign n8820 = n8818 & n8819;
  assign n8821 = n8818 | n8819;
  assign n8822 = ~n8820 & n8821;
  assign n13877 = n8603 | n8605;
  assign n16820 = n8822 & n13877;
  assign n16775 = n8378 | n8603;
  assign n16776 = (n8603 & n8605) | (n8603 & n16775) | (n8605 & n16775);
  assign n16821 = n8822 & n16776;
  assign n16822 = (n16702 & n16820) | (n16702 & n16821) | (n16820 & n16821);
  assign n16823 = n8822 | n13877;
  assign n16824 = n8822 | n16776;
  assign n16825 = (n16702 & n16823) | (n16702 & n16824) | (n16823 & n16824);
  assign n8825 = ~n16822 & n16825;
  assign n8826 = x70 & x94;
  assign n8827 = n8825 & n8826;
  assign n8828 = n8825 | n8826;
  assign n8829 = ~n8827 & n8828;
  assign n13923 = n8610 & n8829;
  assign n16826 = (n8829 & n13828) | (n8829 & n13923) | (n13828 & n13923);
  assign n16827 = (n8612 & n8829) | (n8612 & n13923) | (n8829 & n13923);
  assign n16828 = (n13728 & n16826) | (n13728 & n16827) | (n16826 & n16827);
  assign n13925 = n8610 | n8829;
  assign n16829 = n13828 | n13925;
  assign n16830 = n8612 | n13925;
  assign n16831 = (n13728 & n16829) | (n13728 & n16830) | (n16829 & n16830);
  assign n8832 = ~n16828 & n16831;
  assign n8833 = x69 & x95;
  assign n8834 = n8832 & n8833;
  assign n8835 = n8832 | n8833;
  assign n8836 = ~n8834 & n8835;
  assign n13927 = n8617 & n8836;
  assign n13928 = (n8836 & n13833) | (n8836 & n13927) | (n13833 & n13927);
  assign n13929 = n8617 | n8836;
  assign n13930 = n13833 | n13929;
  assign n8839 = ~n13928 & n13930;
  assign n8840 = x68 & x96;
  assign n8841 = n8839 & n8840;
  assign n8842 = n8839 | n8840;
  assign n8843 = ~n8841 & n8842;
  assign n13931 = n8624 & n8843;
  assign n13932 = (n8843 & n13837) | (n8843 & n13931) | (n13837 & n13931);
  assign n13933 = n8624 | n8843;
  assign n13934 = n13837 | n13933;
  assign n8846 = ~n13932 & n13934;
  assign n8847 = x67 & x97;
  assign n8848 = n8846 & n8847;
  assign n8849 = n8846 | n8847;
  assign n8850 = ~n8848 & n8849;
  assign n13935 = n8631 & n8850;
  assign n13936 = (n8850 & n13841) | (n8850 & n13935) | (n13841 & n13935);
  assign n13937 = n8631 | n8850;
  assign n13938 = n13841 | n13937;
  assign n8853 = ~n13936 & n13938;
  assign n8854 = x66 & x98;
  assign n8855 = n8853 & n8854;
  assign n8856 = n8853 | n8854;
  assign n8857 = ~n8855 & n8856;
  assign n13939 = n8638 & n8857;
  assign n13940 = (n8857 & n13846) | (n8857 & n13939) | (n13846 & n13939);
  assign n13941 = n8638 | n8857;
  assign n13942 = n13846 | n13941;
  assign n8860 = ~n13940 & n13942;
  assign n8861 = x65 & x99;
  assign n8862 = n8860 & n8861;
  assign n8863 = n8860 | n8861;
  assign n8864 = ~n8862 & n8863;
  assign n13874 = n8645 | n8647;
  assign n13943 = n8864 & n13874;
  assign n13944 = n8645 & n8864;
  assign n13945 = (n13768 & n13943) | (n13768 & n13944) | (n13943 & n13944);
  assign n13946 = n8864 | n13874;
  assign n13947 = n8645 | n8864;
  assign n13948 = (n13768 & n13946) | (n13768 & n13947) | (n13946 & n13947);
  assign n8867 = ~n13945 & n13948;
  assign n8868 = x64 & x100;
  assign n8869 = n8867 & n8868;
  assign n8870 = n8867 | n8868;
  assign n8871 = ~n8869 & n8870;
  assign n13872 = n8652 | n8654;
  assign n16832 = n8871 & n13872;
  assign n16833 = n8652 & n8871;
  assign n16834 = (n13766 & n16832) | (n13766 & n16833) | (n16832 & n16833);
  assign n16835 = n8871 | n13872;
  assign n16836 = n8652 | n8871;
  assign n16837 = (n13766 & n16835) | (n13766 & n16836) | (n16835 & n16836);
  assign n8874 = ~n16834 & n16837;
  assign n8875 = x63 & x101;
  assign n8876 = n8874 & n8875;
  assign n8877 = n8874 | n8875;
  assign n8878 = ~n8876 & n8877;
  assign n13870 = n8659 | n8661;
  assign n16838 = n8878 & n13870;
  assign n16839 = n8659 & n8878;
  assign n16840 = (n13764 & n16838) | (n13764 & n16839) | (n16838 & n16839);
  assign n16841 = n8878 | n13870;
  assign n16842 = n8659 | n8878;
  assign n16843 = (n13764 & n16841) | (n13764 & n16842) | (n16841 & n16842);
  assign n8881 = ~n16840 & n16843;
  assign n8882 = x62 & x102;
  assign n8883 = n8881 & n8882;
  assign n8884 = n8881 | n8882;
  assign n8885 = ~n8883 & n8884;
  assign n8886 = n13869 & n8885;
  assign n8887 = n13869 | n8885;
  assign n8888 = ~n8886 & n8887;
  assign n8889 = x61 & x103;
  assign n8890 = n8888 & n8889;
  assign n8891 = n8888 | n8889;
  assign n8892 = ~n8890 & n8891;
  assign n8893 = n13867 & n8892;
  assign n8894 = n13867 | n8892;
  assign n8895 = ~n8893 & n8894;
  assign n8896 = x60 & x104;
  assign n8897 = n8895 & n8896;
  assign n8898 = n8895 | n8896;
  assign n8899 = ~n8897 & n8898;
  assign n8900 = n13865 & n8899;
  assign n8901 = n13865 | n8899;
  assign n8902 = ~n8900 & n8901;
  assign n8903 = x59 & x105;
  assign n8904 = n8902 & n8903;
  assign n8905 = n8902 | n8903;
  assign n8906 = ~n8904 & n8905;
  assign n8907 = n13863 & n8906;
  assign n8908 = n13863 | n8906;
  assign n8909 = ~n8907 & n8908;
  assign n8910 = x58 & x106;
  assign n8911 = n8909 & n8910;
  assign n8912 = n8909 | n8910;
  assign n8913 = ~n8911 & n8912;
  assign n8914 = n13861 & n8913;
  assign n8915 = n13861 | n8913;
  assign n8916 = ~n8914 & n8915;
  assign n8917 = x57 & x107;
  assign n8918 = n8916 & n8917;
  assign n8919 = n8916 | n8917;
  assign n8920 = ~n8918 & n8919;
  assign n8921 = n13859 & n8920;
  assign n8922 = n13859 | n8920;
  assign n8923 = ~n8921 & n8922;
  assign n8924 = x56 & x108;
  assign n8925 = n8923 & n8924;
  assign n8926 = n8923 | n8924;
  assign n8927 = ~n8925 & n8926;
  assign n8928 = n13857 & n8927;
  assign n8929 = n13857 | n8927;
  assign n8930 = ~n8928 & n8929;
  assign n8931 = x55 & x109;
  assign n8932 = n8930 & n8931;
  assign n8933 = n8930 | n8931;
  assign n8934 = ~n8932 & n8933;
  assign n8935 = n13855 & n8934;
  assign n8936 = n13855 | n8934;
  assign n8937 = ~n8935 & n8936;
  assign n8938 = x54 & x110;
  assign n8939 = n8937 & n8938;
  assign n8940 = n8937 | n8938;
  assign n8941 = ~n8939 & n8940;
  assign n8942 = n13853 & n8941;
  assign n8943 = n13853 | n8941;
  assign n8944 = ~n8942 & n8943;
  assign n8945 = x53 & x111;
  assign n8946 = n8944 & n8945;
  assign n8947 = n8944 | n8945;
  assign n8948 = ~n8946 & n8947;
  assign n8949 = n13851 & n8948;
  assign n8950 = n13851 | n8948;
  assign n8951 = ~n8949 & n8950;
  assign n8952 = n8946 | n8949;
  assign n8953 = n8939 | n8942;
  assign n8954 = n8932 | n8935;
  assign n8955 = n8925 | n8928;
  assign n13949 = n8918 | n8920;
  assign n13950 = (n8918 & n13859) | (n8918 & n13949) | (n13859 & n13949);
  assign n13951 = n8911 | n8913;
  assign n13952 = (n8911 & n13861) | (n8911 & n13951) | (n13861 & n13951);
  assign n13953 = n8904 | n8906;
  assign n13954 = (n8904 & n13863) | (n8904 & n13953) | (n13863 & n13953);
  assign n13955 = n8897 | n8899;
  assign n13956 = (n8897 & n13865) | (n8897 & n13955) | (n13865 & n13955);
  assign n13957 = n8890 | n8892;
  assign n13958 = (n8890 & n13867) | (n8890 & n13957) | (n13867 & n13957);
  assign n13871 = (n8659 & n13764) | (n8659 & n13870) | (n13764 & n13870);
  assign n13873 = (n8652 & n13766) | (n8652 & n13872) | (n13766 & n13872);
  assign n13878 = (n16702 & n16776) | (n16702 & n13877) | (n16776 & n13877);
  assign n13968 = n8813 | n8815;
  assign n16844 = n8596 | n8813;
  assign n16845 = (n8813 & n8815) | (n8813 & n16844) | (n8815 & n16844);
  assign n16846 = (n13819 & n13968) | (n13819 & n16845) | (n13968 & n16845);
  assign n16847 = (n13818 & n13968) | (n13818 & n16845) | (n13968 & n16845);
  assign n16848 = (n13662 & n16846) | (n13662 & n16847) | (n16846 & n16847);
  assign n13883 = (n16684 & n16778) | (n16684 & n13882) | (n16778 & n13882);
  assign n16851 = n8554 | n8771;
  assign n16852 = (n8771 & n8773) | (n8771 & n16851) | (n8773 & n16851);
  assign n16853 = n8771 | n8773;
  assign n16854 = (n8771 & n13889) | (n8771 & n16853) | (n13889 & n16853);
  assign n16855 = (n13782 & n16852) | (n13782 & n16854) | (n16852 & n16854);
  assign n16856 = (n16728 & n16852) | (n16728 & n16854) | (n16852 & n16854);
  assign n16857 = (n13560 & n16855) | (n13560 & n16856) | (n16855 & n16856);
  assign n8979 = x79 & x86;
  assign n66387 = n8979 & n66382;
  assign n66388 = n8979 & n66381;
  assign n66389 = (n16740 & n66387) | (n16740 & n66388) | (n66387 & n66388);
  assign n49997 = n8763 & n8979;
  assign n66390 = (n16742 & n49997) | (n16742 & n66388) | (n49997 & n66388);
  assign n49993 = (n16602 & n66389) | (n16602 & n66390) | (n66389 & n66390);
  assign n16859 = (n8766 & n8979) | (n8766 & n49993) | (n8979 & n49993);
  assign n49994 = n8979 & n66382;
  assign n66391 = n8979 & n66380;
  assign n66392 = n8979 & n66379;
  assign n66393 = (n16508 & n66391) | (n16508 & n66392) | (n66391 & n66392);
  assign n49996 = (n16740 & n49994) | (n16740 & n66393) | (n49994 & n66393);
  assign n49998 = (n16742 & n66393) | (n16742 & n49997) | (n66393 & n49997);
  assign n16862 = (n16602 & n49996) | (n16602 & n49998) | (n49996 & n49998);
  assign n16863 = (n16785 & n16859) | (n16785 & n16862) | (n16859 & n16862);
  assign n16864 = (n16787 & n16859) | (n16787 & n16862) | (n16859 & n16862);
  assign n16865 = (n16663 & n16863) | (n16663 & n16864) | (n16863 & n16864);
  assign n66394 = n8979 | n66382;
  assign n66395 = n8979 | n66381;
  assign n66396 = (n16740 & n66394) | (n16740 & n66395) | (n66394 & n66395);
  assign n50005 = n8763 | n8979;
  assign n66397 = (n16742 & n50005) | (n16742 & n66395) | (n50005 & n66395);
  assign n50001 = (n16602 & n66396) | (n16602 & n66397) | (n66396 & n66397);
  assign n16867 = n8766 | n50001;
  assign n50002 = n8979 | n66382;
  assign n66398 = n8979 | n66380;
  assign n66399 = n8979 | n66379;
  assign n66400 = (n16508 & n66398) | (n16508 & n66399) | (n66398 & n66399);
  assign n50004 = (n16740 & n50002) | (n16740 & n66400) | (n50002 & n66400);
  assign n50006 = (n16742 & n66400) | (n16742 & n50005) | (n66400 & n50005);
  assign n16870 = (n16602 & n50004) | (n16602 & n50006) | (n50004 & n50006);
  assign n16871 = (n16785 & n16867) | (n16785 & n16870) | (n16867 & n16870);
  assign n16872 = (n16787 & n16867) | (n16787 & n16870) | (n16867 & n16870);
  assign n16873 = (n16663 & n16871) | (n16663 & n16872) | (n16871 & n16872);
  assign n8982 = ~n16865 & n16873;
  assign n8983 = n16857 & n8982;
  assign n8984 = n16857 | n8982;
  assign n8985 = ~n8983 & n8984;
  assign n8986 = x78 & x87;
  assign n8987 = n8985 & n8986;
  assign n8988 = n8985 | n8986;
  assign n8989 = ~n8987 & n8988;
  assign n13975 = n8778 | n8780;
  assign n13988 = n8989 & n13975;
  assign n13989 = n8778 & n8989;
  assign n13990 = (n16783 & n13988) | (n16783 & n13989) | (n13988 & n13989);
  assign n13991 = n8989 | n13975;
  assign n13992 = n8778 | n8989;
  assign n13993 = (n16783 & n13991) | (n16783 & n13992) | (n13991 & n13992);
  assign n8992 = ~n13990 & n13993;
  assign n8993 = x77 & x88;
  assign n8994 = n8992 & n8993;
  assign n8995 = n8992 | n8993;
  assign n8996 = ~n8994 & n8995;
  assign n13994 = n8785 & n8996;
  assign n16874 = (n8996 & n13904) | (n8996 & n13994) | (n13904 & n13994);
  assign n16875 = (n8996 & n13903) | (n8996 & n13994) | (n13903 & n13994);
  assign n16876 = (n13780 & n16874) | (n13780 & n16875) | (n16874 & n16875);
  assign n13996 = n8785 | n8996;
  assign n16877 = n13904 | n13996;
  assign n16878 = n13903 | n13996;
  assign n16879 = (n13780 & n16877) | (n13780 & n16878) | (n16877 & n16878);
  assign n8999 = ~n16876 & n16879;
  assign n9000 = x76 & x89;
  assign n9001 = n8999 & n9000;
  assign n9002 = n8999 | n9000;
  assign n9003 = ~n9001 & n9002;
  assign n13973 = n8792 | n8794;
  assign n16880 = n9003 & n13973;
  assign n16849 = n8575 | n8792;
  assign n16850 = (n8792 & n8794) | (n8792 & n16849) | (n8794 & n16849);
  assign n16881 = n9003 & n16850;
  assign n16882 = (n13810 & n16880) | (n13810 & n16881) | (n16880 & n16881);
  assign n16883 = n9003 | n13973;
  assign n16884 = n9003 | n16850;
  assign n16885 = (n13810 & n16883) | (n13810 & n16884) | (n16883 & n16884);
  assign n9006 = ~n16882 & n16885;
  assign n9007 = x75 & x90;
  assign n9008 = n9006 & n9007;
  assign n9009 = n9006 | n9007;
  assign n9010 = ~n9008 & n9009;
  assign n13970 = n8799 | n8801;
  assign n13998 = n9010 & n13970;
  assign n13999 = n8799 & n9010;
  assign n14000 = (n13883 & n13998) | (n13883 & n13999) | (n13998 & n13999);
  assign n14001 = n9010 | n13970;
  assign n14002 = n8799 | n9010;
  assign n14003 = (n13883 & n14001) | (n13883 & n14002) | (n14001 & n14002);
  assign n9013 = ~n14000 & n14003;
  assign n9014 = x74 & x91;
  assign n9015 = n9013 & n9014;
  assign n9016 = n9013 | n9014;
  assign n9017 = ~n9015 & n9016;
  assign n14004 = n8806 & n9017;
  assign n16886 = (n9017 & n13913) | (n9017 & n14004) | (n13913 & n14004);
  assign n16887 = (n9017 & n13914) | (n9017 & n14004) | (n13914 & n14004);
  assign n16888 = (n16724 & n16886) | (n16724 & n16887) | (n16886 & n16887);
  assign n14006 = n8806 | n9017;
  assign n16889 = n13913 | n14006;
  assign n16890 = n13914 | n14006;
  assign n16891 = (n16724 & n16889) | (n16724 & n16890) | (n16889 & n16890);
  assign n9020 = ~n16888 & n16891;
  assign n9021 = x73 & x92;
  assign n9022 = n9020 & n9021;
  assign n9023 = n9020 | n9021;
  assign n9024 = ~n9022 & n9023;
  assign n9025 = n16848 & n9024;
  assign n9026 = n16848 | n9024;
  assign n9027 = ~n9025 & n9026;
  assign n9028 = x72 & x93;
  assign n9029 = n9027 & n9028;
  assign n9030 = n9027 | n9028;
  assign n9031 = ~n9029 & n9030;
  assign n13965 = n8820 | n8822;
  assign n14008 = n9031 & n13965;
  assign n14009 = n8820 & n9031;
  assign n14010 = (n13878 & n14008) | (n13878 & n14009) | (n14008 & n14009);
  assign n14011 = n9031 | n13965;
  assign n14012 = n8820 | n9031;
  assign n14013 = (n13878 & n14011) | (n13878 & n14012) | (n14011 & n14012);
  assign n9034 = ~n14010 & n14013;
  assign n9035 = x71 & x94;
  assign n9036 = n9034 & n9035;
  assign n9037 = n9034 | n9035;
  assign n9038 = ~n9036 & n9037;
  assign n14014 = n8827 & n9038;
  assign n14015 = (n9038 & n16828) | (n9038 & n14014) | (n16828 & n14014);
  assign n14016 = n8827 | n9038;
  assign n14017 = n16828 | n14016;
  assign n9041 = ~n14015 & n14017;
  assign n9042 = x70 & x95;
  assign n9043 = n9041 & n9042;
  assign n9044 = n9041 | n9042;
  assign n9045 = ~n9043 & n9044;
  assign n14018 = n8834 & n9045;
  assign n14019 = (n9045 & n13928) | (n9045 & n14018) | (n13928 & n14018);
  assign n14020 = n8834 | n9045;
  assign n14021 = n13928 | n14020;
  assign n9048 = ~n14019 & n14021;
  assign n9049 = x69 & x96;
  assign n9050 = n9048 & n9049;
  assign n9051 = n9048 | n9049;
  assign n9052 = ~n9050 & n9051;
  assign n14022 = n8841 & n9052;
  assign n14023 = (n9052 & n13932) | (n9052 & n14022) | (n13932 & n14022);
  assign n14024 = n8841 | n9052;
  assign n14025 = n13932 | n14024;
  assign n9055 = ~n14023 & n14025;
  assign n9056 = x68 & x97;
  assign n9057 = n9055 & n9056;
  assign n9058 = n9055 | n9056;
  assign n9059 = ~n9057 & n9058;
  assign n14026 = n8848 & n9059;
  assign n14027 = (n9059 & n13936) | (n9059 & n14026) | (n13936 & n14026);
  assign n14028 = n8848 | n9059;
  assign n14029 = n13936 | n14028;
  assign n9062 = ~n14027 & n14029;
  assign n9063 = x67 & x98;
  assign n9064 = n9062 & n9063;
  assign n9065 = n9062 | n9063;
  assign n9066 = ~n9064 & n9065;
  assign n14030 = n8855 & n9066;
  assign n14031 = (n9066 & n13940) | (n9066 & n14030) | (n13940 & n14030);
  assign n14032 = n8855 | n9066;
  assign n14033 = n13940 | n14032;
  assign n9069 = ~n14031 & n14033;
  assign n9070 = x66 & x99;
  assign n9071 = n9069 & n9070;
  assign n9072 = n9069 | n9070;
  assign n9073 = ~n9071 & n9072;
  assign n14034 = n8862 & n9073;
  assign n14035 = (n9073 & n13945) | (n9073 & n14034) | (n13945 & n14034);
  assign n14036 = n8862 | n9073;
  assign n14037 = n13945 | n14036;
  assign n9076 = ~n14035 & n14037;
  assign n9077 = x65 & x100;
  assign n9078 = n9076 & n9077;
  assign n9079 = n9076 | n9077;
  assign n9080 = ~n9078 & n9079;
  assign n13963 = n8869 | n8871;
  assign n14038 = n9080 & n13963;
  assign n14039 = n8869 & n9080;
  assign n14040 = (n13873 & n14038) | (n13873 & n14039) | (n14038 & n14039);
  assign n14041 = n9080 | n13963;
  assign n14042 = n8869 | n9080;
  assign n14043 = (n13873 & n14041) | (n13873 & n14042) | (n14041 & n14042);
  assign n9083 = ~n14040 & n14043;
  assign n9084 = x64 & x101;
  assign n9085 = n9083 & n9084;
  assign n9086 = n9083 | n9084;
  assign n9087 = ~n9085 & n9086;
  assign n13961 = n8876 | n8878;
  assign n16892 = n9087 & n13961;
  assign n16893 = n8876 & n9087;
  assign n16894 = (n13871 & n16892) | (n13871 & n16893) | (n16892 & n16893);
  assign n16895 = n9087 | n13961;
  assign n16896 = n8876 | n9087;
  assign n16897 = (n13871 & n16895) | (n13871 & n16896) | (n16895 & n16896);
  assign n9090 = ~n16894 & n16897;
  assign n9091 = x63 & x102;
  assign n9092 = n9090 & n9091;
  assign n9093 = n9090 | n9091;
  assign n9094 = ~n9092 & n9093;
  assign n13959 = n8883 | n8885;
  assign n16898 = n9094 & n13959;
  assign n16899 = n8883 & n9094;
  assign n16900 = (n13869 & n16898) | (n13869 & n16899) | (n16898 & n16899);
  assign n16901 = n9094 | n13959;
  assign n16902 = n8883 | n9094;
  assign n16903 = (n13869 & n16901) | (n13869 & n16902) | (n16901 & n16902);
  assign n9097 = ~n16900 & n16903;
  assign n9098 = x62 & x103;
  assign n9099 = n9097 & n9098;
  assign n9100 = n9097 | n9098;
  assign n9101 = ~n9099 & n9100;
  assign n9102 = n13958 & n9101;
  assign n9103 = n13958 | n9101;
  assign n9104 = ~n9102 & n9103;
  assign n9105 = x61 & x104;
  assign n9106 = n9104 & n9105;
  assign n9107 = n9104 | n9105;
  assign n9108 = ~n9106 & n9107;
  assign n9109 = n13956 & n9108;
  assign n9110 = n13956 | n9108;
  assign n9111 = ~n9109 & n9110;
  assign n9112 = x60 & x105;
  assign n9113 = n9111 & n9112;
  assign n9114 = n9111 | n9112;
  assign n9115 = ~n9113 & n9114;
  assign n9116 = n13954 & n9115;
  assign n9117 = n13954 | n9115;
  assign n9118 = ~n9116 & n9117;
  assign n9119 = x59 & x106;
  assign n9120 = n9118 & n9119;
  assign n9121 = n9118 | n9119;
  assign n9122 = ~n9120 & n9121;
  assign n9123 = n13952 & n9122;
  assign n9124 = n13952 | n9122;
  assign n9125 = ~n9123 & n9124;
  assign n9126 = x58 & x107;
  assign n9127 = n9125 & n9126;
  assign n9128 = n9125 | n9126;
  assign n9129 = ~n9127 & n9128;
  assign n9130 = n13950 & n9129;
  assign n9131 = n13950 | n9129;
  assign n9132 = ~n9130 & n9131;
  assign n9133 = x57 & x108;
  assign n9134 = n9132 & n9133;
  assign n9135 = n9132 | n9133;
  assign n9136 = ~n9134 & n9135;
  assign n9137 = n8955 & n9136;
  assign n9138 = n8955 | n9136;
  assign n9139 = ~n9137 & n9138;
  assign n9140 = x56 & x109;
  assign n9141 = n9139 & n9140;
  assign n9142 = n9139 | n9140;
  assign n9143 = ~n9141 & n9142;
  assign n9144 = n8954 & n9143;
  assign n9145 = n8954 | n9143;
  assign n9146 = ~n9144 & n9145;
  assign n9147 = x55 & x110;
  assign n9148 = n9146 & n9147;
  assign n9149 = n9146 | n9147;
  assign n9150 = ~n9148 & n9149;
  assign n9151 = n8953 & n9150;
  assign n9152 = n8953 | n9150;
  assign n9153 = ~n9151 & n9152;
  assign n9154 = x54 & x111;
  assign n9155 = n9153 & n9154;
  assign n9156 = n9153 | n9154;
  assign n9157 = ~n9155 & n9156;
  assign n9158 = n8952 & n9157;
  assign n9159 = n8952 | n9157;
  assign n9160 = ~n9158 & n9159;
  assign n9161 = n9155 | n9158;
  assign n9162 = n9148 | n9151;
  assign n9163 = n9141 | n9144;
  assign n14044 = n9134 | n9136;
  assign n14045 = (n8955 & n9134) | (n8955 & n14044) | (n9134 & n14044);
  assign n14046 = n9127 | n9129;
  assign n14047 = (n9127 & n13950) | (n9127 & n14046) | (n13950 & n14046);
  assign n14048 = n9120 | n9122;
  assign n14049 = (n9120 & n13952) | (n9120 & n14048) | (n13952 & n14048);
  assign n14050 = n9113 | n9115;
  assign n14051 = (n9113 & n13954) | (n9113 & n14050) | (n13954 & n14050);
  assign n14052 = n9106 | n9108;
  assign n14053 = (n9106 & n13956) | (n9106 & n14052) | (n13956 & n14052);
  assign n13960 = (n8883 & n13869) | (n8883 & n13959) | (n13869 & n13959);
  assign n13962 = (n8876 & n13871) | (n8876 & n13961) | (n13871 & n13961);
  assign n14066 = n9015 | n9017;
  assign n16906 = n8806 | n9015;
  assign n16907 = (n9015 & n9017) | (n9015 & n16906) | (n9017 & n16906);
  assign n16908 = (n13913 & n14066) | (n13913 & n16907) | (n14066 & n16907);
  assign n16909 = (n13914 & n14066) | (n13914 & n16907) | (n14066 & n16907);
  assign n16910 = (n16724 & n16908) | (n16724 & n16909) | (n16908 & n16909);
  assign n13974 = (n13810 & n16850) | (n13810 & n13973) | (n16850 & n13973);
  assign n14071 = n8994 | n8996;
  assign n16911 = n8785 | n8994;
  assign n16912 = (n8994 & n8996) | (n8994 & n16911) | (n8996 & n16911);
  assign n16913 = (n13904 & n14071) | (n13904 & n16912) | (n14071 & n16912);
  assign n16914 = (n13903 & n14071) | (n13903 & n16912) | (n14071 & n16912);
  assign n16915 = (n13780 & n16913) | (n13780 & n16914) | (n16913 & n16914);
  assign n16916 = n8778 | n8987;
  assign n16917 = (n8987 & n8989) | (n8987 & n16916) | (n8989 & n16916);
  assign n14074 = n8987 | n13988;
  assign n14075 = (n16783 & n16917) | (n16783 & n14074) | (n16917 & n14074);
  assign n9187 = x79 & x87;
  assign n16918 = n9187 & n16865;
  assign n16919 = (n8982 & n9187) | (n8982 & n16918) | (n9187 & n16918);
  assign n14079 = n9187 & n16865;
  assign n14080 = (n16857 & n16919) | (n16857 & n14079) | (n16919 & n14079);
  assign n16920 = n9187 | n16865;
  assign n16921 = n8982 | n16920;
  assign n14082 = n9187 | n16865;
  assign n14083 = (n16857 & n16921) | (n16857 & n14082) | (n16921 & n14082);
  assign n9190 = ~n14080 & n14083;
  assign n9191 = n14075 & n9190;
  assign n9192 = n14075 | n9190;
  assign n9193 = ~n9191 & n9192;
  assign n9194 = x78 & x88;
  assign n9195 = n9193 & n9194;
  assign n9196 = n9193 | n9194;
  assign n9197 = ~n9195 & n9196;
  assign n9198 = n16915 & n9197;
  assign n9199 = n16915 | n9197;
  assign n9200 = ~n9198 & n9199;
  assign n9201 = x77 & x89;
  assign n9202 = n9200 & n9201;
  assign n9203 = n9200 | n9201;
  assign n9204 = ~n9202 & n9203;
  assign n14068 = n9001 | n9003;
  assign n14084 = n9204 & n14068;
  assign n14085 = n9001 & n9204;
  assign n14086 = (n13974 & n14084) | (n13974 & n14085) | (n14084 & n14085);
  assign n14087 = n9204 | n14068;
  assign n14088 = n9001 | n9204;
  assign n14089 = (n13974 & n14087) | (n13974 & n14088) | (n14087 & n14088);
  assign n9207 = ~n14086 & n14089;
  assign n9208 = x76 & x90;
  assign n9209 = n9207 & n9208;
  assign n9210 = n9207 | n9208;
  assign n9211 = ~n9209 & n9210;
  assign n14090 = n9008 & n9211;
  assign n16922 = (n9211 & n13998) | (n9211 & n14090) | (n13998 & n14090);
  assign n16923 = (n9211 & n13999) | (n9211 & n14090) | (n13999 & n14090);
  assign n16924 = (n13883 & n16922) | (n13883 & n16923) | (n16922 & n16923);
  assign n14092 = n9008 | n9211;
  assign n16925 = n13998 | n14092;
  assign n16926 = n13999 | n14092;
  assign n16927 = (n13883 & n16925) | (n13883 & n16926) | (n16925 & n16926);
  assign n9214 = ~n16924 & n16927;
  assign n9215 = x75 & x91;
  assign n9216 = n9214 & n9215;
  assign n9217 = n9214 | n9215;
  assign n9218 = ~n9216 & n9217;
  assign n9219 = n16910 & n9218;
  assign n9220 = n16910 | n9218;
  assign n9221 = ~n9219 & n9220;
  assign n9222 = x74 & x92;
  assign n9223 = n9221 & n9222;
  assign n9224 = n9221 | n9222;
  assign n9225 = ~n9223 & n9224;
  assign n14063 = n9022 | n9024;
  assign n14094 = n9225 & n14063;
  assign n14095 = n9022 & n9225;
  assign n14096 = (n16848 & n14094) | (n16848 & n14095) | (n14094 & n14095);
  assign n14097 = n9225 | n14063;
  assign n14098 = n9022 | n9225;
  assign n14099 = (n16848 & n14097) | (n16848 & n14098) | (n14097 & n14098);
  assign n9228 = ~n14096 & n14099;
  assign n9229 = x73 & x93;
  assign n9230 = n9228 & n9229;
  assign n9231 = n9228 | n9229;
  assign n9232 = ~n9230 & n9231;
  assign n14100 = n9029 & n9232;
  assign n16928 = (n9232 & n14009) | (n9232 & n14100) | (n14009 & n14100);
  assign n16929 = (n9232 & n14008) | (n9232 & n14100) | (n14008 & n14100);
  assign n16930 = (n13878 & n16928) | (n13878 & n16929) | (n16928 & n16929);
  assign n14102 = n9029 | n9232;
  assign n16931 = n14009 | n14102;
  assign n16932 = n14008 | n14102;
  assign n16933 = (n13878 & n16931) | (n13878 & n16932) | (n16931 & n16932);
  assign n9235 = ~n16930 & n16933;
  assign n9236 = x72 & x94;
  assign n9237 = n9235 & n9236;
  assign n9238 = n9235 | n9236;
  assign n9239 = ~n9237 & n9238;
  assign n14061 = n9036 | n9038;
  assign n16934 = n9239 & n14061;
  assign n16904 = n8827 | n9036;
  assign n16905 = (n9036 & n9038) | (n9036 & n16904) | (n9038 & n16904);
  assign n16935 = n9239 & n16905;
  assign n16936 = (n16828 & n16934) | (n16828 & n16935) | (n16934 & n16935);
  assign n16937 = n9239 | n14061;
  assign n16938 = n9239 | n16905;
  assign n16939 = (n16828 & n16937) | (n16828 & n16938) | (n16937 & n16938);
  assign n9242 = ~n16936 & n16939;
  assign n9243 = x71 & x95;
  assign n9244 = n9242 & n9243;
  assign n9245 = n9242 | n9243;
  assign n9246 = ~n9244 & n9245;
  assign n14104 = n9043 & n9246;
  assign n16940 = (n9246 & n14018) | (n9246 & n14104) | (n14018 & n14104);
  assign n16941 = (n9045 & n9246) | (n9045 & n14104) | (n9246 & n14104);
  assign n16942 = (n13928 & n16940) | (n13928 & n16941) | (n16940 & n16941);
  assign n14106 = n9043 | n9246;
  assign n16943 = n14018 | n14106;
  assign n16944 = n9045 | n14106;
  assign n16945 = (n13928 & n16943) | (n13928 & n16944) | (n16943 & n16944);
  assign n9249 = ~n16942 & n16945;
  assign n9250 = x70 & x96;
  assign n9251 = n9249 & n9250;
  assign n9252 = n9249 | n9250;
  assign n9253 = ~n9251 & n9252;
  assign n14108 = n9050 & n9253;
  assign n14109 = (n9253 & n14023) | (n9253 & n14108) | (n14023 & n14108);
  assign n14110 = n9050 | n9253;
  assign n14111 = n14023 | n14110;
  assign n9256 = ~n14109 & n14111;
  assign n9257 = x69 & x97;
  assign n9258 = n9256 & n9257;
  assign n9259 = n9256 | n9257;
  assign n9260 = ~n9258 & n9259;
  assign n14112 = n9057 & n9260;
  assign n14113 = (n9260 & n14027) | (n9260 & n14112) | (n14027 & n14112);
  assign n14114 = n9057 | n9260;
  assign n14115 = n14027 | n14114;
  assign n9263 = ~n14113 & n14115;
  assign n9264 = x68 & x98;
  assign n9265 = n9263 & n9264;
  assign n9266 = n9263 | n9264;
  assign n9267 = ~n9265 & n9266;
  assign n14116 = n9064 & n9267;
  assign n14117 = (n9267 & n14031) | (n9267 & n14116) | (n14031 & n14116);
  assign n14118 = n9064 | n9267;
  assign n14119 = n14031 | n14118;
  assign n9270 = ~n14117 & n14119;
  assign n9271 = x67 & x99;
  assign n9272 = n9270 & n9271;
  assign n9273 = n9270 | n9271;
  assign n9274 = ~n9272 & n9273;
  assign n14120 = n9071 & n9274;
  assign n14121 = (n9274 & n14035) | (n9274 & n14120) | (n14035 & n14120);
  assign n14122 = n9071 | n9274;
  assign n14123 = n14035 | n14122;
  assign n9277 = ~n14121 & n14123;
  assign n9278 = x66 & x100;
  assign n9279 = n9277 & n9278;
  assign n9280 = n9277 | n9278;
  assign n9281 = ~n9279 & n9280;
  assign n14124 = n9078 & n9281;
  assign n14125 = (n9281 & n14040) | (n9281 & n14124) | (n14040 & n14124);
  assign n14126 = n9078 | n9281;
  assign n14127 = n14040 | n14126;
  assign n9284 = ~n14125 & n14127;
  assign n9285 = x65 & x101;
  assign n9286 = n9284 & n9285;
  assign n9287 = n9284 | n9285;
  assign n9288 = ~n9286 & n9287;
  assign n14058 = n9085 | n9087;
  assign n14128 = n9288 & n14058;
  assign n14129 = n9085 & n9288;
  assign n14130 = (n13962 & n14128) | (n13962 & n14129) | (n14128 & n14129);
  assign n14131 = n9288 | n14058;
  assign n14132 = n9085 | n9288;
  assign n14133 = (n13962 & n14131) | (n13962 & n14132) | (n14131 & n14132);
  assign n9291 = ~n14130 & n14133;
  assign n9292 = x64 & x102;
  assign n9293 = n9291 & n9292;
  assign n9294 = n9291 | n9292;
  assign n9295 = ~n9293 & n9294;
  assign n14056 = n9092 | n9094;
  assign n16946 = n9295 & n14056;
  assign n16947 = n9092 & n9295;
  assign n16948 = (n13960 & n16946) | (n13960 & n16947) | (n16946 & n16947);
  assign n16949 = n9295 | n14056;
  assign n16950 = n9092 | n9295;
  assign n16951 = (n13960 & n16949) | (n13960 & n16950) | (n16949 & n16950);
  assign n9298 = ~n16948 & n16951;
  assign n9299 = x63 & x103;
  assign n9300 = n9298 & n9299;
  assign n9301 = n9298 | n9299;
  assign n9302 = ~n9300 & n9301;
  assign n14054 = n9099 | n9101;
  assign n16952 = n9302 & n14054;
  assign n16953 = n9099 & n9302;
  assign n16954 = (n13958 & n16952) | (n13958 & n16953) | (n16952 & n16953);
  assign n16955 = n9302 | n14054;
  assign n16956 = n9099 | n9302;
  assign n16957 = (n13958 & n16955) | (n13958 & n16956) | (n16955 & n16956);
  assign n9305 = ~n16954 & n16957;
  assign n9306 = x62 & x104;
  assign n9307 = n9305 & n9306;
  assign n9308 = n9305 | n9306;
  assign n9309 = ~n9307 & n9308;
  assign n9310 = n14053 & n9309;
  assign n9311 = n14053 | n9309;
  assign n9312 = ~n9310 & n9311;
  assign n9313 = x61 & x105;
  assign n9314 = n9312 & n9313;
  assign n9315 = n9312 | n9313;
  assign n9316 = ~n9314 & n9315;
  assign n9317 = n14051 & n9316;
  assign n9318 = n14051 | n9316;
  assign n9319 = ~n9317 & n9318;
  assign n9320 = x60 & x106;
  assign n9321 = n9319 & n9320;
  assign n9322 = n9319 | n9320;
  assign n9323 = ~n9321 & n9322;
  assign n9324 = n14049 & n9323;
  assign n9325 = n14049 | n9323;
  assign n9326 = ~n9324 & n9325;
  assign n9327 = x59 & x107;
  assign n9328 = n9326 & n9327;
  assign n9329 = n9326 | n9327;
  assign n9330 = ~n9328 & n9329;
  assign n9331 = n14047 & n9330;
  assign n9332 = n14047 | n9330;
  assign n9333 = ~n9331 & n9332;
  assign n9334 = x58 & x108;
  assign n9335 = n9333 & n9334;
  assign n9336 = n9333 | n9334;
  assign n9337 = ~n9335 & n9336;
  assign n9338 = n14045 & n9337;
  assign n9339 = n14045 | n9337;
  assign n9340 = ~n9338 & n9339;
  assign n9341 = x57 & x109;
  assign n9342 = n9340 & n9341;
  assign n9343 = n9340 | n9341;
  assign n9344 = ~n9342 & n9343;
  assign n9345 = n9163 & n9344;
  assign n9346 = n9163 | n9344;
  assign n9347 = ~n9345 & n9346;
  assign n9348 = x56 & x110;
  assign n9349 = n9347 & n9348;
  assign n9350 = n9347 | n9348;
  assign n9351 = ~n9349 & n9350;
  assign n9352 = n9162 & n9351;
  assign n9353 = n9162 | n9351;
  assign n9354 = ~n9352 & n9353;
  assign n9355 = x55 & x111;
  assign n9356 = n9354 & n9355;
  assign n9357 = n9354 | n9355;
  assign n9358 = ~n9356 & n9357;
  assign n9359 = n9161 & n9358;
  assign n9360 = n9161 | n9358;
  assign n9361 = ~n9359 & n9360;
  assign n9362 = n9356 | n9359;
  assign n9363 = n9349 | n9352;
  assign n14134 = n9342 | n9344;
  assign n14135 = (n9163 & n9342) | (n9163 & n14134) | (n9342 & n14134);
  assign n14136 = n9335 | n9337;
  assign n14137 = (n9335 & n14045) | (n9335 & n14136) | (n14045 & n14136);
  assign n14138 = n9328 | n9330;
  assign n14139 = (n9328 & n14047) | (n9328 & n14138) | (n14047 & n14138);
  assign n14140 = n9321 | n9323;
  assign n14141 = (n9321 & n14049) | (n9321 & n14140) | (n14049 & n14140);
  assign n14142 = n9314 | n9316;
  assign n14143 = (n9314 & n14051) | (n9314 & n14142) | (n14051 & n14142);
  assign n14055 = (n9099 & n13958) | (n9099 & n14054) | (n13958 & n14054);
  assign n14057 = (n9092 & n13960) | (n9092 & n14056) | (n13960 & n14056);
  assign n14062 = (n16828 & n16905) | (n16828 & n14061) | (n16905 & n14061);
  assign n14153 = n9230 | n9232;
  assign n16958 = n9029 | n9230;
  assign n16959 = (n9230 & n9232) | (n9230 & n16958) | (n9232 & n16958);
  assign n16960 = (n14009 & n14153) | (n14009 & n16959) | (n14153 & n16959);
  assign n16961 = (n14008 & n14153) | (n14008 & n16959) | (n14153 & n16959);
  assign n16962 = (n13878 & n16960) | (n13878 & n16961) | (n16960 & n16961);
  assign n14158 = n9209 | n9211;
  assign n16963 = n9008 | n9209;
  assign n16964 = (n9209 & n9211) | (n9209 & n16963) | (n9211 & n16963);
  assign n16965 = (n13998 & n14158) | (n13998 & n16964) | (n14158 & n16964);
  assign n16966 = (n13999 & n14158) | (n13999 & n16964) | (n14158 & n16964);
  assign n16967 = (n13883 & n16965) | (n13883 & n16966) | (n16965 & n16966);
  assign n9387 = x79 & x88;
  assign n16969 = n9387 & n16919;
  assign n50007 = n9187 & n9387;
  assign n50008 = n16865 & n50007;
  assign n16971 = (n16857 & n16969) | (n16857 & n50008) | (n16969 & n50008);
  assign n16968 = (n9190 & n9387) | (n9190 & n16971) | (n9387 & n16971);
  assign n14166 = (n14075 & n16968) | (n14075 & n16971) | (n16968 & n16971);
  assign n16973 = n9387 | n16919;
  assign n50009 = n9187 | n9387;
  assign n50010 = (n9387 & n16865) | (n9387 & n50009) | (n16865 & n50009);
  assign n16975 = (n16857 & n16973) | (n16857 & n50010) | (n16973 & n50010);
  assign n16972 = n9190 | n16975;
  assign n14169 = (n14075 & n16972) | (n14075 & n16975) | (n16972 & n16975);
  assign n9390 = ~n14166 & n14169;
  assign n14171 = n9195 & n9390;
  assign n16976 = (n9197 & n9390) | (n9197 & n14171) | (n9390 & n14171);
  assign n14172 = (n16915 & n16976) | (n16915 & n14171) | (n16976 & n14171);
  assign n14174 = n9195 | n9390;
  assign n16977 = n9197 | n14174;
  assign n14175 = (n16915 & n16977) | (n16915 & n14174) | (n16977 & n14174);
  assign n9393 = ~n14172 & n14175;
  assign n9394 = x78 & x89;
  assign n9395 = n9393 & n9394;
  assign n9396 = n9393 | n9394;
  assign n9397 = ~n9395 & n9396;
  assign n14176 = n9202 & n9397;
  assign n16978 = (n9397 & n14085) | (n9397 & n14176) | (n14085 & n14176);
  assign n16979 = (n9397 & n14084) | (n9397 & n14176) | (n14084 & n14176);
  assign n16980 = (n13974 & n16978) | (n13974 & n16979) | (n16978 & n16979);
  assign n14178 = n9202 | n9397;
  assign n16981 = n14085 | n14178;
  assign n16982 = n14084 | n14178;
  assign n16983 = (n13974 & n16981) | (n13974 & n16982) | (n16981 & n16982);
  assign n9400 = ~n16980 & n16983;
  assign n9401 = x77 & x90;
  assign n9402 = n9400 & n9401;
  assign n9403 = n9400 | n9401;
  assign n9404 = ~n9402 & n9403;
  assign n9405 = n16967 & n9404;
  assign n9406 = n16967 | n9404;
  assign n9407 = ~n9405 & n9406;
  assign n9408 = x76 & x91;
  assign n9409 = n9407 & n9408;
  assign n9410 = n9407 | n9408;
  assign n9411 = ~n9409 & n9410;
  assign n14155 = n9216 | n9218;
  assign n14180 = n9411 & n14155;
  assign n14181 = n9216 & n9411;
  assign n14182 = (n16910 & n14180) | (n16910 & n14181) | (n14180 & n14181);
  assign n14183 = n9411 | n14155;
  assign n14184 = n9216 | n9411;
  assign n14185 = (n16910 & n14183) | (n16910 & n14184) | (n14183 & n14184);
  assign n9414 = ~n14182 & n14185;
  assign n9415 = x75 & x92;
  assign n9416 = n9414 & n9415;
  assign n9417 = n9414 | n9415;
  assign n9418 = ~n9416 & n9417;
  assign n14186 = n9223 & n9418;
  assign n16984 = (n9418 & n14095) | (n9418 & n14186) | (n14095 & n14186);
  assign n16985 = (n9418 & n14094) | (n9418 & n14186) | (n14094 & n14186);
  assign n16986 = (n16848 & n16984) | (n16848 & n16985) | (n16984 & n16985);
  assign n14188 = n9223 | n9418;
  assign n16987 = n14095 | n14188;
  assign n16988 = n14094 | n14188;
  assign n16989 = (n16848 & n16987) | (n16848 & n16988) | (n16987 & n16988);
  assign n9421 = ~n16986 & n16989;
  assign n9422 = x74 & x93;
  assign n9423 = n9421 & n9422;
  assign n9424 = n9421 | n9422;
  assign n9425 = ~n9423 & n9424;
  assign n9426 = n16962 & n9425;
  assign n9427 = n16962 | n9425;
  assign n9428 = ~n9426 & n9427;
  assign n9429 = x73 & x94;
  assign n9430 = n9428 & n9429;
  assign n9431 = n9428 | n9429;
  assign n9432 = ~n9430 & n9431;
  assign n14150 = n9237 | n9239;
  assign n14190 = n9432 & n14150;
  assign n14191 = n9237 & n9432;
  assign n14192 = (n14062 & n14190) | (n14062 & n14191) | (n14190 & n14191);
  assign n14193 = n9432 | n14150;
  assign n14194 = n9237 | n9432;
  assign n14195 = (n14062 & n14193) | (n14062 & n14194) | (n14193 & n14194);
  assign n9435 = ~n14192 & n14195;
  assign n9436 = x72 & x95;
  assign n9437 = n9435 & n9436;
  assign n9438 = n9435 | n9436;
  assign n9439 = ~n9437 & n9438;
  assign n14196 = n9244 & n9439;
  assign n14197 = (n9439 & n16942) | (n9439 & n14196) | (n16942 & n14196);
  assign n14198 = n9244 | n9439;
  assign n14199 = n16942 | n14198;
  assign n9442 = ~n14197 & n14199;
  assign n9443 = x71 & x96;
  assign n9444 = n9442 & n9443;
  assign n9445 = n9442 | n9443;
  assign n9446 = ~n9444 & n9445;
  assign n14200 = n9251 & n9446;
  assign n14201 = (n9446 & n14109) | (n9446 & n14200) | (n14109 & n14200);
  assign n14202 = n9251 | n9446;
  assign n14203 = n14109 | n14202;
  assign n9449 = ~n14201 & n14203;
  assign n9450 = x70 & x97;
  assign n9451 = n9449 & n9450;
  assign n9452 = n9449 | n9450;
  assign n9453 = ~n9451 & n9452;
  assign n14204 = n9258 & n9453;
  assign n14205 = (n9453 & n14113) | (n9453 & n14204) | (n14113 & n14204);
  assign n14206 = n9258 | n9453;
  assign n14207 = n14113 | n14206;
  assign n9456 = ~n14205 & n14207;
  assign n9457 = x69 & x98;
  assign n9458 = n9456 & n9457;
  assign n9459 = n9456 | n9457;
  assign n9460 = ~n9458 & n9459;
  assign n14208 = n9265 & n9460;
  assign n14209 = (n9460 & n14117) | (n9460 & n14208) | (n14117 & n14208);
  assign n14210 = n9265 | n9460;
  assign n14211 = n14117 | n14210;
  assign n9463 = ~n14209 & n14211;
  assign n9464 = x68 & x99;
  assign n9465 = n9463 & n9464;
  assign n9466 = n9463 | n9464;
  assign n9467 = ~n9465 & n9466;
  assign n14212 = n9272 & n9467;
  assign n14213 = (n9467 & n14121) | (n9467 & n14212) | (n14121 & n14212);
  assign n14214 = n9272 | n9467;
  assign n14215 = n14121 | n14214;
  assign n9470 = ~n14213 & n14215;
  assign n9471 = x67 & x100;
  assign n9472 = n9470 & n9471;
  assign n9473 = n9470 | n9471;
  assign n9474 = ~n9472 & n9473;
  assign n14216 = n9279 & n9474;
  assign n14217 = (n9474 & n14125) | (n9474 & n14216) | (n14125 & n14216);
  assign n14218 = n9279 | n9474;
  assign n14219 = n14125 | n14218;
  assign n9477 = ~n14217 & n14219;
  assign n9478 = x66 & x101;
  assign n9479 = n9477 & n9478;
  assign n9480 = n9477 | n9478;
  assign n9481 = ~n9479 & n9480;
  assign n14220 = n9286 & n9481;
  assign n14221 = (n9481 & n14130) | (n9481 & n14220) | (n14130 & n14220);
  assign n14222 = n9286 | n9481;
  assign n14223 = n14130 | n14222;
  assign n9484 = ~n14221 & n14223;
  assign n9485 = x65 & x102;
  assign n9486 = n9484 & n9485;
  assign n9487 = n9484 | n9485;
  assign n9488 = ~n9486 & n9487;
  assign n14148 = n9293 | n9295;
  assign n14224 = n9488 & n14148;
  assign n14225 = n9293 & n9488;
  assign n14226 = (n14057 & n14224) | (n14057 & n14225) | (n14224 & n14225);
  assign n14227 = n9488 | n14148;
  assign n14228 = n9293 | n9488;
  assign n14229 = (n14057 & n14227) | (n14057 & n14228) | (n14227 & n14228);
  assign n9491 = ~n14226 & n14229;
  assign n9492 = x64 & x103;
  assign n9493 = n9491 & n9492;
  assign n9494 = n9491 | n9492;
  assign n9495 = ~n9493 & n9494;
  assign n14146 = n9300 | n9302;
  assign n16990 = n9495 & n14146;
  assign n16991 = n9300 & n9495;
  assign n16992 = (n14055 & n16990) | (n14055 & n16991) | (n16990 & n16991);
  assign n16993 = n9495 | n14146;
  assign n16994 = n9300 | n9495;
  assign n16995 = (n14055 & n16993) | (n14055 & n16994) | (n16993 & n16994);
  assign n9498 = ~n16992 & n16995;
  assign n9499 = x63 & x104;
  assign n9500 = n9498 & n9499;
  assign n9501 = n9498 | n9499;
  assign n9502 = ~n9500 & n9501;
  assign n14144 = n9307 | n9309;
  assign n16996 = n9502 & n14144;
  assign n16997 = n9307 & n9502;
  assign n16998 = (n14053 & n16996) | (n14053 & n16997) | (n16996 & n16997);
  assign n16999 = n9502 | n14144;
  assign n17000 = n9307 | n9502;
  assign n17001 = (n14053 & n16999) | (n14053 & n17000) | (n16999 & n17000);
  assign n9505 = ~n16998 & n17001;
  assign n9506 = x62 & x105;
  assign n9507 = n9505 & n9506;
  assign n9508 = n9505 | n9506;
  assign n9509 = ~n9507 & n9508;
  assign n9510 = n14143 & n9509;
  assign n9511 = n14143 | n9509;
  assign n9512 = ~n9510 & n9511;
  assign n9513 = x61 & x106;
  assign n9514 = n9512 & n9513;
  assign n9515 = n9512 | n9513;
  assign n9516 = ~n9514 & n9515;
  assign n9517 = n14141 & n9516;
  assign n9518 = n14141 | n9516;
  assign n9519 = ~n9517 & n9518;
  assign n9520 = x60 & x107;
  assign n9521 = n9519 & n9520;
  assign n9522 = n9519 | n9520;
  assign n9523 = ~n9521 & n9522;
  assign n9524 = n14139 & n9523;
  assign n9525 = n14139 | n9523;
  assign n9526 = ~n9524 & n9525;
  assign n9527 = x59 & x108;
  assign n9528 = n9526 & n9527;
  assign n9529 = n9526 | n9527;
  assign n9530 = ~n9528 & n9529;
  assign n9531 = n14137 & n9530;
  assign n9532 = n14137 | n9530;
  assign n9533 = ~n9531 & n9532;
  assign n9534 = x58 & x109;
  assign n9535 = n9533 & n9534;
  assign n9536 = n9533 | n9534;
  assign n9537 = ~n9535 & n9536;
  assign n9538 = n14135 & n9537;
  assign n9539 = n14135 | n9537;
  assign n9540 = ~n9538 & n9539;
  assign n9541 = x57 & x110;
  assign n9542 = n9540 & n9541;
  assign n9543 = n9540 | n9541;
  assign n9544 = ~n9542 & n9543;
  assign n9545 = n9363 & n9544;
  assign n9546 = n9363 | n9544;
  assign n9547 = ~n9545 & n9546;
  assign n9548 = x56 & x111;
  assign n9549 = n9547 & n9548;
  assign n9550 = n9547 | n9548;
  assign n9551 = ~n9549 & n9550;
  assign n9552 = n9362 & n9551;
  assign n9553 = n9362 | n9551;
  assign n9554 = ~n9552 & n9553;
  assign n9555 = n9549 | n9552;
  assign n14230 = n9542 | n9544;
  assign n14231 = (n9363 & n9542) | (n9363 & n14230) | (n9542 & n14230);
  assign n14232 = n9535 | n9537;
  assign n14233 = (n9535 & n14135) | (n9535 & n14232) | (n14135 & n14232);
  assign n14234 = n9528 | n9530;
  assign n14235 = (n9528 & n14137) | (n9528 & n14234) | (n14137 & n14234);
  assign n14236 = n9521 | n9523;
  assign n14237 = (n9521 & n14139) | (n9521 & n14236) | (n14139 & n14236);
  assign n14238 = n9514 | n9516;
  assign n14239 = (n9514 & n14141) | (n9514 & n14238) | (n14141 & n14238);
  assign n14145 = (n9307 & n14053) | (n9307 & n14144) | (n14053 & n14144);
  assign n14147 = (n9300 & n14055) | (n9300 & n14146) | (n14055 & n14146);
  assign n14252 = n9416 | n9418;
  assign n17004 = n9223 | n9416;
  assign n17005 = (n9416 & n9418) | (n9416 & n17004) | (n9418 & n17004);
  assign n17006 = (n14095 & n14252) | (n14095 & n17005) | (n14252 & n17005);
  assign n17007 = (n14094 & n14252) | (n14094 & n17005) | (n14252 & n17005);
  assign n17008 = (n16848 & n17006) | (n16848 & n17007) | (n17006 & n17007);
  assign n14257 = n9395 | n9397;
  assign n17009 = n9202 | n9395;
  assign n17010 = (n9395 & n9397) | (n9395 & n17009) | (n9397 & n17009);
  assign n17011 = (n14085 & n14257) | (n14085 & n17010) | (n14257 & n17010);
  assign n17012 = (n14084 & n14257) | (n14084 & n17010) | (n14257 & n17010);
  assign n17013 = (n13974 & n17011) | (n13974 & n17012) | (n17011 & n17012);
  assign n9579 = x79 & x89;
  assign n50011 = n9387 & n9579;
  assign n66401 = n16919 & n50011;
  assign n66402 = n9579 & n50007;
  assign n66403 = n16865 & n66402;
  assign n50015 = (n16857 & n66401) | (n16857 & n66403) | (n66401 & n66403);
  assign n50012 = (n9190 & n50015) | (n9190 & n50011) | (n50015 & n50011);
  assign n17016 = (n14075 & n50012) | (n14075 & n50015) | (n50012 & n50015);
  assign n17017 = (n9579 & n16976) | (n9579 & n17016) | (n16976 & n17016);
  assign n50016 = (n9390 & n9579) | (n9390 & n17016) | (n9579 & n17016);
  assign n66404 = n9579 & n50012;
  assign n66405 = n9579 & n50015;
  assign n66406 = (n14075 & n66404) | (n14075 & n66405) | (n66404 & n66405);
  assign n50018 = (n9195 & n50016) | (n9195 & n66406) | (n50016 & n66406);
  assign n17019 = (n16915 & n17017) | (n16915 & n50018) | (n17017 & n50018);
  assign n50019 = n9387 | n9579;
  assign n66407 = (n9579 & n16919) | (n9579 & n50019) | (n16919 & n50019);
  assign n66408 = n9579 | n50007;
  assign n66409 = (n9579 & n16865) | (n9579 & n66408) | (n16865 & n66408);
  assign n50023 = (n16857 & n66407) | (n16857 & n66409) | (n66407 & n66409);
  assign n50020 = (n9190 & n50023) | (n9190 & n50019) | (n50023 & n50019);
  assign n17022 = (n14075 & n50020) | (n14075 & n50023) | (n50020 & n50023);
  assign n17023 = n16976 | n17022;
  assign n50024 = n9390 | n17022;
  assign n50025 = (n9195 & n17022) | (n9195 & n50024) | (n17022 & n50024);
  assign n17025 = (n16915 & n17023) | (n16915 & n50025) | (n17023 & n50025);
  assign n9582 = ~n17019 & n17025;
  assign n9583 = n17013 & n9582;
  assign n9584 = n17013 | n9582;
  assign n9585 = ~n9583 & n9584;
  assign n9586 = x78 & x90;
  assign n9587 = n9585 & n9586;
  assign n9588 = n9585 | n9586;
  assign n9589 = ~n9587 & n9588;
  assign n14254 = n9402 | n9404;
  assign n14263 = n9589 & n14254;
  assign n14264 = n9402 & n9589;
  assign n14265 = (n16967 & n14263) | (n16967 & n14264) | (n14263 & n14264);
  assign n14266 = n9589 | n14254;
  assign n14267 = n9402 | n9589;
  assign n14268 = (n16967 & n14266) | (n16967 & n14267) | (n14266 & n14267);
  assign n9592 = ~n14265 & n14268;
  assign n9593 = x77 & x91;
  assign n9594 = n9592 & n9593;
  assign n9595 = n9592 | n9593;
  assign n9596 = ~n9594 & n9595;
  assign n14269 = n9409 & n9596;
  assign n17026 = (n9596 & n14181) | (n9596 & n14269) | (n14181 & n14269);
  assign n17027 = (n9596 & n14180) | (n9596 & n14269) | (n14180 & n14269);
  assign n17028 = (n16910 & n17026) | (n16910 & n17027) | (n17026 & n17027);
  assign n14271 = n9409 | n9596;
  assign n17029 = n14181 | n14271;
  assign n17030 = n14180 | n14271;
  assign n17031 = (n16910 & n17029) | (n16910 & n17030) | (n17029 & n17030);
  assign n9599 = ~n17028 & n17031;
  assign n9600 = x76 & x92;
  assign n9601 = n9599 & n9600;
  assign n9602 = n9599 | n9600;
  assign n9603 = ~n9601 & n9602;
  assign n9604 = n17008 & n9603;
  assign n9605 = n17008 | n9603;
  assign n9606 = ~n9604 & n9605;
  assign n9607 = x75 & x93;
  assign n9608 = n9606 & n9607;
  assign n9609 = n9606 | n9607;
  assign n9610 = ~n9608 & n9609;
  assign n14249 = n9423 | n9425;
  assign n14273 = n9610 & n14249;
  assign n14274 = n9423 & n9610;
  assign n14275 = (n16962 & n14273) | (n16962 & n14274) | (n14273 & n14274);
  assign n14276 = n9610 | n14249;
  assign n14277 = n9423 | n9610;
  assign n14278 = (n16962 & n14276) | (n16962 & n14277) | (n14276 & n14277);
  assign n9613 = ~n14275 & n14278;
  assign n9614 = x74 & x94;
  assign n9615 = n9613 & n9614;
  assign n9616 = n9613 | n9614;
  assign n9617 = ~n9615 & n9616;
  assign n14279 = n9430 & n9617;
  assign n17032 = (n9617 & n14191) | (n9617 & n14279) | (n14191 & n14279);
  assign n17033 = (n9617 & n14190) | (n9617 & n14279) | (n14190 & n14279);
  assign n17034 = (n14062 & n17032) | (n14062 & n17033) | (n17032 & n17033);
  assign n14281 = n9430 | n9617;
  assign n17035 = n14191 | n14281;
  assign n17036 = n14190 | n14281;
  assign n17037 = (n14062 & n17035) | (n14062 & n17036) | (n17035 & n17036);
  assign n9620 = ~n17034 & n17037;
  assign n9621 = x73 & x95;
  assign n9622 = n9620 & n9621;
  assign n9623 = n9620 | n9621;
  assign n9624 = ~n9622 & n9623;
  assign n14247 = n9437 | n9439;
  assign n17038 = n9624 & n14247;
  assign n17002 = n9244 | n9437;
  assign n17003 = (n9437 & n9439) | (n9437 & n17002) | (n9439 & n17002);
  assign n17039 = n9624 & n17003;
  assign n17040 = (n16942 & n17038) | (n16942 & n17039) | (n17038 & n17039);
  assign n17041 = n9624 | n14247;
  assign n17042 = n9624 | n17003;
  assign n17043 = (n16942 & n17041) | (n16942 & n17042) | (n17041 & n17042);
  assign n9627 = ~n17040 & n17043;
  assign n9628 = x72 & x96;
  assign n9629 = n9627 & n9628;
  assign n9630 = n9627 | n9628;
  assign n9631 = ~n9629 & n9630;
  assign n14283 = n9444 & n9631;
  assign n17044 = (n9631 & n14200) | (n9631 & n14283) | (n14200 & n14283);
  assign n17045 = (n9446 & n9631) | (n9446 & n14283) | (n9631 & n14283);
  assign n17046 = (n14109 & n17044) | (n14109 & n17045) | (n17044 & n17045);
  assign n14285 = n9444 | n9631;
  assign n17047 = n14200 | n14285;
  assign n17048 = n9446 | n14285;
  assign n17049 = (n14109 & n17047) | (n14109 & n17048) | (n17047 & n17048);
  assign n9634 = ~n17046 & n17049;
  assign n9635 = x71 & x97;
  assign n9636 = n9634 & n9635;
  assign n9637 = n9634 | n9635;
  assign n9638 = ~n9636 & n9637;
  assign n14287 = n9451 & n9638;
  assign n14288 = (n9638 & n14205) | (n9638 & n14287) | (n14205 & n14287);
  assign n14289 = n9451 | n9638;
  assign n14290 = n14205 | n14289;
  assign n9641 = ~n14288 & n14290;
  assign n9642 = x70 & x98;
  assign n9643 = n9641 & n9642;
  assign n9644 = n9641 | n9642;
  assign n9645 = ~n9643 & n9644;
  assign n14291 = n9458 & n9645;
  assign n14292 = (n9645 & n14209) | (n9645 & n14291) | (n14209 & n14291);
  assign n14293 = n9458 | n9645;
  assign n14294 = n14209 | n14293;
  assign n9648 = ~n14292 & n14294;
  assign n9649 = x69 & x99;
  assign n9650 = n9648 & n9649;
  assign n9651 = n9648 | n9649;
  assign n9652 = ~n9650 & n9651;
  assign n14295 = n9465 & n9652;
  assign n14296 = (n9652 & n14213) | (n9652 & n14295) | (n14213 & n14295);
  assign n14297 = n9465 | n9652;
  assign n14298 = n14213 | n14297;
  assign n9655 = ~n14296 & n14298;
  assign n9656 = x68 & x100;
  assign n9657 = n9655 & n9656;
  assign n9658 = n9655 | n9656;
  assign n9659 = ~n9657 & n9658;
  assign n14299 = n9472 & n9659;
  assign n14300 = (n9659 & n14217) | (n9659 & n14299) | (n14217 & n14299);
  assign n14301 = n9472 | n9659;
  assign n14302 = n14217 | n14301;
  assign n9662 = ~n14300 & n14302;
  assign n9663 = x67 & x101;
  assign n9664 = n9662 & n9663;
  assign n9665 = n9662 | n9663;
  assign n9666 = ~n9664 & n9665;
  assign n14303 = n9479 & n9666;
  assign n14304 = (n9666 & n14221) | (n9666 & n14303) | (n14221 & n14303);
  assign n14305 = n9479 | n9666;
  assign n14306 = n14221 | n14305;
  assign n9669 = ~n14304 & n14306;
  assign n9670 = x66 & x102;
  assign n9671 = n9669 & n9670;
  assign n9672 = n9669 | n9670;
  assign n9673 = ~n9671 & n9672;
  assign n14307 = n9486 & n9673;
  assign n14308 = (n9673 & n14226) | (n9673 & n14307) | (n14226 & n14307);
  assign n14309 = n9486 | n9673;
  assign n14310 = n14226 | n14309;
  assign n9676 = ~n14308 & n14310;
  assign n9677 = x65 & x103;
  assign n9678 = n9676 & n9677;
  assign n9679 = n9676 | n9677;
  assign n9680 = ~n9678 & n9679;
  assign n14244 = n9493 | n9495;
  assign n14311 = n9680 & n14244;
  assign n14312 = n9493 & n9680;
  assign n14313 = (n14147 & n14311) | (n14147 & n14312) | (n14311 & n14312);
  assign n14314 = n9680 | n14244;
  assign n14315 = n9493 | n9680;
  assign n14316 = (n14147 & n14314) | (n14147 & n14315) | (n14314 & n14315);
  assign n9683 = ~n14313 & n14316;
  assign n9684 = x64 & x104;
  assign n9685 = n9683 & n9684;
  assign n9686 = n9683 | n9684;
  assign n9687 = ~n9685 & n9686;
  assign n14242 = n9500 | n9502;
  assign n17050 = n9687 & n14242;
  assign n17051 = n9500 & n9687;
  assign n17052 = (n14145 & n17050) | (n14145 & n17051) | (n17050 & n17051);
  assign n17053 = n9687 | n14242;
  assign n17054 = n9500 | n9687;
  assign n17055 = (n14145 & n17053) | (n14145 & n17054) | (n17053 & n17054);
  assign n9690 = ~n17052 & n17055;
  assign n9691 = x63 & x105;
  assign n9692 = n9690 & n9691;
  assign n9693 = n9690 | n9691;
  assign n9694 = ~n9692 & n9693;
  assign n14240 = n9507 | n9509;
  assign n17056 = n9694 & n14240;
  assign n17057 = n9507 & n9694;
  assign n17058 = (n14143 & n17056) | (n14143 & n17057) | (n17056 & n17057);
  assign n17059 = n9694 | n14240;
  assign n17060 = n9507 | n9694;
  assign n17061 = (n14143 & n17059) | (n14143 & n17060) | (n17059 & n17060);
  assign n9697 = ~n17058 & n17061;
  assign n9698 = x62 & x106;
  assign n9699 = n9697 & n9698;
  assign n9700 = n9697 | n9698;
  assign n9701 = ~n9699 & n9700;
  assign n9702 = n14239 & n9701;
  assign n9703 = n14239 | n9701;
  assign n9704 = ~n9702 & n9703;
  assign n9705 = x61 & x107;
  assign n9706 = n9704 & n9705;
  assign n9707 = n9704 | n9705;
  assign n9708 = ~n9706 & n9707;
  assign n9709 = n14237 & n9708;
  assign n9710 = n14237 | n9708;
  assign n9711 = ~n9709 & n9710;
  assign n9712 = x60 & x108;
  assign n9713 = n9711 & n9712;
  assign n9714 = n9711 | n9712;
  assign n9715 = ~n9713 & n9714;
  assign n9716 = n14235 & n9715;
  assign n9717 = n14235 | n9715;
  assign n9718 = ~n9716 & n9717;
  assign n9719 = x59 & x109;
  assign n9720 = n9718 & n9719;
  assign n9721 = n9718 | n9719;
  assign n9722 = ~n9720 & n9721;
  assign n9723 = n14233 & n9722;
  assign n9724 = n14233 | n9722;
  assign n9725 = ~n9723 & n9724;
  assign n9726 = x58 & x110;
  assign n9727 = n9725 & n9726;
  assign n9728 = n9725 | n9726;
  assign n9729 = ~n9727 & n9728;
  assign n9730 = n14231 & n9729;
  assign n9731 = n14231 | n9729;
  assign n9732 = ~n9730 & n9731;
  assign n9733 = x57 & x111;
  assign n9734 = n9732 & n9733;
  assign n9735 = n9732 | n9733;
  assign n9736 = ~n9734 & n9735;
  assign n9737 = n9555 & n9736;
  assign n9738 = n9555 | n9736;
  assign n9739 = ~n9737 & n9738;
  assign n14317 = n9734 | n9736;
  assign n14318 = (n9555 & n9734) | (n9555 & n14317) | (n9734 & n14317);
  assign n14319 = n9727 | n9729;
  assign n14320 = (n9727 & n14231) | (n9727 & n14319) | (n14231 & n14319);
  assign n14321 = n9720 | n9722;
  assign n14322 = (n9720 & n14233) | (n9720 & n14321) | (n14233 & n14321);
  assign n14323 = n9713 | n9715;
  assign n14324 = (n9713 & n14235) | (n9713 & n14323) | (n14235 & n14323);
  assign n14325 = n9706 | n9708;
  assign n14326 = (n9706 & n14237) | (n9706 & n14325) | (n14237 & n14325);
  assign n14241 = (n9507 & n14143) | (n9507 & n14240) | (n14143 & n14240);
  assign n14243 = (n9500 & n14145) | (n9500 & n14242) | (n14145 & n14242);
  assign n14248 = (n16942 & n17003) | (n16942 & n14247) | (n17003 & n14247);
  assign n14336 = n9615 | n9617;
  assign n17062 = n9430 | n9615;
  assign n17063 = (n9615 & n9617) | (n9615 & n17062) | (n9617 & n17062);
  assign n17064 = (n14191 & n14336) | (n14191 & n17063) | (n14336 & n17063);
  assign n17065 = (n14190 & n14336) | (n14190 & n17063) | (n14336 & n17063);
  assign n17066 = (n14062 & n17064) | (n14062 & n17065) | (n17064 & n17065);
  assign n14341 = n9594 | n9596;
  assign n17067 = n9409 | n9594;
  assign n17068 = (n9594 & n9596) | (n9594 & n17067) | (n9596 & n17067);
  assign n17069 = (n14181 & n14341) | (n14181 & n17068) | (n14341 & n17068);
  assign n17070 = (n14180 & n14341) | (n14180 & n17068) | (n14341 & n17068);
  assign n17071 = (n16910 & n17069) | (n16910 & n17070) | (n17069 & n17070);
  assign n9763 = x79 & x90;
  assign n17072 = n9763 & n17019;
  assign n17073 = (n9582 & n9763) | (n9582 & n17072) | (n9763 & n17072);
  assign n14346 = n9763 & n17019;
  assign n14347 = (n17013 & n17073) | (n17013 & n14346) | (n17073 & n14346);
  assign n17074 = n9763 | n17019;
  assign n17075 = n9582 | n17074;
  assign n14349 = n9763 | n17019;
  assign n14350 = (n17013 & n17075) | (n17013 & n14349) | (n17075 & n14349);
  assign n9766 = ~n14347 & n14350;
  assign n14351 = n9587 & n9766;
  assign n17076 = (n9766 & n14264) | (n9766 & n14351) | (n14264 & n14351);
  assign n17077 = (n9766 & n14263) | (n9766 & n14351) | (n14263 & n14351);
  assign n17078 = (n16967 & n17076) | (n16967 & n17077) | (n17076 & n17077);
  assign n14353 = n9587 | n9766;
  assign n17079 = n14264 | n14353;
  assign n17080 = n14263 | n14353;
  assign n17081 = (n16967 & n17079) | (n16967 & n17080) | (n17079 & n17080);
  assign n9769 = ~n17078 & n17081;
  assign n9770 = x78 & x91;
  assign n9771 = n9769 & n9770;
  assign n9772 = n9769 | n9770;
  assign n9773 = ~n9771 & n9772;
  assign n9774 = n17071 & n9773;
  assign n9775 = n17071 | n9773;
  assign n9776 = ~n9774 & n9775;
  assign n9777 = x77 & x92;
  assign n9778 = n9776 & n9777;
  assign n9779 = n9776 | n9777;
  assign n9780 = ~n9778 & n9779;
  assign n14338 = n9601 | n9603;
  assign n14355 = n9780 & n14338;
  assign n14356 = n9601 & n9780;
  assign n14357 = (n17008 & n14355) | (n17008 & n14356) | (n14355 & n14356);
  assign n14358 = n9780 | n14338;
  assign n14359 = n9601 | n9780;
  assign n14360 = (n17008 & n14358) | (n17008 & n14359) | (n14358 & n14359);
  assign n9783 = ~n14357 & n14360;
  assign n9784 = x76 & x93;
  assign n9785 = n9783 & n9784;
  assign n9786 = n9783 | n9784;
  assign n9787 = ~n9785 & n9786;
  assign n14361 = n9608 & n9787;
  assign n17082 = (n9787 & n14274) | (n9787 & n14361) | (n14274 & n14361);
  assign n17083 = (n9787 & n14273) | (n9787 & n14361) | (n14273 & n14361);
  assign n17084 = (n16962 & n17082) | (n16962 & n17083) | (n17082 & n17083);
  assign n14363 = n9608 | n9787;
  assign n17085 = n14274 | n14363;
  assign n17086 = n14273 | n14363;
  assign n17087 = (n16962 & n17085) | (n16962 & n17086) | (n17085 & n17086);
  assign n9790 = ~n17084 & n17087;
  assign n9791 = x75 & x94;
  assign n9792 = n9790 & n9791;
  assign n9793 = n9790 | n9791;
  assign n9794 = ~n9792 & n9793;
  assign n9795 = n17066 & n9794;
  assign n9796 = n17066 | n9794;
  assign n9797 = ~n9795 & n9796;
  assign n9798 = x74 & x95;
  assign n9799 = n9797 & n9798;
  assign n9800 = n9797 | n9798;
  assign n9801 = ~n9799 & n9800;
  assign n14333 = n9622 | n9624;
  assign n14365 = n9801 & n14333;
  assign n14366 = n9622 & n9801;
  assign n14367 = (n14248 & n14365) | (n14248 & n14366) | (n14365 & n14366);
  assign n14368 = n9801 | n14333;
  assign n14369 = n9622 | n9801;
  assign n14370 = (n14248 & n14368) | (n14248 & n14369) | (n14368 & n14369);
  assign n9804 = ~n14367 & n14370;
  assign n9805 = x73 & x96;
  assign n9806 = n9804 & n9805;
  assign n9807 = n9804 | n9805;
  assign n9808 = ~n9806 & n9807;
  assign n14371 = n9629 & n9808;
  assign n14372 = (n9808 & n17046) | (n9808 & n14371) | (n17046 & n14371);
  assign n14373 = n9629 | n9808;
  assign n14374 = n17046 | n14373;
  assign n9811 = ~n14372 & n14374;
  assign n9812 = x72 & x97;
  assign n9813 = n9811 & n9812;
  assign n9814 = n9811 | n9812;
  assign n9815 = ~n9813 & n9814;
  assign n14375 = n9636 & n9815;
  assign n14376 = (n9815 & n14288) | (n9815 & n14375) | (n14288 & n14375);
  assign n14377 = n9636 | n9815;
  assign n14378 = n14288 | n14377;
  assign n9818 = ~n14376 & n14378;
  assign n9819 = x71 & x98;
  assign n9820 = n9818 & n9819;
  assign n9821 = n9818 | n9819;
  assign n9822 = ~n9820 & n9821;
  assign n14379 = n9643 & n9822;
  assign n14380 = (n9822 & n14292) | (n9822 & n14379) | (n14292 & n14379);
  assign n14381 = n9643 | n9822;
  assign n14382 = n14292 | n14381;
  assign n9825 = ~n14380 & n14382;
  assign n9826 = x70 & x99;
  assign n9827 = n9825 & n9826;
  assign n9828 = n9825 | n9826;
  assign n9829 = ~n9827 & n9828;
  assign n14383 = n9650 & n9829;
  assign n14384 = (n9829 & n14296) | (n9829 & n14383) | (n14296 & n14383);
  assign n14385 = n9650 | n9829;
  assign n14386 = n14296 | n14385;
  assign n9832 = ~n14384 & n14386;
  assign n9833 = x69 & x100;
  assign n9834 = n9832 & n9833;
  assign n9835 = n9832 | n9833;
  assign n9836 = ~n9834 & n9835;
  assign n14387 = n9657 & n9836;
  assign n14388 = (n9836 & n14300) | (n9836 & n14387) | (n14300 & n14387);
  assign n14389 = n9657 | n9836;
  assign n14390 = n14300 | n14389;
  assign n9839 = ~n14388 & n14390;
  assign n9840 = x68 & x101;
  assign n9841 = n9839 & n9840;
  assign n9842 = n9839 | n9840;
  assign n9843 = ~n9841 & n9842;
  assign n14391 = n9664 & n9843;
  assign n14392 = (n9843 & n14304) | (n9843 & n14391) | (n14304 & n14391);
  assign n14393 = n9664 | n9843;
  assign n14394 = n14304 | n14393;
  assign n9846 = ~n14392 & n14394;
  assign n9847 = x67 & x102;
  assign n9848 = n9846 & n9847;
  assign n9849 = n9846 | n9847;
  assign n9850 = ~n9848 & n9849;
  assign n14395 = n9671 & n9850;
  assign n14396 = (n9850 & n14308) | (n9850 & n14395) | (n14308 & n14395);
  assign n14397 = n9671 | n9850;
  assign n14398 = n14308 | n14397;
  assign n9853 = ~n14396 & n14398;
  assign n9854 = x66 & x103;
  assign n9855 = n9853 & n9854;
  assign n9856 = n9853 | n9854;
  assign n9857 = ~n9855 & n9856;
  assign n14399 = n9678 & n9857;
  assign n14400 = (n9857 & n14313) | (n9857 & n14399) | (n14313 & n14399);
  assign n14401 = n9678 | n9857;
  assign n14402 = n14313 | n14401;
  assign n9860 = ~n14400 & n14402;
  assign n9861 = x65 & x104;
  assign n9862 = n9860 & n9861;
  assign n9863 = n9860 | n9861;
  assign n9864 = ~n9862 & n9863;
  assign n14331 = n9685 | n9687;
  assign n14403 = n9864 & n14331;
  assign n14404 = n9685 & n9864;
  assign n14405 = (n14243 & n14403) | (n14243 & n14404) | (n14403 & n14404);
  assign n14406 = n9864 | n14331;
  assign n14407 = n9685 | n9864;
  assign n14408 = (n14243 & n14406) | (n14243 & n14407) | (n14406 & n14407);
  assign n9867 = ~n14405 & n14408;
  assign n9868 = x64 & x105;
  assign n9869 = n9867 & n9868;
  assign n9870 = n9867 | n9868;
  assign n9871 = ~n9869 & n9870;
  assign n14329 = n9692 | n9694;
  assign n17088 = n9871 & n14329;
  assign n17089 = n9692 & n9871;
  assign n17090 = (n14241 & n17088) | (n14241 & n17089) | (n17088 & n17089);
  assign n17091 = n9871 | n14329;
  assign n17092 = n9692 | n9871;
  assign n17093 = (n14241 & n17091) | (n14241 & n17092) | (n17091 & n17092);
  assign n9874 = ~n17090 & n17093;
  assign n9875 = x63 & x106;
  assign n9876 = n9874 & n9875;
  assign n9877 = n9874 | n9875;
  assign n9878 = ~n9876 & n9877;
  assign n14327 = n9699 | n9701;
  assign n17094 = n9878 & n14327;
  assign n17095 = n9699 & n9878;
  assign n17096 = (n14239 & n17094) | (n14239 & n17095) | (n17094 & n17095);
  assign n17097 = n9878 | n14327;
  assign n17098 = n9699 | n9878;
  assign n17099 = (n14239 & n17097) | (n14239 & n17098) | (n17097 & n17098);
  assign n9881 = ~n17096 & n17099;
  assign n9882 = x62 & x107;
  assign n9883 = n9881 & n9882;
  assign n9884 = n9881 | n9882;
  assign n9885 = ~n9883 & n9884;
  assign n9886 = n14326 & n9885;
  assign n9887 = n14326 | n9885;
  assign n9888 = ~n9886 & n9887;
  assign n9889 = x61 & x108;
  assign n9890 = n9888 & n9889;
  assign n9891 = n9888 | n9889;
  assign n9892 = ~n9890 & n9891;
  assign n9893 = n14324 & n9892;
  assign n9894 = n14324 | n9892;
  assign n9895 = ~n9893 & n9894;
  assign n9896 = x60 & x109;
  assign n9897 = n9895 & n9896;
  assign n9898 = n9895 | n9896;
  assign n9899 = ~n9897 & n9898;
  assign n9900 = n14322 & n9899;
  assign n9901 = n14322 | n9899;
  assign n9902 = ~n9900 & n9901;
  assign n9903 = x59 & x110;
  assign n9904 = n9902 & n9903;
  assign n9905 = n9902 | n9903;
  assign n9906 = ~n9904 & n9905;
  assign n9907 = n14320 & n9906;
  assign n9908 = n14320 | n9906;
  assign n9909 = ~n9907 & n9908;
  assign n9910 = x58 & x111;
  assign n9911 = n9909 & n9910;
  assign n9912 = n9909 | n9910;
  assign n9913 = ~n9911 & n9912;
  assign n9914 = n14318 & n9913;
  assign n9915 = n14318 | n9913;
  assign n9916 = ~n9914 & n9915;
  assign n14409 = n9911 | n9913;
  assign n14410 = (n9911 & n14318) | (n9911 & n14409) | (n14318 & n14409);
  assign n14411 = n9904 | n9906;
  assign n14412 = (n9904 & n14320) | (n9904 & n14411) | (n14320 & n14411);
  assign n14413 = n9897 | n9899;
  assign n14414 = (n9897 & n14322) | (n9897 & n14413) | (n14322 & n14413);
  assign n14415 = n9890 | n9892;
  assign n14416 = (n9890 & n14324) | (n9890 & n14415) | (n14324 & n14415);
  assign n14328 = (n9699 & n14239) | (n9699 & n14327) | (n14239 & n14327);
  assign n14330 = (n9692 & n14241) | (n9692 & n14329) | (n14241 & n14329);
  assign n14429 = n9785 | n9787;
  assign n17102 = n9608 | n9785;
  assign n17103 = (n9785 & n9787) | (n9785 & n17102) | (n9787 & n17102);
  assign n17104 = (n14274 & n14429) | (n14274 & n17103) | (n14429 & n17103);
  assign n17105 = (n14273 & n14429) | (n14273 & n17103) | (n14429 & n17103);
  assign n17106 = (n16962 & n17104) | (n16962 & n17105) | (n17104 & n17105);
  assign n9939 = x79 & x91;
  assign n14434 = n9766 | n14347;
  assign n17107 = (n9587 & n14347) | (n9587 & n14434) | (n14347 & n14434);
  assign n14436 = n9939 & n17107;
  assign n50026 = n9939 & n17073;
  assign n66410 = n9763 & n9939;
  assign n66411 = n17019 & n66410;
  assign n50028 = (n17013 & n50026) | (n17013 & n66411) | (n50026 & n66411);
  assign n17109 = (n9766 & n9939) | (n9766 & n50028) | (n9939 & n50028);
  assign n17110 = (n14264 & n14436) | (n14264 & n17109) | (n14436 & n17109);
  assign n17111 = (n14263 & n14436) | (n14263 & n17109) | (n14436 & n17109);
  assign n17112 = (n16967 & n17110) | (n16967 & n17111) | (n17110 & n17111);
  assign n14439 = n9939 | n17107;
  assign n50029 = n9939 | n17073;
  assign n66412 = n9763 | n9939;
  assign n66413 = (n9939 & n17019) | (n9939 & n66412) | (n17019 & n66412);
  assign n50031 = (n17013 & n50029) | (n17013 & n66413) | (n50029 & n66413);
  assign n17114 = n9766 | n50031;
  assign n17115 = (n14264 & n14439) | (n14264 & n17114) | (n14439 & n17114);
  assign n17116 = (n14263 & n14439) | (n14263 & n17114) | (n14439 & n17114);
  assign n17117 = (n16967 & n17115) | (n16967 & n17116) | (n17115 & n17116);
  assign n9942 = ~n17112 & n17117;
  assign n14443 = n9771 & n9942;
  assign n17118 = (n9773 & n9942) | (n9773 & n14443) | (n9942 & n14443);
  assign n14444 = (n17071 & n17118) | (n17071 & n14443) | (n17118 & n14443);
  assign n14446 = n9771 | n9942;
  assign n17119 = n9773 | n14446;
  assign n14447 = (n17071 & n17119) | (n17071 & n14446) | (n17119 & n14446);
  assign n9945 = ~n14444 & n14447;
  assign n9946 = x78 & x92;
  assign n9947 = n9945 & n9946;
  assign n9948 = n9945 | n9946;
  assign n9949 = ~n9947 & n9948;
  assign n14448 = n9778 & n9949;
  assign n17120 = (n9949 & n14356) | (n9949 & n14448) | (n14356 & n14448);
  assign n17121 = (n9949 & n14355) | (n9949 & n14448) | (n14355 & n14448);
  assign n17122 = (n17008 & n17120) | (n17008 & n17121) | (n17120 & n17121);
  assign n14450 = n9778 | n9949;
  assign n17123 = n14356 | n14450;
  assign n17124 = n14355 | n14450;
  assign n17125 = (n17008 & n17123) | (n17008 & n17124) | (n17123 & n17124);
  assign n9952 = ~n17122 & n17125;
  assign n9953 = x77 & x93;
  assign n9954 = n9952 & n9953;
  assign n9955 = n9952 | n9953;
  assign n9956 = ~n9954 & n9955;
  assign n9957 = n17106 & n9956;
  assign n9958 = n17106 | n9956;
  assign n9959 = ~n9957 & n9958;
  assign n9960 = x76 & x94;
  assign n9961 = n9959 & n9960;
  assign n9962 = n9959 | n9960;
  assign n9963 = ~n9961 & n9962;
  assign n14426 = n9792 | n9794;
  assign n14452 = n9963 & n14426;
  assign n14453 = n9792 & n9963;
  assign n14454 = (n17066 & n14452) | (n17066 & n14453) | (n14452 & n14453);
  assign n14455 = n9963 | n14426;
  assign n14456 = n9792 | n9963;
  assign n14457 = (n17066 & n14455) | (n17066 & n14456) | (n14455 & n14456);
  assign n9966 = ~n14454 & n14457;
  assign n9967 = x75 & x95;
  assign n9968 = n9966 & n9967;
  assign n9969 = n9966 | n9967;
  assign n9970 = ~n9968 & n9969;
  assign n14458 = n9799 & n9970;
  assign n17126 = (n9970 & n14366) | (n9970 & n14458) | (n14366 & n14458);
  assign n17127 = (n9970 & n14365) | (n9970 & n14458) | (n14365 & n14458);
  assign n17128 = (n14248 & n17126) | (n14248 & n17127) | (n17126 & n17127);
  assign n14460 = n9799 | n9970;
  assign n17129 = n14366 | n14460;
  assign n17130 = n14365 | n14460;
  assign n17131 = (n14248 & n17129) | (n14248 & n17130) | (n17129 & n17130);
  assign n9973 = ~n17128 & n17131;
  assign n9974 = x74 & x96;
  assign n9975 = n9973 & n9974;
  assign n9976 = n9973 | n9974;
  assign n9977 = ~n9975 & n9976;
  assign n14424 = n9806 | n9808;
  assign n17132 = n9977 & n14424;
  assign n17100 = n9629 | n9806;
  assign n17101 = (n9806 & n9808) | (n9806 & n17100) | (n9808 & n17100);
  assign n17133 = n9977 & n17101;
  assign n17134 = (n17046 & n17132) | (n17046 & n17133) | (n17132 & n17133);
  assign n17135 = n9977 | n14424;
  assign n17136 = n9977 | n17101;
  assign n17137 = (n17046 & n17135) | (n17046 & n17136) | (n17135 & n17136);
  assign n9980 = ~n17134 & n17137;
  assign n9981 = x73 & x97;
  assign n9982 = n9980 & n9981;
  assign n9983 = n9980 | n9981;
  assign n9984 = ~n9982 & n9983;
  assign n14462 = n9813 & n9984;
  assign n17138 = (n9984 & n14375) | (n9984 & n14462) | (n14375 & n14462);
  assign n17139 = (n9815 & n9984) | (n9815 & n14462) | (n9984 & n14462);
  assign n17140 = (n14288 & n17138) | (n14288 & n17139) | (n17138 & n17139);
  assign n14464 = n9813 | n9984;
  assign n17141 = n14375 | n14464;
  assign n17142 = n9815 | n14464;
  assign n17143 = (n14288 & n17141) | (n14288 & n17142) | (n17141 & n17142);
  assign n9987 = ~n17140 & n17143;
  assign n9988 = x72 & x98;
  assign n9989 = n9987 & n9988;
  assign n9990 = n9987 | n9988;
  assign n9991 = ~n9989 & n9990;
  assign n14466 = n9820 & n9991;
  assign n14467 = (n9991 & n14380) | (n9991 & n14466) | (n14380 & n14466);
  assign n14468 = n9820 | n9991;
  assign n14469 = n14380 | n14468;
  assign n9994 = ~n14467 & n14469;
  assign n9995 = x71 & x99;
  assign n9996 = n9994 & n9995;
  assign n9997 = n9994 | n9995;
  assign n9998 = ~n9996 & n9997;
  assign n14470 = n9827 & n9998;
  assign n14471 = (n9998 & n14384) | (n9998 & n14470) | (n14384 & n14470);
  assign n14472 = n9827 | n9998;
  assign n14473 = n14384 | n14472;
  assign n10001 = ~n14471 & n14473;
  assign n10002 = x70 & x100;
  assign n10003 = n10001 & n10002;
  assign n10004 = n10001 | n10002;
  assign n10005 = ~n10003 & n10004;
  assign n14474 = n9834 & n10005;
  assign n14475 = (n10005 & n14388) | (n10005 & n14474) | (n14388 & n14474);
  assign n14476 = n9834 | n10005;
  assign n14477 = n14388 | n14476;
  assign n10008 = ~n14475 & n14477;
  assign n10009 = x69 & x101;
  assign n10010 = n10008 & n10009;
  assign n10011 = n10008 | n10009;
  assign n10012 = ~n10010 & n10011;
  assign n14478 = n9841 & n10012;
  assign n14479 = (n10012 & n14392) | (n10012 & n14478) | (n14392 & n14478);
  assign n14480 = n9841 | n10012;
  assign n14481 = n14392 | n14480;
  assign n10015 = ~n14479 & n14481;
  assign n10016 = x68 & x102;
  assign n10017 = n10015 & n10016;
  assign n10018 = n10015 | n10016;
  assign n10019 = ~n10017 & n10018;
  assign n14482 = n9848 & n10019;
  assign n14483 = (n10019 & n14396) | (n10019 & n14482) | (n14396 & n14482);
  assign n14484 = n9848 | n10019;
  assign n14485 = n14396 | n14484;
  assign n10022 = ~n14483 & n14485;
  assign n10023 = x67 & x103;
  assign n10024 = n10022 & n10023;
  assign n10025 = n10022 | n10023;
  assign n10026 = ~n10024 & n10025;
  assign n14486 = n9855 & n10026;
  assign n14487 = (n10026 & n14400) | (n10026 & n14486) | (n14400 & n14486);
  assign n14488 = n9855 | n10026;
  assign n14489 = n14400 | n14488;
  assign n10029 = ~n14487 & n14489;
  assign n10030 = x66 & x104;
  assign n10031 = n10029 & n10030;
  assign n10032 = n10029 | n10030;
  assign n10033 = ~n10031 & n10032;
  assign n14490 = n9862 & n10033;
  assign n14491 = (n10033 & n14405) | (n10033 & n14490) | (n14405 & n14490);
  assign n14492 = n9862 | n10033;
  assign n14493 = n14405 | n14492;
  assign n10036 = ~n14491 & n14493;
  assign n10037 = x65 & x105;
  assign n10038 = n10036 & n10037;
  assign n10039 = n10036 | n10037;
  assign n10040 = ~n10038 & n10039;
  assign n14421 = n9869 | n9871;
  assign n14494 = n10040 & n14421;
  assign n14495 = n9869 & n10040;
  assign n14496 = (n14330 & n14494) | (n14330 & n14495) | (n14494 & n14495);
  assign n14497 = n10040 | n14421;
  assign n14498 = n9869 | n10040;
  assign n14499 = (n14330 & n14497) | (n14330 & n14498) | (n14497 & n14498);
  assign n10043 = ~n14496 & n14499;
  assign n10044 = x64 & x106;
  assign n10045 = n10043 & n10044;
  assign n10046 = n10043 | n10044;
  assign n10047 = ~n10045 & n10046;
  assign n14419 = n9876 | n9878;
  assign n17144 = n10047 & n14419;
  assign n17145 = n9876 & n10047;
  assign n17146 = (n14328 & n17144) | (n14328 & n17145) | (n17144 & n17145);
  assign n17147 = n10047 | n14419;
  assign n17148 = n9876 | n10047;
  assign n17149 = (n14328 & n17147) | (n14328 & n17148) | (n17147 & n17148);
  assign n10050 = ~n17146 & n17149;
  assign n10051 = x63 & x107;
  assign n10052 = n10050 & n10051;
  assign n10053 = n10050 | n10051;
  assign n10054 = ~n10052 & n10053;
  assign n14417 = n9883 | n9885;
  assign n17150 = n10054 & n14417;
  assign n17151 = n9883 & n10054;
  assign n17152 = (n14326 & n17150) | (n14326 & n17151) | (n17150 & n17151);
  assign n17153 = n10054 | n14417;
  assign n17154 = n9883 | n10054;
  assign n17155 = (n14326 & n17153) | (n14326 & n17154) | (n17153 & n17154);
  assign n10057 = ~n17152 & n17155;
  assign n10058 = x62 & x108;
  assign n10059 = n10057 & n10058;
  assign n10060 = n10057 | n10058;
  assign n10061 = ~n10059 & n10060;
  assign n10062 = n14416 & n10061;
  assign n10063 = n14416 | n10061;
  assign n10064 = ~n10062 & n10063;
  assign n10065 = x61 & x109;
  assign n10066 = n10064 & n10065;
  assign n10067 = n10064 | n10065;
  assign n10068 = ~n10066 & n10067;
  assign n10069 = n14414 & n10068;
  assign n10070 = n14414 | n10068;
  assign n10071 = ~n10069 & n10070;
  assign n10072 = x60 & x110;
  assign n10073 = n10071 & n10072;
  assign n10074 = n10071 | n10072;
  assign n10075 = ~n10073 & n10074;
  assign n10076 = n14412 & n10075;
  assign n10077 = n14412 | n10075;
  assign n10078 = ~n10076 & n10077;
  assign n10079 = x59 & x111;
  assign n10080 = n10078 & n10079;
  assign n10081 = n10078 | n10079;
  assign n10082 = ~n10080 & n10081;
  assign n10083 = n14410 & n10082;
  assign n10084 = n14410 | n10082;
  assign n10085 = ~n10083 & n10084;
  assign n14500 = n10080 | n10082;
  assign n14501 = (n10080 & n14410) | (n10080 & n14500) | (n14410 & n14500);
  assign n14502 = n10073 | n10075;
  assign n14503 = (n10073 & n14412) | (n10073 & n14502) | (n14412 & n14502);
  assign n14504 = n10066 | n10068;
  assign n14505 = (n10066 & n14414) | (n10066 & n14504) | (n14414 & n14504);
  assign n14418 = (n9883 & n14326) | (n9883 & n14417) | (n14326 & n14417);
  assign n14420 = (n9876 & n14328) | (n9876 & n14419) | (n14328 & n14419);
  assign n14425 = (n17046 & n17101) | (n17046 & n14424) | (n17101 & n14424);
  assign n14515 = n9968 | n9970;
  assign n17156 = n9799 | n9968;
  assign n17157 = (n9968 & n9970) | (n9968 & n17156) | (n9970 & n17156);
  assign n17158 = (n14366 & n14515) | (n14366 & n17157) | (n14515 & n17157);
  assign n17159 = (n14365 & n14515) | (n14365 & n17157) | (n14515 & n17157);
  assign n17160 = (n14248 & n17158) | (n14248 & n17159) | (n17158 & n17159);
  assign n14520 = n9947 | n9949;
  assign n17161 = n9778 | n9947;
  assign n17162 = (n9947 & n9949) | (n9947 & n17161) | (n9949 & n17161);
  assign n17163 = (n14356 & n14520) | (n14356 & n17162) | (n14520 & n17162);
  assign n17164 = (n14355 & n14520) | (n14355 & n17162) | (n14520 & n17162);
  assign n17165 = (n17008 & n17163) | (n17008 & n17164) | (n17163 & n17164);
  assign n10107 = x79 & x92;
  assign n14522 = n10107 & n17112;
  assign n17166 = (n10107 & n14522) | (n10107 & n17118) | (n14522 & n17118);
  assign n50032 = (n9942 & n10107) | (n9942 & n14522) | (n10107 & n14522);
  assign n66414 = n10107 & n17112;
  assign n50034 = (n9771 & n50032) | (n9771 & n66414) | (n50032 & n66414);
  assign n17168 = (n17071 & n17166) | (n17071 & n50034) | (n17166 & n50034);
  assign n14524 = n10107 | n17112;
  assign n17169 = n14524 | n17118;
  assign n50035 = n9942 | n14524;
  assign n50036 = (n9771 & n14524) | (n9771 & n50035) | (n14524 & n50035);
  assign n17171 = (n17071 & n17169) | (n17071 & n50036) | (n17169 & n50036);
  assign n10110 = ~n17168 & n17171;
  assign n10111 = n17165 & n10110;
  assign n10112 = n17165 | n10110;
  assign n10113 = ~n10111 & n10112;
  assign n10114 = x78 & x93;
  assign n10115 = n10113 & n10114;
  assign n10116 = n10113 | n10114;
  assign n10117 = ~n10115 & n10116;
  assign n14517 = n9954 | n9956;
  assign n14526 = n10117 & n14517;
  assign n14527 = n9954 & n10117;
  assign n14528 = (n17106 & n14526) | (n17106 & n14527) | (n14526 & n14527);
  assign n14529 = n10117 | n14517;
  assign n14530 = n9954 | n10117;
  assign n14531 = (n17106 & n14529) | (n17106 & n14530) | (n14529 & n14530);
  assign n10120 = ~n14528 & n14531;
  assign n10121 = x77 & x94;
  assign n10122 = n10120 & n10121;
  assign n10123 = n10120 | n10121;
  assign n10124 = ~n10122 & n10123;
  assign n14532 = n9961 & n10124;
  assign n17172 = (n10124 & n14453) | (n10124 & n14532) | (n14453 & n14532);
  assign n17173 = (n10124 & n14452) | (n10124 & n14532) | (n14452 & n14532);
  assign n17174 = (n17066 & n17172) | (n17066 & n17173) | (n17172 & n17173);
  assign n14534 = n9961 | n10124;
  assign n17175 = n14453 | n14534;
  assign n17176 = n14452 | n14534;
  assign n17177 = (n17066 & n17175) | (n17066 & n17176) | (n17175 & n17176);
  assign n10127 = ~n17174 & n17177;
  assign n10128 = x76 & x95;
  assign n10129 = n10127 & n10128;
  assign n10130 = n10127 | n10128;
  assign n10131 = ~n10129 & n10130;
  assign n10132 = n17160 & n10131;
  assign n10133 = n17160 | n10131;
  assign n10134 = ~n10132 & n10133;
  assign n10135 = x75 & x96;
  assign n10136 = n10134 & n10135;
  assign n10137 = n10134 | n10135;
  assign n10138 = ~n10136 & n10137;
  assign n14512 = n9975 | n9977;
  assign n14536 = n10138 & n14512;
  assign n14537 = n9975 & n10138;
  assign n14538 = (n14425 & n14536) | (n14425 & n14537) | (n14536 & n14537);
  assign n14539 = n10138 | n14512;
  assign n14540 = n9975 | n10138;
  assign n14541 = (n14425 & n14539) | (n14425 & n14540) | (n14539 & n14540);
  assign n10141 = ~n14538 & n14541;
  assign n10142 = x74 & x97;
  assign n10143 = n10141 & n10142;
  assign n10144 = n10141 | n10142;
  assign n10145 = ~n10143 & n10144;
  assign n14542 = n9982 & n10145;
  assign n14543 = (n10145 & n17140) | (n10145 & n14542) | (n17140 & n14542);
  assign n14544 = n9982 | n10145;
  assign n14545 = n17140 | n14544;
  assign n10148 = ~n14543 & n14545;
  assign n10149 = x73 & x98;
  assign n10150 = n10148 & n10149;
  assign n10151 = n10148 | n10149;
  assign n10152 = ~n10150 & n10151;
  assign n14546 = n9989 & n10152;
  assign n14547 = (n10152 & n14467) | (n10152 & n14546) | (n14467 & n14546);
  assign n14548 = n9989 | n10152;
  assign n14549 = n14467 | n14548;
  assign n10155 = ~n14547 & n14549;
  assign n10156 = x72 & x99;
  assign n10157 = n10155 & n10156;
  assign n10158 = n10155 | n10156;
  assign n10159 = ~n10157 & n10158;
  assign n14550 = n9996 & n10159;
  assign n14551 = (n10159 & n14471) | (n10159 & n14550) | (n14471 & n14550);
  assign n14552 = n9996 | n10159;
  assign n14553 = n14471 | n14552;
  assign n10162 = ~n14551 & n14553;
  assign n10163 = x71 & x100;
  assign n10164 = n10162 & n10163;
  assign n10165 = n10162 | n10163;
  assign n10166 = ~n10164 & n10165;
  assign n14554 = n10003 & n10166;
  assign n14555 = (n10166 & n14475) | (n10166 & n14554) | (n14475 & n14554);
  assign n14556 = n10003 | n10166;
  assign n14557 = n14475 | n14556;
  assign n10169 = ~n14555 & n14557;
  assign n10170 = x70 & x101;
  assign n10171 = n10169 & n10170;
  assign n10172 = n10169 | n10170;
  assign n10173 = ~n10171 & n10172;
  assign n14558 = n10010 & n10173;
  assign n14559 = (n10173 & n14479) | (n10173 & n14558) | (n14479 & n14558);
  assign n14560 = n10010 | n10173;
  assign n14561 = n14479 | n14560;
  assign n10176 = ~n14559 & n14561;
  assign n10177 = x69 & x102;
  assign n10178 = n10176 & n10177;
  assign n10179 = n10176 | n10177;
  assign n10180 = ~n10178 & n10179;
  assign n14562 = n10017 & n10180;
  assign n14563 = (n10180 & n14483) | (n10180 & n14562) | (n14483 & n14562);
  assign n14564 = n10017 | n10180;
  assign n14565 = n14483 | n14564;
  assign n10183 = ~n14563 & n14565;
  assign n10184 = x68 & x103;
  assign n10185 = n10183 & n10184;
  assign n10186 = n10183 | n10184;
  assign n10187 = ~n10185 & n10186;
  assign n14566 = n10024 & n10187;
  assign n14567 = (n10187 & n14487) | (n10187 & n14566) | (n14487 & n14566);
  assign n14568 = n10024 | n10187;
  assign n14569 = n14487 | n14568;
  assign n10190 = ~n14567 & n14569;
  assign n10191 = x67 & x104;
  assign n10192 = n10190 & n10191;
  assign n10193 = n10190 | n10191;
  assign n10194 = ~n10192 & n10193;
  assign n14570 = n10031 & n10194;
  assign n14571 = (n10194 & n14491) | (n10194 & n14570) | (n14491 & n14570);
  assign n14572 = n10031 | n10194;
  assign n14573 = n14491 | n14572;
  assign n10197 = ~n14571 & n14573;
  assign n10198 = x66 & x105;
  assign n10199 = n10197 & n10198;
  assign n10200 = n10197 | n10198;
  assign n10201 = ~n10199 & n10200;
  assign n14574 = n10038 & n10201;
  assign n14575 = (n10201 & n14496) | (n10201 & n14574) | (n14496 & n14574);
  assign n14576 = n10038 | n10201;
  assign n14577 = n14496 | n14576;
  assign n10204 = ~n14575 & n14577;
  assign n10205 = x65 & x106;
  assign n10206 = n10204 & n10205;
  assign n10207 = n10204 | n10205;
  assign n10208 = ~n10206 & n10207;
  assign n14510 = n10045 | n10047;
  assign n14578 = n10208 & n14510;
  assign n14579 = n10045 & n10208;
  assign n14580 = (n14420 & n14578) | (n14420 & n14579) | (n14578 & n14579);
  assign n14581 = n10208 | n14510;
  assign n14582 = n10045 | n10208;
  assign n14583 = (n14420 & n14581) | (n14420 & n14582) | (n14581 & n14582);
  assign n10211 = ~n14580 & n14583;
  assign n10212 = x64 & x107;
  assign n10213 = n10211 & n10212;
  assign n10214 = n10211 | n10212;
  assign n10215 = ~n10213 & n10214;
  assign n14508 = n10052 | n10054;
  assign n17178 = n10215 & n14508;
  assign n17179 = n10052 & n10215;
  assign n17180 = (n14418 & n17178) | (n14418 & n17179) | (n17178 & n17179);
  assign n17181 = n10215 | n14508;
  assign n17182 = n10052 | n10215;
  assign n17183 = (n14418 & n17181) | (n14418 & n17182) | (n17181 & n17182);
  assign n10218 = ~n17180 & n17183;
  assign n10219 = x63 & x108;
  assign n10220 = n10218 & n10219;
  assign n10221 = n10218 | n10219;
  assign n10222 = ~n10220 & n10221;
  assign n14506 = n10059 | n10061;
  assign n17184 = n10222 & n14506;
  assign n17185 = n10059 & n10222;
  assign n17186 = (n14416 & n17184) | (n14416 & n17185) | (n17184 & n17185);
  assign n17187 = n10222 | n14506;
  assign n17188 = n10059 | n10222;
  assign n17189 = (n14416 & n17187) | (n14416 & n17188) | (n17187 & n17188);
  assign n10225 = ~n17186 & n17189;
  assign n10226 = x62 & x109;
  assign n10227 = n10225 & n10226;
  assign n10228 = n10225 | n10226;
  assign n10229 = ~n10227 & n10228;
  assign n10230 = n14505 & n10229;
  assign n10231 = n14505 | n10229;
  assign n10232 = ~n10230 & n10231;
  assign n10233 = x61 & x110;
  assign n10234 = n10232 & n10233;
  assign n10235 = n10232 | n10233;
  assign n10236 = ~n10234 & n10235;
  assign n10237 = n14503 & n10236;
  assign n10238 = n14503 | n10236;
  assign n10239 = ~n10237 & n10238;
  assign n10240 = x60 & x111;
  assign n10241 = n10239 & n10240;
  assign n10242 = n10239 | n10240;
  assign n10243 = ~n10241 & n10242;
  assign n10244 = n14501 & n10243;
  assign n10245 = n14501 | n10243;
  assign n10246 = ~n10244 & n10245;
  assign n14584 = n10241 | n10243;
  assign n14585 = (n10241 & n14501) | (n10241 & n14584) | (n14501 & n14584);
  assign n14586 = n10234 | n10236;
  assign n14587 = (n10234 & n14503) | (n10234 & n14586) | (n14503 & n14586);
  assign n14507 = (n10059 & n14416) | (n10059 & n14506) | (n14416 & n14506);
  assign n14509 = (n10052 & n14418) | (n10052 & n14508) | (n14418 & n14508);
  assign n14600 = n10122 | n10124;
  assign n17192 = n9961 | n10122;
  assign n17193 = (n10122 & n10124) | (n10122 & n17192) | (n10124 & n17192);
  assign n17194 = (n14453 & n14600) | (n14453 & n17193) | (n14600 & n17193);
  assign n17195 = (n14452 & n14600) | (n14452 & n17193) | (n14600 & n17193);
  assign n17196 = (n17066 & n17194) | (n17066 & n17195) | (n17194 & n17195);
  assign n10267 = x79 & x93;
  assign n50040 = n10107 & n10267;
  assign n66415 = n17112 & n50040;
  assign n50041 = (n17118 & n66415) | (n17118 & n50040) | (n66415 & n50040);
  assign n50037 = n10267 & n50034;
  assign n50038 = (n17071 & n50041) | (n17071 & n50037) | (n50041 & n50037);
  assign n17198 = (n10110 & n10267) | (n10110 & n50038) | (n10267 & n50038);
  assign n17200 = n10267 & n50034;
  assign n17201 = (n17071 & n50041) | (n17071 & n17200) | (n50041 & n17200);
  assign n14606 = (n17165 & n17198) | (n17165 & n17201) | (n17198 & n17201);
  assign n50045 = n10107 | n10267;
  assign n66416 = (n10267 & n17112) | (n10267 & n50045) | (n17112 & n50045);
  assign n50046 = (n17118 & n66416) | (n17118 & n50045) | (n66416 & n50045);
  assign n50042 = n10267 | n50034;
  assign n50043 = (n17071 & n50046) | (n17071 & n50042) | (n50046 & n50042);
  assign n17203 = n10110 | n50043;
  assign n17205 = n10267 | n50034;
  assign n17206 = (n17071 & n50046) | (n17071 & n17205) | (n50046 & n17205);
  assign n14609 = (n17165 & n17203) | (n17165 & n17206) | (n17203 & n17206);
  assign n10270 = ~n14606 & n14609;
  assign n14610 = n10115 & n10270;
  assign n17207 = (n10270 & n14527) | (n10270 & n14610) | (n14527 & n14610);
  assign n17208 = (n10270 & n14526) | (n10270 & n14610) | (n14526 & n14610);
  assign n17209 = (n17106 & n17207) | (n17106 & n17208) | (n17207 & n17208);
  assign n14612 = n10115 | n10270;
  assign n17210 = n14527 | n14612;
  assign n17211 = n14526 | n14612;
  assign n17212 = (n17106 & n17210) | (n17106 & n17211) | (n17210 & n17211);
  assign n10273 = ~n17209 & n17212;
  assign n10274 = x78 & x94;
  assign n10275 = n10273 & n10274;
  assign n10276 = n10273 | n10274;
  assign n10277 = ~n10275 & n10276;
  assign n10278 = n17196 & n10277;
  assign n10279 = n17196 | n10277;
  assign n10280 = ~n10278 & n10279;
  assign n10281 = x77 & x95;
  assign n10282 = n10280 & n10281;
  assign n10283 = n10280 | n10281;
  assign n10284 = ~n10282 & n10283;
  assign n14597 = n10129 | n10131;
  assign n14614 = n10284 & n14597;
  assign n14615 = n10129 & n10284;
  assign n14616 = (n17160 & n14614) | (n17160 & n14615) | (n14614 & n14615);
  assign n14617 = n10284 | n14597;
  assign n14618 = n10129 | n10284;
  assign n14619 = (n17160 & n14617) | (n17160 & n14618) | (n14617 & n14618);
  assign n10287 = ~n14616 & n14619;
  assign n10288 = x76 & x96;
  assign n10289 = n10287 & n10288;
  assign n10290 = n10287 | n10288;
  assign n10291 = ~n10289 & n10290;
  assign n14620 = n10136 & n10291;
  assign n17213 = (n10291 & n14537) | (n10291 & n14620) | (n14537 & n14620);
  assign n17214 = (n10291 & n14536) | (n10291 & n14620) | (n14536 & n14620);
  assign n17215 = (n14425 & n17213) | (n14425 & n17214) | (n17213 & n17214);
  assign n14622 = n10136 | n10291;
  assign n17216 = n14537 | n14622;
  assign n17217 = n14536 | n14622;
  assign n17218 = (n14425 & n17216) | (n14425 & n17217) | (n17216 & n17217);
  assign n10294 = ~n17215 & n17218;
  assign n10295 = x75 & x97;
  assign n10296 = n10294 & n10295;
  assign n10297 = n10294 | n10295;
  assign n10298 = ~n10296 & n10297;
  assign n14595 = n10143 | n10145;
  assign n17219 = n10298 & n14595;
  assign n17190 = n9982 | n10143;
  assign n17191 = (n10143 & n10145) | (n10143 & n17190) | (n10145 & n17190);
  assign n17220 = n10298 & n17191;
  assign n17221 = (n17140 & n17219) | (n17140 & n17220) | (n17219 & n17220);
  assign n17222 = n10298 | n14595;
  assign n17223 = n10298 | n17191;
  assign n17224 = (n17140 & n17222) | (n17140 & n17223) | (n17222 & n17223);
  assign n10301 = ~n17221 & n17224;
  assign n10302 = x74 & x98;
  assign n10303 = n10301 & n10302;
  assign n10304 = n10301 | n10302;
  assign n10305 = ~n10303 & n10304;
  assign n14624 = n10150 & n10305;
  assign n17225 = (n10305 & n14546) | (n10305 & n14624) | (n14546 & n14624);
  assign n17226 = (n10152 & n10305) | (n10152 & n14624) | (n10305 & n14624);
  assign n17227 = (n14467 & n17225) | (n14467 & n17226) | (n17225 & n17226);
  assign n14626 = n10150 | n10305;
  assign n17228 = n14546 | n14626;
  assign n17229 = n10152 | n14626;
  assign n17230 = (n14467 & n17228) | (n14467 & n17229) | (n17228 & n17229);
  assign n10308 = ~n17227 & n17230;
  assign n10309 = x73 & x99;
  assign n10310 = n10308 & n10309;
  assign n10311 = n10308 | n10309;
  assign n10312 = ~n10310 & n10311;
  assign n14628 = n10157 & n10312;
  assign n14629 = (n10312 & n14551) | (n10312 & n14628) | (n14551 & n14628);
  assign n14630 = n10157 | n10312;
  assign n14631 = n14551 | n14630;
  assign n10315 = ~n14629 & n14631;
  assign n10316 = x72 & x100;
  assign n10317 = n10315 & n10316;
  assign n10318 = n10315 | n10316;
  assign n10319 = ~n10317 & n10318;
  assign n14632 = n10164 & n10319;
  assign n14633 = (n10319 & n14555) | (n10319 & n14632) | (n14555 & n14632);
  assign n14634 = n10164 | n10319;
  assign n14635 = n14555 | n14634;
  assign n10322 = ~n14633 & n14635;
  assign n10323 = x71 & x101;
  assign n10324 = n10322 & n10323;
  assign n10325 = n10322 | n10323;
  assign n10326 = ~n10324 & n10325;
  assign n14636 = n10171 & n10326;
  assign n14637 = (n10326 & n14559) | (n10326 & n14636) | (n14559 & n14636);
  assign n14638 = n10171 | n10326;
  assign n14639 = n14559 | n14638;
  assign n10329 = ~n14637 & n14639;
  assign n10330 = x70 & x102;
  assign n10331 = n10329 & n10330;
  assign n10332 = n10329 | n10330;
  assign n10333 = ~n10331 & n10332;
  assign n14640 = n10178 & n10333;
  assign n14641 = (n10333 & n14563) | (n10333 & n14640) | (n14563 & n14640);
  assign n14642 = n10178 | n10333;
  assign n14643 = n14563 | n14642;
  assign n10336 = ~n14641 & n14643;
  assign n10337 = x69 & x103;
  assign n10338 = n10336 & n10337;
  assign n10339 = n10336 | n10337;
  assign n10340 = ~n10338 & n10339;
  assign n14644 = n10185 & n10340;
  assign n14645 = (n10340 & n14567) | (n10340 & n14644) | (n14567 & n14644);
  assign n14646 = n10185 | n10340;
  assign n14647 = n14567 | n14646;
  assign n10343 = ~n14645 & n14647;
  assign n10344 = x68 & x104;
  assign n10345 = n10343 & n10344;
  assign n10346 = n10343 | n10344;
  assign n10347 = ~n10345 & n10346;
  assign n14648 = n10192 & n10347;
  assign n14649 = (n10347 & n14571) | (n10347 & n14648) | (n14571 & n14648);
  assign n14650 = n10192 | n10347;
  assign n14651 = n14571 | n14650;
  assign n10350 = ~n14649 & n14651;
  assign n10351 = x67 & x105;
  assign n10352 = n10350 & n10351;
  assign n10353 = n10350 | n10351;
  assign n10354 = ~n10352 & n10353;
  assign n14652 = n10199 & n10354;
  assign n14653 = (n10354 & n14575) | (n10354 & n14652) | (n14575 & n14652);
  assign n14654 = n10199 | n10354;
  assign n14655 = n14575 | n14654;
  assign n10357 = ~n14653 & n14655;
  assign n10358 = x66 & x106;
  assign n10359 = n10357 & n10358;
  assign n10360 = n10357 | n10358;
  assign n10361 = ~n10359 & n10360;
  assign n14656 = n10206 & n10361;
  assign n14657 = (n10361 & n14580) | (n10361 & n14656) | (n14580 & n14656);
  assign n14658 = n10206 | n10361;
  assign n14659 = n14580 | n14658;
  assign n10364 = ~n14657 & n14659;
  assign n10365 = x65 & x107;
  assign n10366 = n10364 & n10365;
  assign n10367 = n10364 | n10365;
  assign n10368 = ~n10366 & n10367;
  assign n14592 = n10213 | n10215;
  assign n14660 = n10368 & n14592;
  assign n14661 = n10213 & n10368;
  assign n14662 = (n14509 & n14660) | (n14509 & n14661) | (n14660 & n14661);
  assign n14663 = n10368 | n14592;
  assign n14664 = n10213 | n10368;
  assign n14665 = (n14509 & n14663) | (n14509 & n14664) | (n14663 & n14664);
  assign n10371 = ~n14662 & n14665;
  assign n10372 = x64 & x108;
  assign n10373 = n10371 & n10372;
  assign n10374 = n10371 | n10372;
  assign n10375 = ~n10373 & n10374;
  assign n14590 = n10220 | n10222;
  assign n17231 = n10375 & n14590;
  assign n17232 = n10220 & n10375;
  assign n17233 = (n14507 & n17231) | (n14507 & n17232) | (n17231 & n17232);
  assign n17234 = n10375 | n14590;
  assign n17235 = n10220 | n10375;
  assign n17236 = (n14507 & n17234) | (n14507 & n17235) | (n17234 & n17235);
  assign n10378 = ~n17233 & n17236;
  assign n10379 = x63 & x109;
  assign n10380 = n10378 & n10379;
  assign n10381 = n10378 | n10379;
  assign n10382 = ~n10380 & n10381;
  assign n14588 = n10227 | n10229;
  assign n17237 = n10382 & n14588;
  assign n17238 = n10227 & n10382;
  assign n17239 = (n14505 & n17237) | (n14505 & n17238) | (n17237 & n17238);
  assign n17240 = n10382 | n14588;
  assign n17241 = n10227 | n10382;
  assign n17242 = (n14505 & n17240) | (n14505 & n17241) | (n17240 & n17241);
  assign n10385 = ~n17239 & n17242;
  assign n10386 = x62 & x110;
  assign n10387 = n10385 & n10386;
  assign n10388 = n10385 | n10386;
  assign n10389 = ~n10387 & n10388;
  assign n10390 = n14587 & n10389;
  assign n10391 = n14587 | n10389;
  assign n10392 = ~n10390 & n10391;
  assign n10393 = x61 & x111;
  assign n10394 = n10392 & n10393;
  assign n10395 = n10392 | n10393;
  assign n10396 = ~n10394 & n10395;
  assign n10397 = n14585 & n10396;
  assign n10398 = n14585 | n10396;
  assign n10399 = ~n10397 & n10398;
  assign n14666 = n10394 | n10396;
  assign n14667 = (n10394 & n14585) | (n10394 & n14666) | (n14585 & n14666);
  assign n14589 = (n10227 & n14505) | (n10227 & n14588) | (n14505 & n14588);
  assign n14591 = (n10220 & n14507) | (n10220 & n14590) | (n14507 & n14590);
  assign n14596 = (n17140 & n17191) | (n17140 & n14595) | (n17191 & n14595);
  assign n14677 = n10289 | n10291;
  assign n17243 = n10136 | n10289;
  assign n17244 = (n10289 & n10291) | (n10289 & n17243) | (n10291 & n17243);
  assign n17245 = (n14537 & n14677) | (n14537 & n17244) | (n14677 & n17244);
  assign n17246 = (n14536 & n14677) | (n14536 & n17244) | (n14677 & n17244);
  assign n17247 = (n14425 & n17245) | (n14425 & n17246) | (n17245 & n17246);
  assign n10419 = x79 & x94;
  assign n14682 = n10270 | n14606;
  assign n17248 = (n10115 & n14606) | (n10115 & n14682) | (n14606 & n14682);
  assign n14684 = n10419 & n17248;
  assign n66417 = n10419 & n50038;
  assign n66418 = n10267 & n10419;
  assign n66419 = (n10110 & n66417) | (n10110 & n66418) | (n66417 & n66418);
  assign n66420 = n10419 & n50041;
  assign n66421 = n10419 & n17200;
  assign n66422 = (n17071 & n66420) | (n17071 & n66421) | (n66420 & n66421);
  assign n50049 = (n17165 & n66419) | (n17165 & n66422) | (n66419 & n66422);
  assign n17250 = (n10270 & n10419) | (n10270 & n50049) | (n10419 & n50049);
  assign n17251 = (n14527 & n14684) | (n14527 & n17250) | (n14684 & n17250);
  assign n17252 = (n14526 & n14684) | (n14526 & n17250) | (n14684 & n17250);
  assign n17253 = (n17106 & n17251) | (n17106 & n17252) | (n17251 & n17252);
  assign n14687 = n10419 | n17248;
  assign n66423 = n10419 | n50038;
  assign n66424 = n10267 | n10419;
  assign n66425 = (n10110 & n66423) | (n10110 & n66424) | (n66423 & n66424);
  assign n66426 = n10419 | n50041;
  assign n66427 = n10419 | n17200;
  assign n66428 = (n17071 & n66426) | (n17071 & n66427) | (n66426 & n66427);
  assign n50052 = (n17165 & n66425) | (n17165 & n66428) | (n66425 & n66428);
  assign n17255 = n10270 | n50052;
  assign n17256 = (n14527 & n14687) | (n14527 & n17255) | (n14687 & n17255);
  assign n17257 = (n14526 & n14687) | (n14526 & n17255) | (n14687 & n17255);
  assign n17258 = (n17106 & n17256) | (n17106 & n17257) | (n17256 & n17257);
  assign n10422 = ~n17253 & n17258;
  assign n14691 = n10275 & n10422;
  assign n17259 = (n10277 & n10422) | (n10277 & n14691) | (n10422 & n14691);
  assign n14692 = (n17196 & n17259) | (n17196 & n14691) | (n17259 & n14691);
  assign n14694 = n10275 | n10422;
  assign n17260 = n10277 | n14694;
  assign n14695 = (n17196 & n17260) | (n17196 & n14694) | (n17260 & n14694);
  assign n10425 = ~n14692 & n14695;
  assign n10426 = x78 & x95;
  assign n10427 = n10425 & n10426;
  assign n10428 = n10425 | n10426;
  assign n10429 = ~n10427 & n10428;
  assign n14696 = n10282 & n10429;
  assign n17261 = (n10429 & n14615) | (n10429 & n14696) | (n14615 & n14696);
  assign n17262 = (n10429 & n14614) | (n10429 & n14696) | (n14614 & n14696);
  assign n17263 = (n17160 & n17261) | (n17160 & n17262) | (n17261 & n17262);
  assign n14698 = n10282 | n10429;
  assign n17264 = n14615 | n14698;
  assign n17265 = n14614 | n14698;
  assign n17266 = (n17160 & n17264) | (n17160 & n17265) | (n17264 & n17265);
  assign n10432 = ~n17263 & n17266;
  assign n10433 = x77 & x96;
  assign n10434 = n10432 & n10433;
  assign n10435 = n10432 | n10433;
  assign n10436 = ~n10434 & n10435;
  assign n10437 = n17247 & n10436;
  assign n10438 = n17247 | n10436;
  assign n10439 = ~n10437 & n10438;
  assign n10440 = x76 & x97;
  assign n10441 = n10439 & n10440;
  assign n10442 = n10439 | n10440;
  assign n10443 = ~n10441 & n10442;
  assign n14674 = n10296 | n10298;
  assign n14700 = n10443 & n14674;
  assign n14701 = n10296 & n10443;
  assign n14702 = (n14596 & n14700) | (n14596 & n14701) | (n14700 & n14701);
  assign n14703 = n10443 | n14674;
  assign n14704 = n10296 | n10443;
  assign n14705 = (n14596 & n14703) | (n14596 & n14704) | (n14703 & n14704);
  assign n10446 = ~n14702 & n14705;
  assign n10447 = x75 & x98;
  assign n10448 = n10446 & n10447;
  assign n10449 = n10446 | n10447;
  assign n10450 = ~n10448 & n10449;
  assign n14706 = n10303 & n10450;
  assign n14707 = (n10450 & n17227) | (n10450 & n14706) | (n17227 & n14706);
  assign n14708 = n10303 | n10450;
  assign n14709 = n17227 | n14708;
  assign n10453 = ~n14707 & n14709;
  assign n10454 = x74 & x99;
  assign n10455 = n10453 & n10454;
  assign n10456 = n10453 | n10454;
  assign n10457 = ~n10455 & n10456;
  assign n14710 = n10310 & n10457;
  assign n14711 = (n10457 & n14629) | (n10457 & n14710) | (n14629 & n14710);
  assign n14712 = n10310 | n10457;
  assign n14713 = n14629 | n14712;
  assign n10460 = ~n14711 & n14713;
  assign n10461 = x73 & x100;
  assign n10462 = n10460 & n10461;
  assign n10463 = n10460 | n10461;
  assign n10464 = ~n10462 & n10463;
  assign n14714 = n10317 & n10464;
  assign n14715 = (n10464 & n14633) | (n10464 & n14714) | (n14633 & n14714);
  assign n14716 = n10317 | n10464;
  assign n14717 = n14633 | n14716;
  assign n10467 = ~n14715 & n14717;
  assign n10468 = x72 & x101;
  assign n10469 = n10467 & n10468;
  assign n10470 = n10467 | n10468;
  assign n10471 = ~n10469 & n10470;
  assign n14718 = n10324 & n10471;
  assign n14719 = (n10471 & n14637) | (n10471 & n14718) | (n14637 & n14718);
  assign n14720 = n10324 | n10471;
  assign n14721 = n14637 | n14720;
  assign n10474 = ~n14719 & n14721;
  assign n10475 = x71 & x102;
  assign n10476 = n10474 & n10475;
  assign n10477 = n10474 | n10475;
  assign n10478 = ~n10476 & n10477;
  assign n14722 = n10331 & n10478;
  assign n14723 = (n10478 & n14641) | (n10478 & n14722) | (n14641 & n14722);
  assign n14724 = n10331 | n10478;
  assign n14725 = n14641 | n14724;
  assign n10481 = ~n14723 & n14725;
  assign n10482 = x70 & x103;
  assign n10483 = n10481 & n10482;
  assign n10484 = n10481 | n10482;
  assign n10485 = ~n10483 & n10484;
  assign n14726 = n10338 & n10485;
  assign n14727 = (n10485 & n14645) | (n10485 & n14726) | (n14645 & n14726);
  assign n14728 = n10338 | n10485;
  assign n14729 = n14645 | n14728;
  assign n10488 = ~n14727 & n14729;
  assign n10489 = x69 & x104;
  assign n10490 = n10488 & n10489;
  assign n10491 = n10488 | n10489;
  assign n10492 = ~n10490 & n10491;
  assign n14730 = n10345 & n10492;
  assign n14731 = (n10492 & n14649) | (n10492 & n14730) | (n14649 & n14730);
  assign n14732 = n10345 | n10492;
  assign n14733 = n14649 | n14732;
  assign n10495 = ~n14731 & n14733;
  assign n10496 = x68 & x105;
  assign n10497 = n10495 & n10496;
  assign n10498 = n10495 | n10496;
  assign n10499 = ~n10497 & n10498;
  assign n14734 = n10352 & n10499;
  assign n14735 = (n10499 & n14653) | (n10499 & n14734) | (n14653 & n14734);
  assign n14736 = n10352 | n10499;
  assign n14737 = n14653 | n14736;
  assign n10502 = ~n14735 & n14737;
  assign n10503 = x67 & x106;
  assign n10504 = n10502 & n10503;
  assign n10505 = n10502 | n10503;
  assign n10506 = ~n10504 & n10505;
  assign n14738 = n10359 & n10506;
  assign n14739 = (n10506 & n14657) | (n10506 & n14738) | (n14657 & n14738);
  assign n14740 = n10359 | n10506;
  assign n14741 = n14657 | n14740;
  assign n10509 = ~n14739 & n14741;
  assign n10510 = x66 & x107;
  assign n10511 = n10509 & n10510;
  assign n10512 = n10509 | n10510;
  assign n10513 = ~n10511 & n10512;
  assign n14742 = n10366 & n10513;
  assign n14743 = (n10513 & n14662) | (n10513 & n14742) | (n14662 & n14742);
  assign n14744 = n10366 | n10513;
  assign n14745 = n14662 | n14744;
  assign n10516 = ~n14743 & n14745;
  assign n10517 = x65 & x108;
  assign n10518 = n10516 & n10517;
  assign n10519 = n10516 | n10517;
  assign n10520 = ~n10518 & n10519;
  assign n14672 = n10373 | n10375;
  assign n14746 = n10520 & n14672;
  assign n14747 = n10373 & n10520;
  assign n14748 = (n14591 & n14746) | (n14591 & n14747) | (n14746 & n14747);
  assign n14749 = n10520 | n14672;
  assign n14750 = n10373 | n10520;
  assign n14751 = (n14591 & n14749) | (n14591 & n14750) | (n14749 & n14750);
  assign n10523 = ~n14748 & n14751;
  assign n10524 = x64 & x109;
  assign n10525 = n10523 & n10524;
  assign n10526 = n10523 | n10524;
  assign n10527 = ~n10525 & n10526;
  assign n14670 = n10380 | n10382;
  assign n17267 = n10527 & n14670;
  assign n17268 = n10380 & n10527;
  assign n17269 = (n14589 & n17267) | (n14589 & n17268) | (n17267 & n17268);
  assign n17270 = n10527 | n14670;
  assign n17271 = n10380 | n10527;
  assign n17272 = (n14589 & n17270) | (n14589 & n17271) | (n17270 & n17271);
  assign n10530 = ~n17269 & n17272;
  assign n10531 = x63 & x110;
  assign n10532 = n10530 & n10531;
  assign n10533 = n10530 | n10531;
  assign n10534 = ~n10532 & n10533;
  assign n14668 = n10387 | n10389;
  assign n17273 = n10534 & n14668;
  assign n17274 = n10387 & n10534;
  assign n17275 = (n14587 & n17273) | (n14587 & n17274) | (n17273 & n17274);
  assign n17276 = n10534 | n14668;
  assign n17277 = n10387 | n10534;
  assign n17278 = (n14587 & n17276) | (n14587 & n17277) | (n17276 & n17277);
  assign n10537 = ~n17275 & n17278;
  assign n10538 = x62 & x111;
  assign n10539 = n10537 & n10538;
  assign n10540 = n10537 | n10538;
  assign n10541 = ~n10539 & n10540;
  assign n10542 = n14667 & n10541;
  assign n10543 = n14667 | n10541;
  assign n10544 = ~n10542 & n10543;
  assign n14669 = (n10387 & n14587) | (n10387 & n14668) | (n14587 & n14668);
  assign n14671 = (n10380 & n14589) | (n10380 & n14670) | (n14589 & n14670);
  assign n14764 = n10427 | n10429;
  assign n17281 = n10282 | n10427;
  assign n17282 = (n10427 & n10429) | (n10427 & n17281) | (n10429 & n17281);
  assign n17283 = (n14615 & n14764) | (n14615 & n17282) | (n14764 & n17282);
  assign n17284 = (n14614 & n14764) | (n14614 & n17282) | (n14764 & n17282);
  assign n17285 = (n17160 & n17283) | (n17160 & n17284) | (n17283 & n17284);
  assign n10563 = x79 & x95;
  assign n14766 = n10563 & n17253;
  assign n17286 = (n10563 & n14766) | (n10563 & n17259) | (n14766 & n17259);
  assign n50053 = (n10422 & n10563) | (n10422 & n14766) | (n10563 & n14766);
  assign n66429 = n10563 & n17253;
  assign n50055 = (n10275 & n50053) | (n10275 & n66429) | (n50053 & n66429);
  assign n17288 = (n17196 & n17286) | (n17196 & n50055) | (n17286 & n50055);
  assign n14768 = n10563 | n17253;
  assign n17289 = n14768 | n17259;
  assign n50056 = n10422 | n14768;
  assign n50057 = (n10275 & n14768) | (n10275 & n50056) | (n14768 & n50056);
  assign n17291 = (n17196 & n17289) | (n17196 & n50057) | (n17289 & n50057);
  assign n10566 = ~n17288 & n17291;
  assign n10567 = n17285 & n10566;
  assign n10568 = n17285 | n10566;
  assign n10569 = ~n10567 & n10568;
  assign n10570 = x78 & x96;
  assign n10571 = n10569 & n10570;
  assign n10572 = n10569 | n10570;
  assign n10573 = ~n10571 & n10572;
  assign n14761 = n10434 | n10436;
  assign n14770 = n10573 & n14761;
  assign n14771 = n10434 & n10573;
  assign n14772 = (n17247 & n14770) | (n17247 & n14771) | (n14770 & n14771);
  assign n14773 = n10573 | n14761;
  assign n14774 = n10434 | n10573;
  assign n14775 = (n17247 & n14773) | (n17247 & n14774) | (n14773 & n14774);
  assign n10576 = ~n14772 & n14775;
  assign n10577 = x77 & x97;
  assign n10578 = n10576 & n10577;
  assign n10579 = n10576 | n10577;
  assign n10580 = ~n10578 & n10579;
  assign n14776 = n10441 & n10580;
  assign n17292 = (n10580 & n14701) | (n10580 & n14776) | (n14701 & n14776);
  assign n17293 = (n10580 & n14700) | (n10580 & n14776) | (n14700 & n14776);
  assign n17294 = (n14596 & n17292) | (n14596 & n17293) | (n17292 & n17293);
  assign n14778 = n10441 | n10580;
  assign n17295 = n14701 | n14778;
  assign n17296 = n14700 | n14778;
  assign n17297 = (n14596 & n17295) | (n14596 & n17296) | (n17295 & n17296);
  assign n10583 = ~n17294 & n17297;
  assign n10584 = x76 & x98;
  assign n10585 = n10583 & n10584;
  assign n10586 = n10583 | n10584;
  assign n10587 = ~n10585 & n10586;
  assign n14759 = n10448 | n10450;
  assign n17298 = n10587 & n14759;
  assign n17279 = n10303 | n10448;
  assign n17280 = (n10448 & n10450) | (n10448 & n17279) | (n10450 & n17279);
  assign n17299 = n10587 & n17280;
  assign n17300 = (n17227 & n17298) | (n17227 & n17299) | (n17298 & n17299);
  assign n17301 = n10587 | n14759;
  assign n17302 = n10587 | n17280;
  assign n17303 = (n17227 & n17301) | (n17227 & n17302) | (n17301 & n17302);
  assign n10590 = ~n17300 & n17303;
  assign n10591 = x75 & x99;
  assign n10592 = n10590 & n10591;
  assign n10593 = n10590 | n10591;
  assign n10594 = ~n10592 & n10593;
  assign n14780 = n10455 & n10594;
  assign n17304 = (n10594 & n14710) | (n10594 & n14780) | (n14710 & n14780);
  assign n17305 = (n10457 & n10594) | (n10457 & n14780) | (n10594 & n14780);
  assign n17306 = (n14629 & n17304) | (n14629 & n17305) | (n17304 & n17305);
  assign n14782 = n10455 | n10594;
  assign n17307 = n14710 | n14782;
  assign n17308 = n10457 | n14782;
  assign n17309 = (n14629 & n17307) | (n14629 & n17308) | (n17307 & n17308);
  assign n10597 = ~n17306 & n17309;
  assign n10598 = x74 & x100;
  assign n10599 = n10597 & n10598;
  assign n10600 = n10597 | n10598;
  assign n10601 = ~n10599 & n10600;
  assign n14784 = n10462 & n10601;
  assign n14785 = (n10601 & n14715) | (n10601 & n14784) | (n14715 & n14784);
  assign n14786 = n10462 | n10601;
  assign n14787 = n14715 | n14786;
  assign n10604 = ~n14785 & n14787;
  assign n10605 = x73 & x101;
  assign n10606 = n10604 & n10605;
  assign n10607 = n10604 | n10605;
  assign n10608 = ~n10606 & n10607;
  assign n14788 = n10469 & n10608;
  assign n14789 = (n10608 & n14719) | (n10608 & n14788) | (n14719 & n14788);
  assign n14790 = n10469 | n10608;
  assign n14791 = n14719 | n14790;
  assign n10611 = ~n14789 & n14791;
  assign n10612 = x72 & x102;
  assign n10613 = n10611 & n10612;
  assign n10614 = n10611 | n10612;
  assign n10615 = ~n10613 & n10614;
  assign n14792 = n10476 & n10615;
  assign n14793 = (n10615 & n14723) | (n10615 & n14792) | (n14723 & n14792);
  assign n14794 = n10476 | n10615;
  assign n14795 = n14723 | n14794;
  assign n10618 = ~n14793 & n14795;
  assign n10619 = x71 & x103;
  assign n10620 = n10618 & n10619;
  assign n10621 = n10618 | n10619;
  assign n10622 = ~n10620 & n10621;
  assign n14796 = n10483 & n10622;
  assign n14797 = (n10622 & n14727) | (n10622 & n14796) | (n14727 & n14796);
  assign n14798 = n10483 | n10622;
  assign n14799 = n14727 | n14798;
  assign n10625 = ~n14797 & n14799;
  assign n10626 = x70 & x104;
  assign n10627 = n10625 & n10626;
  assign n10628 = n10625 | n10626;
  assign n10629 = ~n10627 & n10628;
  assign n14800 = n10490 & n10629;
  assign n14801 = (n10629 & n14731) | (n10629 & n14800) | (n14731 & n14800);
  assign n14802 = n10490 | n10629;
  assign n14803 = n14731 | n14802;
  assign n10632 = ~n14801 & n14803;
  assign n10633 = x69 & x105;
  assign n10634 = n10632 & n10633;
  assign n10635 = n10632 | n10633;
  assign n10636 = ~n10634 & n10635;
  assign n14804 = n10497 & n10636;
  assign n14805 = (n10636 & n14735) | (n10636 & n14804) | (n14735 & n14804);
  assign n14806 = n10497 | n10636;
  assign n14807 = n14735 | n14806;
  assign n10639 = ~n14805 & n14807;
  assign n10640 = x68 & x106;
  assign n10641 = n10639 & n10640;
  assign n10642 = n10639 | n10640;
  assign n10643 = ~n10641 & n10642;
  assign n14808 = n10504 & n10643;
  assign n14809 = (n10643 & n14739) | (n10643 & n14808) | (n14739 & n14808);
  assign n14810 = n10504 | n10643;
  assign n14811 = n14739 | n14810;
  assign n10646 = ~n14809 & n14811;
  assign n10647 = x67 & x107;
  assign n10648 = n10646 & n10647;
  assign n10649 = n10646 | n10647;
  assign n10650 = ~n10648 & n10649;
  assign n14812 = n10511 & n10650;
  assign n14813 = (n10650 & n14743) | (n10650 & n14812) | (n14743 & n14812);
  assign n14814 = n10511 | n10650;
  assign n14815 = n14743 | n14814;
  assign n10653 = ~n14813 & n14815;
  assign n10654 = x66 & x108;
  assign n10655 = n10653 & n10654;
  assign n10656 = n10653 | n10654;
  assign n10657 = ~n10655 & n10656;
  assign n14816 = n10518 & n10657;
  assign n14817 = (n10657 & n14748) | (n10657 & n14816) | (n14748 & n14816);
  assign n14818 = n10518 | n10657;
  assign n14819 = n14748 | n14818;
  assign n10660 = ~n14817 & n14819;
  assign n10661 = x65 & x109;
  assign n10662 = n10660 & n10661;
  assign n10663 = n10660 | n10661;
  assign n10664 = ~n10662 & n10663;
  assign n14756 = n10525 | n10527;
  assign n14820 = n10664 & n14756;
  assign n14821 = n10525 & n10664;
  assign n14822 = (n14671 & n14820) | (n14671 & n14821) | (n14820 & n14821);
  assign n14823 = n10664 | n14756;
  assign n14824 = n10525 | n10664;
  assign n14825 = (n14671 & n14823) | (n14671 & n14824) | (n14823 & n14824);
  assign n10667 = ~n14822 & n14825;
  assign n10668 = x64 & x110;
  assign n10669 = n10667 & n10668;
  assign n10670 = n10667 | n10668;
  assign n10671 = ~n10669 & n10670;
  assign n14754 = n10532 | n10534;
  assign n17310 = n10671 & n14754;
  assign n17311 = n10532 & n10671;
  assign n17312 = (n14669 & n17310) | (n14669 & n17311) | (n17310 & n17311);
  assign n17313 = n10671 | n14754;
  assign n17314 = n10532 | n10671;
  assign n17315 = (n14669 & n17313) | (n14669 & n17314) | (n17313 & n17314);
  assign n10674 = ~n17312 & n17315;
  assign n10675 = x63 & x111;
  assign n10676 = n10674 & n10675;
  assign n10677 = n10674 | n10675;
  assign n10678 = ~n10676 & n10677;
  assign n14752 = n10539 | n10541;
  assign n17316 = n10678 & n14752;
  assign n17317 = n10539 & n10678;
  assign n17318 = (n14667 & n17316) | (n14667 & n17317) | (n17316 & n17317);
  assign n17319 = n10678 | n14752;
  assign n17320 = n10539 | n10678;
  assign n17321 = (n14667 & n17319) | (n14667 & n17320) | (n17319 & n17320);
  assign n10681 = ~n17318 & n17321;
  assign n14753 = (n10539 & n14667) | (n10539 & n14752) | (n14667 & n14752);
  assign n14755 = (n10532 & n14669) | (n10532 & n14754) | (n14669 & n14754);
  assign n14760 = (n17227 & n17280) | (n17227 & n14759) | (n17280 & n14759);
  assign n14833 = n10578 | n10580;
  assign n17322 = n10441 | n10578;
  assign n17323 = (n10578 & n10580) | (n10578 & n17322) | (n10580 & n17322);
  assign n17324 = (n14701 & n14833) | (n14701 & n17323) | (n14833 & n17323);
  assign n17325 = (n14700 & n14833) | (n14700 & n17323) | (n14833 & n17323);
  assign n17326 = (n14596 & n17324) | (n14596 & n17325) | (n17324 & n17325);
  assign n10699 = x79 & x96;
  assign n50061 = n10563 & n10699;
  assign n66430 = n17253 & n50061;
  assign n50062 = (n17259 & n66430) | (n17259 & n50061) | (n66430 & n50061);
  assign n50058 = n10699 & n50055;
  assign n50059 = (n17196 & n50062) | (n17196 & n50058) | (n50062 & n50058);
  assign n17328 = (n10566 & n10699) | (n10566 & n50059) | (n10699 & n50059);
  assign n17330 = n10699 & n50055;
  assign n17331 = (n17196 & n50062) | (n17196 & n17330) | (n50062 & n17330);
  assign n14839 = (n17285 & n17328) | (n17285 & n17331) | (n17328 & n17331);
  assign n50066 = n10563 | n10699;
  assign n66431 = (n10699 & n17253) | (n10699 & n50066) | (n17253 & n50066);
  assign n50067 = (n17259 & n66431) | (n17259 & n50066) | (n66431 & n50066);
  assign n50063 = n10699 | n50055;
  assign n50064 = (n17196 & n50067) | (n17196 & n50063) | (n50067 & n50063);
  assign n17333 = n10566 | n50064;
  assign n17335 = n10699 | n50055;
  assign n17336 = (n17196 & n50067) | (n17196 & n17335) | (n50067 & n17335);
  assign n14842 = (n17285 & n17333) | (n17285 & n17336) | (n17333 & n17336);
  assign n10702 = ~n14839 & n14842;
  assign n14843 = n10571 & n10702;
  assign n17337 = (n10702 & n14771) | (n10702 & n14843) | (n14771 & n14843);
  assign n17338 = (n10702 & n14770) | (n10702 & n14843) | (n14770 & n14843);
  assign n17339 = (n17247 & n17337) | (n17247 & n17338) | (n17337 & n17338);
  assign n14845 = n10571 | n10702;
  assign n17340 = n14771 | n14845;
  assign n17341 = n14770 | n14845;
  assign n17342 = (n17247 & n17340) | (n17247 & n17341) | (n17340 & n17341);
  assign n10705 = ~n17339 & n17342;
  assign n10706 = x78 & x97;
  assign n10707 = n10705 & n10706;
  assign n10708 = n10705 | n10706;
  assign n10709 = ~n10707 & n10708;
  assign n10710 = n17326 & n10709;
  assign n10711 = n17326 | n10709;
  assign n10712 = ~n10710 & n10711;
  assign n10713 = x77 & x98;
  assign n10714 = n10712 & n10713;
  assign n10715 = n10712 | n10713;
  assign n10716 = ~n10714 & n10715;
  assign n14830 = n10585 | n10587;
  assign n14847 = n10716 & n14830;
  assign n14848 = n10585 & n10716;
  assign n14849 = (n14760 & n14847) | (n14760 & n14848) | (n14847 & n14848);
  assign n14850 = n10716 | n14830;
  assign n14851 = n10585 | n10716;
  assign n14852 = (n14760 & n14850) | (n14760 & n14851) | (n14850 & n14851);
  assign n10719 = ~n14849 & n14852;
  assign n10720 = x76 & x99;
  assign n10721 = n10719 & n10720;
  assign n10722 = n10719 | n10720;
  assign n10723 = ~n10721 & n10722;
  assign n14853 = n10592 & n10723;
  assign n14854 = (n10723 & n17306) | (n10723 & n14853) | (n17306 & n14853);
  assign n14855 = n10592 | n10723;
  assign n14856 = n17306 | n14855;
  assign n10726 = ~n14854 & n14856;
  assign n10727 = x75 & x100;
  assign n10728 = n10726 & n10727;
  assign n10729 = n10726 | n10727;
  assign n10730 = ~n10728 & n10729;
  assign n14857 = n10599 & n10730;
  assign n14858 = (n10730 & n14785) | (n10730 & n14857) | (n14785 & n14857);
  assign n14859 = n10599 | n10730;
  assign n14860 = n14785 | n14859;
  assign n10733 = ~n14858 & n14860;
  assign n10734 = x74 & x101;
  assign n10735 = n10733 & n10734;
  assign n10736 = n10733 | n10734;
  assign n10737 = ~n10735 & n10736;
  assign n14861 = n10606 & n10737;
  assign n14862 = (n10737 & n14789) | (n10737 & n14861) | (n14789 & n14861);
  assign n14863 = n10606 | n10737;
  assign n14864 = n14789 | n14863;
  assign n10740 = ~n14862 & n14864;
  assign n10741 = x73 & x102;
  assign n10742 = n10740 & n10741;
  assign n10743 = n10740 | n10741;
  assign n10744 = ~n10742 & n10743;
  assign n14865 = n10613 & n10744;
  assign n14866 = (n10744 & n14793) | (n10744 & n14865) | (n14793 & n14865);
  assign n14867 = n10613 | n10744;
  assign n14868 = n14793 | n14867;
  assign n10747 = ~n14866 & n14868;
  assign n10748 = x72 & x103;
  assign n10749 = n10747 & n10748;
  assign n10750 = n10747 | n10748;
  assign n10751 = ~n10749 & n10750;
  assign n14869 = n10620 & n10751;
  assign n14870 = (n10751 & n14797) | (n10751 & n14869) | (n14797 & n14869);
  assign n14871 = n10620 | n10751;
  assign n14872 = n14797 | n14871;
  assign n10754 = ~n14870 & n14872;
  assign n10755 = x71 & x104;
  assign n10756 = n10754 & n10755;
  assign n10757 = n10754 | n10755;
  assign n10758 = ~n10756 & n10757;
  assign n14873 = n10627 & n10758;
  assign n14874 = (n10758 & n14801) | (n10758 & n14873) | (n14801 & n14873);
  assign n14875 = n10627 | n10758;
  assign n14876 = n14801 | n14875;
  assign n10761 = ~n14874 & n14876;
  assign n10762 = x70 & x105;
  assign n10763 = n10761 & n10762;
  assign n10764 = n10761 | n10762;
  assign n10765 = ~n10763 & n10764;
  assign n14877 = n10634 & n10765;
  assign n14878 = (n10765 & n14805) | (n10765 & n14877) | (n14805 & n14877);
  assign n14879 = n10634 | n10765;
  assign n14880 = n14805 | n14879;
  assign n10768 = ~n14878 & n14880;
  assign n10769 = x69 & x106;
  assign n10770 = n10768 & n10769;
  assign n10771 = n10768 | n10769;
  assign n10772 = ~n10770 & n10771;
  assign n14881 = n10641 & n10772;
  assign n14882 = (n10772 & n14809) | (n10772 & n14881) | (n14809 & n14881);
  assign n14883 = n10641 | n10772;
  assign n14884 = n14809 | n14883;
  assign n10775 = ~n14882 & n14884;
  assign n10776 = x68 & x107;
  assign n10777 = n10775 & n10776;
  assign n10778 = n10775 | n10776;
  assign n10779 = ~n10777 & n10778;
  assign n14885 = n10648 & n10779;
  assign n14886 = (n10779 & n14813) | (n10779 & n14885) | (n14813 & n14885);
  assign n14887 = n10648 | n10779;
  assign n14888 = n14813 | n14887;
  assign n10782 = ~n14886 & n14888;
  assign n10783 = x67 & x108;
  assign n10784 = n10782 & n10783;
  assign n10785 = n10782 | n10783;
  assign n10786 = ~n10784 & n10785;
  assign n14889 = n10655 & n10786;
  assign n14890 = (n10786 & n14817) | (n10786 & n14889) | (n14817 & n14889);
  assign n14891 = n10655 | n10786;
  assign n14892 = n14817 | n14891;
  assign n10789 = ~n14890 & n14892;
  assign n10790 = x66 & x109;
  assign n10791 = n10789 & n10790;
  assign n10792 = n10789 | n10790;
  assign n10793 = ~n10791 & n10792;
  assign n14893 = n10662 & n10793;
  assign n14894 = (n10793 & n14822) | (n10793 & n14893) | (n14822 & n14893);
  assign n14895 = n10662 | n10793;
  assign n14896 = n14822 | n14895;
  assign n10796 = ~n14894 & n14896;
  assign n10797 = x65 & x110;
  assign n10798 = n10796 & n10797;
  assign n10799 = n10796 | n10797;
  assign n10800 = ~n10798 & n10799;
  assign n14828 = n10669 | n10671;
  assign n14897 = n10800 & n14828;
  assign n14898 = n10669 & n10800;
  assign n14899 = (n14755 & n14897) | (n14755 & n14898) | (n14897 & n14898);
  assign n14900 = n10800 | n14828;
  assign n14901 = n10669 | n10800;
  assign n14902 = (n14755 & n14900) | (n14755 & n14901) | (n14900 & n14901);
  assign n10803 = ~n14899 & n14902;
  assign n10804 = x64 & x111;
  assign n10805 = n10803 & n10804;
  assign n10806 = n10803 | n10804;
  assign n10807 = ~n10805 & n10806;
  assign n14826 = n10676 | n10678;
  assign n17343 = n10807 & n14826;
  assign n17344 = n10676 & n10807;
  assign n17345 = (n14753 & n17343) | (n14753 & n17344) | (n17343 & n17344);
  assign n17346 = n10807 | n14826;
  assign n17347 = n10676 | n10807;
  assign n17348 = (n14753 & n17346) | (n14753 & n17347) | (n17346 & n17347);
  assign n10810 = ~n17345 & n17348;
  assign n14827 = (n10676 & n14753) | (n10676 & n14826) | (n14753 & n14826);
  assign n10827 = x79 & x97;
  assign n14911 = n10702 | n14839;
  assign n17351 = (n10571 & n14839) | (n10571 & n14911) | (n14839 & n14911);
  assign n14913 = n10827 & n17351;
  assign n66432 = n10827 & n50059;
  assign n66433 = n10699 & n10827;
  assign n66434 = (n10566 & n66432) | (n10566 & n66433) | (n66432 & n66433);
  assign n66435 = n10827 & n50062;
  assign n66436 = n10827 & n17330;
  assign n66437 = (n17196 & n66435) | (n17196 & n66436) | (n66435 & n66436);
  assign n50070 = (n17285 & n66434) | (n17285 & n66437) | (n66434 & n66437);
  assign n17353 = (n10702 & n10827) | (n10702 & n50070) | (n10827 & n50070);
  assign n17354 = (n14771 & n14913) | (n14771 & n17353) | (n14913 & n17353);
  assign n17355 = (n14770 & n14913) | (n14770 & n17353) | (n14913 & n17353);
  assign n17356 = (n17247 & n17354) | (n17247 & n17355) | (n17354 & n17355);
  assign n14916 = n10827 | n17351;
  assign n66438 = n10827 | n50059;
  assign n66439 = n10699 | n10827;
  assign n66440 = (n10566 & n66438) | (n10566 & n66439) | (n66438 & n66439);
  assign n66441 = n10827 | n50062;
  assign n66442 = n10827 | n17330;
  assign n66443 = (n17196 & n66441) | (n17196 & n66442) | (n66441 & n66442);
  assign n50073 = (n17285 & n66440) | (n17285 & n66443) | (n66440 & n66443);
  assign n17358 = n10702 | n50073;
  assign n17359 = (n14771 & n14916) | (n14771 & n17358) | (n14916 & n17358);
  assign n17360 = (n14770 & n14916) | (n14770 & n17358) | (n14916 & n17358);
  assign n17361 = (n17247 & n17359) | (n17247 & n17360) | (n17359 & n17360);
  assign n10830 = ~n17356 & n17361;
  assign n14920 = n10707 & n10830;
  assign n17362 = (n10709 & n10830) | (n10709 & n14920) | (n10830 & n14920);
  assign n14921 = (n17326 & n17362) | (n17326 & n14920) | (n17362 & n14920);
  assign n14923 = n10707 | n10830;
  assign n17363 = n10709 | n14923;
  assign n14924 = (n17326 & n17363) | (n17326 & n14923) | (n17363 & n14923);
  assign n10833 = ~n14921 & n14924;
  assign n10834 = x78 & x98;
  assign n10835 = n10833 & n10834;
  assign n10836 = n10833 | n10834;
  assign n10837 = ~n10835 & n10836;
  assign n14925 = n10714 & n10837;
  assign n17364 = (n10837 & n14848) | (n10837 & n14925) | (n14848 & n14925);
  assign n17365 = (n10837 & n14847) | (n10837 & n14925) | (n14847 & n14925);
  assign n17366 = (n14760 & n17364) | (n14760 & n17365) | (n17364 & n17365);
  assign n14927 = n10714 | n10837;
  assign n17367 = n14848 | n14927;
  assign n17368 = n14847 | n14927;
  assign n17369 = (n14760 & n17367) | (n14760 & n17368) | (n17367 & n17368);
  assign n10840 = ~n17366 & n17369;
  assign n10841 = x77 & x99;
  assign n10842 = n10840 & n10841;
  assign n10843 = n10840 | n10841;
  assign n10844 = ~n10842 & n10843;
  assign n14906 = n10721 | n10723;
  assign n17370 = n10844 & n14906;
  assign n17349 = n10592 | n10721;
  assign n17350 = (n10721 & n10723) | (n10721 & n17349) | (n10723 & n17349);
  assign n17371 = n10844 & n17350;
  assign n17372 = (n17306 & n17370) | (n17306 & n17371) | (n17370 & n17371);
  assign n17373 = n10844 | n14906;
  assign n17374 = n10844 | n17350;
  assign n17375 = (n17306 & n17373) | (n17306 & n17374) | (n17373 & n17374);
  assign n10847 = ~n17372 & n17375;
  assign n10848 = x76 & x100;
  assign n10849 = n10847 & n10848;
  assign n10850 = n10847 | n10848;
  assign n10851 = ~n10849 & n10850;
  assign n14929 = n10728 & n10851;
  assign n17376 = (n10851 & n14857) | (n10851 & n14929) | (n14857 & n14929);
  assign n17377 = (n10730 & n10851) | (n10730 & n14929) | (n10851 & n14929);
  assign n17378 = (n14785 & n17376) | (n14785 & n17377) | (n17376 & n17377);
  assign n14931 = n10728 | n10851;
  assign n17379 = n14857 | n14931;
  assign n17380 = n10730 | n14931;
  assign n17381 = (n14785 & n17379) | (n14785 & n17380) | (n17379 & n17380);
  assign n10854 = ~n17378 & n17381;
  assign n10855 = x75 & x101;
  assign n10856 = n10854 & n10855;
  assign n10857 = n10854 | n10855;
  assign n10858 = ~n10856 & n10857;
  assign n14933 = n10735 & n10858;
  assign n14934 = (n10858 & n14862) | (n10858 & n14933) | (n14862 & n14933);
  assign n14935 = n10735 | n10858;
  assign n14936 = n14862 | n14935;
  assign n10861 = ~n14934 & n14936;
  assign n10862 = x74 & x102;
  assign n10863 = n10861 & n10862;
  assign n10864 = n10861 | n10862;
  assign n10865 = ~n10863 & n10864;
  assign n14937 = n10742 & n10865;
  assign n14938 = (n10865 & n14866) | (n10865 & n14937) | (n14866 & n14937);
  assign n14939 = n10742 | n10865;
  assign n14940 = n14866 | n14939;
  assign n10868 = ~n14938 & n14940;
  assign n10869 = x73 & x103;
  assign n10870 = n10868 & n10869;
  assign n10871 = n10868 | n10869;
  assign n10872 = ~n10870 & n10871;
  assign n14941 = n10749 & n10872;
  assign n14942 = (n10872 & n14870) | (n10872 & n14941) | (n14870 & n14941);
  assign n14943 = n10749 | n10872;
  assign n14944 = n14870 | n14943;
  assign n10875 = ~n14942 & n14944;
  assign n10876 = x72 & x104;
  assign n10877 = n10875 & n10876;
  assign n10878 = n10875 | n10876;
  assign n10879 = ~n10877 & n10878;
  assign n14945 = n10756 & n10879;
  assign n14946 = (n10879 & n14874) | (n10879 & n14945) | (n14874 & n14945);
  assign n14947 = n10756 | n10879;
  assign n14948 = n14874 | n14947;
  assign n10882 = ~n14946 & n14948;
  assign n10883 = x71 & x105;
  assign n10884 = n10882 & n10883;
  assign n10885 = n10882 | n10883;
  assign n10886 = ~n10884 & n10885;
  assign n14949 = n10763 & n10886;
  assign n14950 = (n10886 & n14878) | (n10886 & n14949) | (n14878 & n14949);
  assign n14951 = n10763 | n10886;
  assign n14952 = n14878 | n14951;
  assign n10889 = ~n14950 & n14952;
  assign n10890 = x70 & x106;
  assign n10891 = n10889 & n10890;
  assign n10892 = n10889 | n10890;
  assign n10893 = ~n10891 & n10892;
  assign n14953 = n10770 & n10893;
  assign n14954 = (n10893 & n14882) | (n10893 & n14953) | (n14882 & n14953);
  assign n14955 = n10770 | n10893;
  assign n14956 = n14882 | n14955;
  assign n10896 = ~n14954 & n14956;
  assign n10897 = x69 & x107;
  assign n10898 = n10896 & n10897;
  assign n10899 = n10896 | n10897;
  assign n10900 = ~n10898 & n10899;
  assign n14957 = n10777 & n10900;
  assign n14958 = (n10900 & n14886) | (n10900 & n14957) | (n14886 & n14957);
  assign n14959 = n10777 | n10900;
  assign n14960 = n14886 | n14959;
  assign n10903 = ~n14958 & n14960;
  assign n10904 = x68 & x108;
  assign n10905 = n10903 & n10904;
  assign n10906 = n10903 | n10904;
  assign n10907 = ~n10905 & n10906;
  assign n14961 = n10784 & n10907;
  assign n14962 = (n10907 & n14890) | (n10907 & n14961) | (n14890 & n14961);
  assign n14963 = n10784 | n10907;
  assign n14964 = n14890 | n14963;
  assign n10910 = ~n14962 & n14964;
  assign n10911 = x67 & x109;
  assign n10912 = n10910 & n10911;
  assign n10913 = n10910 | n10911;
  assign n10914 = ~n10912 & n10913;
  assign n14965 = n10791 & n10914;
  assign n14966 = (n10914 & n14894) | (n10914 & n14965) | (n14894 & n14965);
  assign n14967 = n10791 | n10914;
  assign n14968 = n14894 | n14967;
  assign n10917 = ~n14966 & n14968;
  assign n10918 = x66 & x110;
  assign n10919 = n10917 & n10918;
  assign n10920 = n10917 | n10918;
  assign n10921 = ~n10919 & n10920;
  assign n14969 = n10798 & n10921;
  assign n14970 = (n10921 & n14899) | (n10921 & n14969) | (n14899 & n14969);
  assign n14971 = n10798 | n10921;
  assign n14972 = n14899 | n14971;
  assign n10924 = ~n14970 & n14972;
  assign n10925 = x65 & x111;
  assign n10926 = n10924 & n10925;
  assign n10927 = n10924 | n10925;
  assign n10928 = ~n10926 & n10927;
  assign n14903 = n10805 | n10807;
  assign n14973 = n10928 & n14903;
  assign n14974 = n10805 & n10928;
  assign n14975 = (n14827 & n14973) | (n14827 & n14974) | (n14973 & n14974);
  assign n14976 = n10928 | n14903;
  assign n14977 = n10805 | n10928;
  assign n14978 = (n14827 & n14976) | (n14827 & n14977) | (n14976 & n14977);
  assign n10931 = ~n14975 & n14978;
  assign n14907 = (n17306 & n17350) | (n17306 & n14906) | (n17350 & n14906);
  assign n14982 = n10835 | n10837;
  assign n17382 = n10714 | n10835;
  assign n17383 = (n10835 & n10837) | (n10835 & n17382) | (n10837 & n17382);
  assign n17384 = (n14848 & n14982) | (n14848 & n17383) | (n14982 & n17383);
  assign n17385 = (n14847 & n14982) | (n14847 & n17383) | (n14982 & n17383);
  assign n17386 = (n14760 & n17384) | (n14760 & n17385) | (n17384 & n17385);
  assign n10947 = x79 & x98;
  assign n14984 = n10947 & n17356;
  assign n17387 = (n10947 & n14984) | (n10947 & n17362) | (n14984 & n17362);
  assign n50074 = (n10830 & n10947) | (n10830 & n14984) | (n10947 & n14984);
  assign n66444 = n10947 & n17356;
  assign n50076 = (n10707 & n50074) | (n10707 & n66444) | (n50074 & n66444);
  assign n17389 = (n17326 & n17387) | (n17326 & n50076) | (n17387 & n50076);
  assign n14986 = n10947 | n17356;
  assign n17390 = n14986 | n17362;
  assign n50077 = n10830 | n14986;
  assign n50078 = (n10707 & n14986) | (n10707 & n50077) | (n14986 & n50077);
  assign n17392 = (n17326 & n17390) | (n17326 & n50078) | (n17390 & n50078);
  assign n10950 = ~n17389 & n17392;
  assign n10951 = n17386 & n10950;
  assign n10952 = n17386 | n10950;
  assign n10953 = ~n10951 & n10952;
  assign n10954 = x78 & x99;
  assign n10955 = n10953 & n10954;
  assign n10956 = n10953 | n10954;
  assign n10957 = ~n10955 & n10956;
  assign n14979 = n10842 | n10844;
  assign n14988 = n10957 & n14979;
  assign n14989 = n10842 & n10957;
  assign n14990 = (n14907 & n14988) | (n14907 & n14989) | (n14988 & n14989);
  assign n14991 = n10957 | n14979;
  assign n14992 = n10842 | n10957;
  assign n14993 = (n14907 & n14991) | (n14907 & n14992) | (n14991 & n14992);
  assign n10960 = ~n14990 & n14993;
  assign n10961 = x77 & x100;
  assign n10962 = n10960 & n10961;
  assign n10963 = n10960 | n10961;
  assign n10964 = ~n10962 & n10963;
  assign n14994 = n10849 & n10964;
  assign n14995 = (n10964 & n17378) | (n10964 & n14994) | (n17378 & n14994);
  assign n14996 = n10849 | n10964;
  assign n14997 = n17378 | n14996;
  assign n10967 = ~n14995 & n14997;
  assign n10968 = x76 & x101;
  assign n10969 = n10967 & n10968;
  assign n10970 = n10967 | n10968;
  assign n10971 = ~n10969 & n10970;
  assign n14998 = n10856 & n10971;
  assign n14999 = (n10971 & n14934) | (n10971 & n14998) | (n14934 & n14998);
  assign n15000 = n10856 | n10971;
  assign n15001 = n14934 | n15000;
  assign n10974 = ~n14999 & n15001;
  assign n10975 = x75 & x102;
  assign n10976 = n10974 & n10975;
  assign n10977 = n10974 | n10975;
  assign n10978 = ~n10976 & n10977;
  assign n15002 = n10863 & n10978;
  assign n15003 = (n10978 & n14938) | (n10978 & n15002) | (n14938 & n15002);
  assign n15004 = n10863 | n10978;
  assign n15005 = n14938 | n15004;
  assign n10981 = ~n15003 & n15005;
  assign n10982 = x74 & x103;
  assign n10983 = n10981 & n10982;
  assign n10984 = n10981 | n10982;
  assign n10985 = ~n10983 & n10984;
  assign n15006 = n10870 & n10985;
  assign n15007 = (n10985 & n14942) | (n10985 & n15006) | (n14942 & n15006);
  assign n15008 = n10870 | n10985;
  assign n15009 = n14942 | n15008;
  assign n10988 = ~n15007 & n15009;
  assign n10989 = x73 & x104;
  assign n10990 = n10988 & n10989;
  assign n10991 = n10988 | n10989;
  assign n10992 = ~n10990 & n10991;
  assign n15010 = n10877 & n10992;
  assign n15011 = (n10992 & n14946) | (n10992 & n15010) | (n14946 & n15010);
  assign n15012 = n10877 | n10992;
  assign n15013 = n14946 | n15012;
  assign n10995 = ~n15011 & n15013;
  assign n10996 = x72 & x105;
  assign n10997 = n10995 & n10996;
  assign n10998 = n10995 | n10996;
  assign n10999 = ~n10997 & n10998;
  assign n15014 = n10884 & n10999;
  assign n15015 = (n10999 & n14950) | (n10999 & n15014) | (n14950 & n15014);
  assign n15016 = n10884 | n10999;
  assign n15017 = n14950 | n15016;
  assign n11002 = ~n15015 & n15017;
  assign n11003 = x71 & x106;
  assign n11004 = n11002 & n11003;
  assign n11005 = n11002 | n11003;
  assign n11006 = ~n11004 & n11005;
  assign n15018 = n10891 & n11006;
  assign n15019 = (n11006 & n14954) | (n11006 & n15018) | (n14954 & n15018);
  assign n15020 = n10891 | n11006;
  assign n15021 = n14954 | n15020;
  assign n11009 = ~n15019 & n15021;
  assign n11010 = x70 & x107;
  assign n11011 = n11009 & n11010;
  assign n11012 = n11009 | n11010;
  assign n11013 = ~n11011 & n11012;
  assign n15022 = n10898 & n11013;
  assign n15023 = (n11013 & n14958) | (n11013 & n15022) | (n14958 & n15022);
  assign n15024 = n10898 | n11013;
  assign n15025 = n14958 | n15024;
  assign n11016 = ~n15023 & n15025;
  assign n11017 = x69 & x108;
  assign n11018 = n11016 & n11017;
  assign n11019 = n11016 | n11017;
  assign n11020 = ~n11018 & n11019;
  assign n15026 = n10905 & n11020;
  assign n15027 = (n11020 & n14962) | (n11020 & n15026) | (n14962 & n15026);
  assign n15028 = n10905 | n11020;
  assign n15029 = n14962 | n15028;
  assign n11023 = ~n15027 & n15029;
  assign n11024 = x68 & x109;
  assign n11025 = n11023 & n11024;
  assign n11026 = n11023 | n11024;
  assign n11027 = ~n11025 & n11026;
  assign n15030 = n10912 & n11027;
  assign n15031 = (n11027 & n14966) | (n11027 & n15030) | (n14966 & n15030);
  assign n15032 = n10912 | n11027;
  assign n15033 = n14966 | n15032;
  assign n11030 = ~n15031 & n15033;
  assign n11031 = x67 & x110;
  assign n11032 = n11030 & n11031;
  assign n11033 = n11030 | n11031;
  assign n11034 = ~n11032 & n11033;
  assign n15034 = n10919 & n11034;
  assign n15035 = (n11034 & n14970) | (n11034 & n15034) | (n14970 & n15034);
  assign n15036 = n10919 | n11034;
  assign n15037 = n14970 | n15036;
  assign n11037 = ~n15035 & n15037;
  assign n11038 = x66 & x111;
  assign n11039 = n11037 & n11038;
  assign n11040 = n11037 | n11038;
  assign n11041 = ~n11039 & n11040;
  assign n15038 = n10926 & n11041;
  assign n15039 = (n11041 & n14975) | (n11041 & n15038) | (n14975 & n15038);
  assign n15040 = n10926 | n11041;
  assign n15041 = n14975 | n15040;
  assign n11044 = ~n15039 & n15041;
  assign n11059 = x79 & x99;
  assign n50082 = n10947 & n11059;
  assign n66445 = n17356 & n50082;
  assign n50083 = (n17362 & n66445) | (n17362 & n50082) | (n66445 & n50082);
  assign n50079 = n11059 & n50076;
  assign n50080 = (n17326 & n50083) | (n17326 & n50079) | (n50083 & n50079);
  assign n17396 = (n10950 & n11059) | (n10950 & n50080) | (n11059 & n50080);
  assign n17398 = n11059 & n50076;
  assign n17399 = (n17326 & n50083) | (n17326 & n17398) | (n50083 & n17398);
  assign n15049 = (n17386 & n17396) | (n17386 & n17399) | (n17396 & n17399);
  assign n50087 = n10947 | n11059;
  assign n66446 = (n11059 & n17356) | (n11059 & n50087) | (n17356 & n50087);
  assign n50088 = (n17362 & n66446) | (n17362 & n50087) | (n66446 & n50087);
  assign n50084 = n11059 | n50076;
  assign n50085 = (n17326 & n50088) | (n17326 & n50084) | (n50088 & n50084);
  assign n17401 = n10950 | n50085;
  assign n17403 = n11059 | n50076;
  assign n17404 = (n17326 & n50088) | (n17326 & n17403) | (n50088 & n17403);
  assign n15052 = (n17386 & n17401) | (n17386 & n17404) | (n17401 & n17404);
  assign n11062 = ~n15049 & n15052;
  assign n15053 = n10955 & n11062;
  assign n17405 = (n11062 & n14989) | (n11062 & n15053) | (n14989 & n15053);
  assign n17406 = (n11062 & n14988) | (n11062 & n15053) | (n14988 & n15053);
  assign n17407 = (n14907 & n17405) | (n14907 & n17406) | (n17405 & n17406);
  assign n15055 = n10955 | n11062;
  assign n17408 = n14989 | n15055;
  assign n17409 = n14988 | n15055;
  assign n17410 = (n14907 & n17408) | (n14907 & n17409) | (n17408 & n17409);
  assign n11065 = ~n17407 & n17410;
  assign n11066 = x78 & x100;
  assign n11067 = n11065 & n11066;
  assign n11068 = n11065 | n11066;
  assign n11069 = ~n11067 & n11068;
  assign n15043 = n10962 | n10964;
  assign n17411 = n11069 & n15043;
  assign n17393 = n10849 | n10962;
  assign n17394 = (n10962 & n10964) | (n10962 & n17393) | (n10964 & n17393);
  assign n17412 = n11069 & n17394;
  assign n17413 = (n17378 & n17411) | (n17378 & n17412) | (n17411 & n17412);
  assign n17414 = n11069 | n15043;
  assign n17415 = n11069 | n17394;
  assign n17416 = (n17378 & n17414) | (n17378 & n17415) | (n17414 & n17415);
  assign n11072 = ~n17413 & n17416;
  assign n11073 = x77 & x101;
  assign n11074 = n11072 & n11073;
  assign n11075 = n11072 | n11073;
  assign n11076 = ~n11074 & n11075;
  assign n15057 = n10969 & n11076;
  assign n17417 = (n11076 & n14998) | (n11076 & n15057) | (n14998 & n15057);
  assign n17418 = (n10971 & n11076) | (n10971 & n15057) | (n11076 & n15057);
  assign n17419 = (n14934 & n17417) | (n14934 & n17418) | (n17417 & n17418);
  assign n15059 = n10969 | n11076;
  assign n17420 = n14998 | n15059;
  assign n17421 = n10971 | n15059;
  assign n17422 = (n14934 & n17420) | (n14934 & n17421) | (n17420 & n17421);
  assign n11079 = ~n17419 & n17422;
  assign n11080 = x76 & x102;
  assign n11081 = n11079 & n11080;
  assign n11082 = n11079 | n11080;
  assign n11083 = ~n11081 & n11082;
  assign n15061 = n10976 & n11083;
  assign n15062 = (n11083 & n15003) | (n11083 & n15061) | (n15003 & n15061);
  assign n15063 = n10976 | n11083;
  assign n15064 = n15003 | n15063;
  assign n11086 = ~n15062 & n15064;
  assign n11087 = x75 & x103;
  assign n11088 = n11086 & n11087;
  assign n11089 = n11086 | n11087;
  assign n11090 = ~n11088 & n11089;
  assign n15065 = n10983 & n11090;
  assign n15066 = (n11090 & n15007) | (n11090 & n15065) | (n15007 & n15065);
  assign n15067 = n10983 | n11090;
  assign n15068 = n15007 | n15067;
  assign n11093 = ~n15066 & n15068;
  assign n11094 = x74 & x104;
  assign n11095 = n11093 & n11094;
  assign n11096 = n11093 | n11094;
  assign n11097 = ~n11095 & n11096;
  assign n15069 = n10990 & n11097;
  assign n15070 = (n11097 & n15011) | (n11097 & n15069) | (n15011 & n15069);
  assign n15071 = n10990 | n11097;
  assign n15072 = n15011 | n15071;
  assign n11100 = ~n15070 & n15072;
  assign n11101 = x73 & x105;
  assign n11102 = n11100 & n11101;
  assign n11103 = n11100 | n11101;
  assign n11104 = ~n11102 & n11103;
  assign n15073 = n10997 & n11104;
  assign n15074 = (n11104 & n15015) | (n11104 & n15073) | (n15015 & n15073);
  assign n15075 = n10997 | n11104;
  assign n15076 = n15015 | n15075;
  assign n11107 = ~n15074 & n15076;
  assign n11108 = x72 & x106;
  assign n11109 = n11107 & n11108;
  assign n11110 = n11107 | n11108;
  assign n11111 = ~n11109 & n11110;
  assign n15077 = n11004 & n11111;
  assign n15078 = (n11111 & n15019) | (n11111 & n15077) | (n15019 & n15077);
  assign n15079 = n11004 | n11111;
  assign n15080 = n15019 | n15079;
  assign n11114 = ~n15078 & n15080;
  assign n11115 = x71 & x107;
  assign n11116 = n11114 & n11115;
  assign n11117 = n11114 | n11115;
  assign n11118 = ~n11116 & n11117;
  assign n15081 = n11011 & n11118;
  assign n15082 = (n11118 & n15023) | (n11118 & n15081) | (n15023 & n15081);
  assign n15083 = n11011 | n11118;
  assign n15084 = n15023 | n15083;
  assign n11121 = ~n15082 & n15084;
  assign n11122 = x70 & x108;
  assign n11123 = n11121 & n11122;
  assign n11124 = n11121 | n11122;
  assign n11125 = ~n11123 & n11124;
  assign n15085 = n11018 & n11125;
  assign n15086 = (n11125 & n15027) | (n11125 & n15085) | (n15027 & n15085);
  assign n15087 = n11018 | n11125;
  assign n15088 = n15027 | n15087;
  assign n11128 = ~n15086 & n15088;
  assign n11129 = x69 & x109;
  assign n11130 = n11128 & n11129;
  assign n11131 = n11128 | n11129;
  assign n11132 = ~n11130 & n11131;
  assign n15089 = n11025 & n11132;
  assign n15090 = (n11132 & n15031) | (n11132 & n15089) | (n15031 & n15089);
  assign n15091 = n11025 | n11132;
  assign n15092 = n15031 | n15091;
  assign n11135 = ~n15090 & n15092;
  assign n11136 = x68 & x110;
  assign n11137 = n11135 & n11136;
  assign n11138 = n11135 | n11136;
  assign n11139 = ~n11137 & n11138;
  assign n15093 = n11032 & n11139;
  assign n15094 = (n11139 & n15035) | (n11139 & n15093) | (n15035 & n15093);
  assign n15095 = n11032 | n11139;
  assign n15096 = n15035 | n15095;
  assign n11142 = ~n15094 & n15096;
  assign n11143 = x67 & x111;
  assign n11144 = n11142 & n11143;
  assign n11145 = n11142 | n11143;
  assign n11146 = ~n11144 & n11145;
  assign n15097 = n11039 & n11146;
  assign n15098 = (n11146 & n15039) | (n11146 & n15097) | (n15039 & n15097);
  assign n15099 = n11039 | n11146;
  assign n15100 = n15039 | n15099;
  assign n11149 = ~n15098 & n15100;
  assign n11163 = x79 & x100;
  assign n15104 = n11062 | n15049;
  assign n17423 = (n10955 & n15049) | (n10955 & n15104) | (n15049 & n15104);
  assign n15106 = n11163 & n17423;
  assign n66447 = n11163 & n50080;
  assign n66448 = n11059 & n11163;
  assign n66449 = (n10950 & n66447) | (n10950 & n66448) | (n66447 & n66448);
  assign n66450 = n11163 & n50083;
  assign n66451 = n11163 & n17398;
  assign n66452 = (n17326 & n66450) | (n17326 & n66451) | (n66450 & n66451);
  assign n50091 = (n17386 & n66449) | (n17386 & n66452) | (n66449 & n66452);
  assign n17425 = (n11062 & n11163) | (n11062 & n50091) | (n11163 & n50091);
  assign n17426 = (n14989 & n15106) | (n14989 & n17425) | (n15106 & n17425);
  assign n17427 = (n14988 & n15106) | (n14988 & n17425) | (n15106 & n17425);
  assign n17428 = (n14907 & n17426) | (n14907 & n17427) | (n17426 & n17427);
  assign n15109 = n11163 | n17423;
  assign n66453 = n11163 | n50080;
  assign n66454 = n11059 | n11163;
  assign n66455 = (n10950 & n66453) | (n10950 & n66454) | (n66453 & n66454);
  assign n66456 = n11163 | n50083;
  assign n66457 = n11163 | n17398;
  assign n66458 = (n17326 & n66456) | (n17326 & n66457) | (n66456 & n66457);
  assign n50094 = (n17386 & n66455) | (n17386 & n66458) | (n66455 & n66458);
  assign n17430 = n11062 | n50094;
  assign n17431 = (n14989 & n15109) | (n14989 & n17430) | (n15109 & n17430);
  assign n17432 = (n14988 & n15109) | (n14988 & n17430) | (n15109 & n17430);
  assign n17433 = (n14907 & n17431) | (n14907 & n17432) | (n17431 & n17432);
  assign n11166 = ~n17428 & n17433;
  assign n15113 = n11067 & n11166;
  assign n17434 = (n11069 & n11166) | (n11069 & n15113) | (n11166 & n15113);
  assign n17435 = (n15043 & n15113) | (n15043 & n17434) | (n15113 & n17434);
  assign n17436 = (n15113 & n17394) | (n15113 & n17434) | (n17394 & n17434);
  assign n17437 = (n17378 & n17435) | (n17378 & n17436) | (n17435 & n17436);
  assign n15116 = n11067 | n11166;
  assign n17438 = n11069 | n15116;
  assign n17439 = (n15043 & n15116) | (n15043 & n17438) | (n15116 & n17438);
  assign n17440 = (n15116 & n17394) | (n15116 & n17438) | (n17394 & n17438);
  assign n17441 = (n17378 & n17439) | (n17378 & n17440) | (n17439 & n17440);
  assign n11169 = ~n17437 & n17441;
  assign n11170 = x78 & x101;
  assign n11171 = n11169 & n11170;
  assign n11172 = n11169 | n11170;
  assign n11173 = ~n11171 & n11172;
  assign n15118 = n11074 & n11173;
  assign n15119 = (n11173 & n17419) | (n11173 & n15118) | (n17419 & n15118);
  assign n15120 = n11074 | n11173;
  assign n15121 = n17419 | n15120;
  assign n11176 = ~n15119 & n15121;
  assign n11177 = x77 & x102;
  assign n11178 = n11176 & n11177;
  assign n11179 = n11176 | n11177;
  assign n11180 = ~n11178 & n11179;
  assign n15122 = n11081 & n11180;
  assign n15123 = (n11180 & n15062) | (n11180 & n15122) | (n15062 & n15122);
  assign n15124 = n11081 | n11180;
  assign n15125 = n15062 | n15124;
  assign n11183 = ~n15123 & n15125;
  assign n11184 = x76 & x103;
  assign n11185 = n11183 & n11184;
  assign n11186 = n11183 | n11184;
  assign n11187 = ~n11185 & n11186;
  assign n15126 = n11088 & n11187;
  assign n15127 = (n11187 & n15066) | (n11187 & n15126) | (n15066 & n15126);
  assign n15128 = n11088 | n11187;
  assign n15129 = n15066 | n15128;
  assign n11190 = ~n15127 & n15129;
  assign n11191 = x75 & x104;
  assign n11192 = n11190 & n11191;
  assign n11193 = n11190 | n11191;
  assign n11194 = ~n11192 & n11193;
  assign n15130 = n11095 & n11194;
  assign n15131 = (n11194 & n15070) | (n11194 & n15130) | (n15070 & n15130);
  assign n15132 = n11095 | n11194;
  assign n15133 = n15070 | n15132;
  assign n11197 = ~n15131 & n15133;
  assign n11198 = x74 & x105;
  assign n11199 = n11197 & n11198;
  assign n11200 = n11197 | n11198;
  assign n11201 = ~n11199 & n11200;
  assign n15134 = n11102 & n11201;
  assign n15135 = (n11201 & n15074) | (n11201 & n15134) | (n15074 & n15134);
  assign n15136 = n11102 | n11201;
  assign n15137 = n15074 | n15136;
  assign n11204 = ~n15135 & n15137;
  assign n11205 = x73 & x106;
  assign n11206 = n11204 & n11205;
  assign n11207 = n11204 | n11205;
  assign n11208 = ~n11206 & n11207;
  assign n15138 = n11109 & n11208;
  assign n15139 = (n11208 & n15078) | (n11208 & n15138) | (n15078 & n15138);
  assign n15140 = n11109 | n11208;
  assign n15141 = n15078 | n15140;
  assign n11211 = ~n15139 & n15141;
  assign n11212 = x72 & x107;
  assign n11213 = n11211 & n11212;
  assign n11214 = n11211 | n11212;
  assign n11215 = ~n11213 & n11214;
  assign n15142 = n11116 & n11215;
  assign n15143 = (n11215 & n15082) | (n11215 & n15142) | (n15082 & n15142);
  assign n15144 = n11116 | n11215;
  assign n15145 = n15082 | n15144;
  assign n11218 = ~n15143 & n15145;
  assign n11219 = x71 & x108;
  assign n11220 = n11218 & n11219;
  assign n11221 = n11218 | n11219;
  assign n11222 = ~n11220 & n11221;
  assign n15146 = n11123 & n11222;
  assign n15147 = (n11222 & n15086) | (n11222 & n15146) | (n15086 & n15146);
  assign n15148 = n11123 | n11222;
  assign n15149 = n15086 | n15148;
  assign n11225 = ~n15147 & n15149;
  assign n11226 = x70 & x109;
  assign n11227 = n11225 & n11226;
  assign n11228 = n11225 | n11226;
  assign n11229 = ~n11227 & n11228;
  assign n15150 = n11130 & n11229;
  assign n15151 = (n11229 & n15090) | (n11229 & n15150) | (n15090 & n15150);
  assign n15152 = n11130 | n11229;
  assign n15153 = n15090 | n15152;
  assign n11232 = ~n15151 & n15153;
  assign n11233 = x69 & x110;
  assign n11234 = n11232 & n11233;
  assign n11235 = n11232 | n11233;
  assign n11236 = ~n11234 & n11235;
  assign n15154 = n11137 & n11236;
  assign n15155 = (n11236 & n15094) | (n11236 & n15154) | (n15094 & n15154);
  assign n15156 = n11137 | n11236;
  assign n15157 = n15094 | n15156;
  assign n11239 = ~n15155 & n15157;
  assign n11240 = x68 & x111;
  assign n11241 = n11239 & n11240;
  assign n11242 = n11239 | n11240;
  assign n11243 = ~n11241 & n11242;
  assign n15158 = n11144 & n11243;
  assign n15159 = (n11243 & n15098) | (n11243 & n15158) | (n15098 & n15158);
  assign n15160 = n11144 | n11243;
  assign n15161 = n15098 | n15160;
  assign n11246 = ~n15159 & n15161;
  assign n11259 = x79 & x101;
  assign n15165 = n11259 & n17428;
  assign n15166 = (n11259 & n17437) | (n11259 & n15165) | (n17437 & n15165);
  assign n15167 = n11259 | n17428;
  assign n15168 = n17437 | n15167;
  assign n11262 = ~n15166 & n15168;
  assign n50095 = n11171 & n11262;
  assign n50096 = (n11173 & n11262) | (n11173 & n50095) | (n11262 & n50095);
  assign n17442 = n11074 | n11171;
  assign n17443 = (n11171 & n11173) | (n11171 & n17442) | (n11173 & n17442);
  assign n17445 = n11262 & n17443;
  assign n17446 = (n17419 & n50096) | (n17419 & n17445) | (n50096 & n17445);
  assign n50097 = n11171 | n11262;
  assign n50098 = n11173 | n50097;
  assign n17448 = n11262 | n17443;
  assign n17449 = (n17419 & n50098) | (n17419 & n17448) | (n50098 & n17448);
  assign n11265 = ~n17446 & n17449;
  assign n11266 = x78 & x102;
  assign n11267 = n11265 & n11266;
  assign n11268 = n11265 | n11266;
  assign n11269 = ~n11267 & n11268;
  assign n15169 = n11178 & n11269;
  assign n17450 = (n11269 & n15122) | (n11269 & n15169) | (n15122 & n15169);
  assign n17451 = (n11180 & n11269) | (n11180 & n15169) | (n11269 & n15169);
  assign n17452 = (n15062 & n17450) | (n15062 & n17451) | (n17450 & n17451);
  assign n15171 = n11178 | n11269;
  assign n17453 = n15122 | n15171;
  assign n17454 = n11180 | n15171;
  assign n17455 = (n15062 & n17453) | (n15062 & n17454) | (n17453 & n17454);
  assign n11272 = ~n17452 & n17455;
  assign n11273 = x77 & x103;
  assign n11274 = n11272 & n11273;
  assign n11275 = n11272 | n11273;
  assign n11276 = ~n11274 & n11275;
  assign n15173 = n11185 & n11276;
  assign n15174 = (n11276 & n15127) | (n11276 & n15173) | (n15127 & n15173);
  assign n15175 = n11185 | n11276;
  assign n15176 = n15127 | n15175;
  assign n11279 = ~n15174 & n15176;
  assign n11280 = x76 & x104;
  assign n11281 = n11279 & n11280;
  assign n11282 = n11279 | n11280;
  assign n11283 = ~n11281 & n11282;
  assign n15177 = n11192 & n11283;
  assign n15178 = (n11283 & n15131) | (n11283 & n15177) | (n15131 & n15177);
  assign n15179 = n11192 | n11283;
  assign n15180 = n15131 | n15179;
  assign n11286 = ~n15178 & n15180;
  assign n11287 = x75 & x105;
  assign n11288 = n11286 & n11287;
  assign n11289 = n11286 | n11287;
  assign n11290 = ~n11288 & n11289;
  assign n15181 = n11199 & n11290;
  assign n15182 = (n11290 & n15135) | (n11290 & n15181) | (n15135 & n15181);
  assign n15183 = n11199 | n11290;
  assign n15184 = n15135 | n15183;
  assign n11293 = ~n15182 & n15184;
  assign n11294 = x74 & x106;
  assign n11295 = n11293 & n11294;
  assign n11296 = n11293 | n11294;
  assign n11297 = ~n11295 & n11296;
  assign n15185 = n11206 & n11297;
  assign n15186 = (n11297 & n15139) | (n11297 & n15185) | (n15139 & n15185);
  assign n15187 = n11206 | n11297;
  assign n15188 = n15139 | n15187;
  assign n11300 = ~n15186 & n15188;
  assign n11301 = x73 & x107;
  assign n11302 = n11300 & n11301;
  assign n11303 = n11300 | n11301;
  assign n11304 = ~n11302 & n11303;
  assign n15189 = n11213 & n11304;
  assign n15190 = (n11304 & n15143) | (n11304 & n15189) | (n15143 & n15189);
  assign n15191 = n11213 | n11304;
  assign n15192 = n15143 | n15191;
  assign n11307 = ~n15190 & n15192;
  assign n11308 = x72 & x108;
  assign n11309 = n11307 & n11308;
  assign n11310 = n11307 | n11308;
  assign n11311 = ~n11309 & n11310;
  assign n15193 = n11220 & n11311;
  assign n15194 = (n11311 & n15147) | (n11311 & n15193) | (n15147 & n15193);
  assign n15195 = n11220 | n11311;
  assign n15196 = n15147 | n15195;
  assign n11314 = ~n15194 & n15196;
  assign n11315 = x71 & x109;
  assign n11316 = n11314 & n11315;
  assign n11317 = n11314 | n11315;
  assign n11318 = ~n11316 & n11317;
  assign n15197 = n11227 & n11318;
  assign n15198 = (n11318 & n15151) | (n11318 & n15197) | (n15151 & n15197);
  assign n15199 = n11227 | n11318;
  assign n15200 = n15151 | n15199;
  assign n11321 = ~n15198 & n15200;
  assign n11322 = x70 & x110;
  assign n11323 = n11321 & n11322;
  assign n11324 = n11321 | n11322;
  assign n11325 = ~n11323 & n11324;
  assign n15201 = n11234 & n11325;
  assign n15202 = (n11325 & n15155) | (n11325 & n15201) | (n15155 & n15201);
  assign n15203 = n11234 | n11325;
  assign n15204 = n15155 | n15203;
  assign n11328 = ~n15202 & n15204;
  assign n11329 = x69 & x111;
  assign n11330 = n11328 & n11329;
  assign n11331 = n11328 | n11329;
  assign n11332 = ~n11330 & n11331;
  assign n15205 = n11241 & n11332;
  assign n15206 = (n11332 & n15159) | (n11332 & n15205) | (n15159 & n15205);
  assign n15207 = n11241 | n11332;
  assign n15208 = n15159 | n15207;
  assign n11335 = ~n15206 & n15208;
  assign n15163 = n11171 | n11173;
  assign n11347 = x79 & x102;
  assign n17458 = n11259 & n11347;
  assign n50099 = n17428 & n17458;
  assign n17459 = (n17437 & n50099) | (n17437 & n17458) | (n50099 & n17458);
  assign n17456 = (n11262 & n11347) | (n11262 & n17459) | (n11347 & n17459);
  assign n17460 = (n15163 & n17456) | (n15163 & n17459) | (n17456 & n17459);
  assign n17461 = (n17443 & n17456) | (n17443 & n17459) | (n17456 & n17459);
  assign n17462 = (n17419 & n17460) | (n17419 & n17461) | (n17460 & n17461);
  assign n17465 = n11259 | n11347;
  assign n50100 = (n11347 & n17428) | (n11347 & n17465) | (n17428 & n17465);
  assign n17466 = (n17437 & n50100) | (n17437 & n17465) | (n50100 & n17465);
  assign n17463 = n11262 | n17466;
  assign n17467 = (n15163 & n17463) | (n15163 & n17466) | (n17463 & n17466);
  assign n17468 = (n17443 & n17463) | (n17443 & n17466) | (n17463 & n17466);
  assign n17469 = (n17419 & n17467) | (n17419 & n17468) | (n17467 & n17468);
  assign n11350 = ~n17462 & n17469;
  assign n15217 = n11267 & n11350;
  assign n15218 = (n11350 & n17452) | (n11350 & n15217) | (n17452 & n15217);
  assign n15219 = n11267 | n11350;
  assign n15220 = n17452 | n15219;
  assign n11353 = ~n15218 & n15220;
  assign n11354 = x78 & x103;
  assign n11355 = n11353 & n11354;
  assign n11356 = n11353 | n11354;
  assign n11357 = ~n11355 & n11356;
  assign n15221 = n11274 & n11357;
  assign n15222 = (n11357 & n15174) | (n11357 & n15221) | (n15174 & n15221);
  assign n15223 = n11274 | n11357;
  assign n15224 = n15174 | n15223;
  assign n11360 = ~n15222 & n15224;
  assign n11361 = x77 & x104;
  assign n11362 = n11360 & n11361;
  assign n11363 = n11360 | n11361;
  assign n11364 = ~n11362 & n11363;
  assign n15225 = n11281 & n11364;
  assign n15226 = (n11364 & n15178) | (n11364 & n15225) | (n15178 & n15225);
  assign n15227 = n11281 | n11364;
  assign n15228 = n15178 | n15227;
  assign n11367 = ~n15226 & n15228;
  assign n11368 = x76 & x105;
  assign n11369 = n11367 & n11368;
  assign n11370 = n11367 | n11368;
  assign n11371 = ~n11369 & n11370;
  assign n15229 = n11288 & n11371;
  assign n15230 = (n11371 & n15182) | (n11371 & n15229) | (n15182 & n15229);
  assign n15231 = n11288 | n11371;
  assign n15232 = n15182 | n15231;
  assign n11374 = ~n15230 & n15232;
  assign n11375 = x75 & x106;
  assign n11376 = n11374 & n11375;
  assign n11377 = n11374 | n11375;
  assign n11378 = ~n11376 & n11377;
  assign n15233 = n11295 & n11378;
  assign n15234 = (n11378 & n15186) | (n11378 & n15233) | (n15186 & n15233);
  assign n15235 = n11295 | n11378;
  assign n15236 = n15186 | n15235;
  assign n11381 = ~n15234 & n15236;
  assign n11382 = x74 & x107;
  assign n11383 = n11381 & n11382;
  assign n11384 = n11381 | n11382;
  assign n11385 = ~n11383 & n11384;
  assign n15237 = n11302 & n11385;
  assign n15238 = (n11385 & n15190) | (n11385 & n15237) | (n15190 & n15237);
  assign n15239 = n11302 | n11385;
  assign n15240 = n15190 | n15239;
  assign n11388 = ~n15238 & n15240;
  assign n11389 = x73 & x108;
  assign n11390 = n11388 & n11389;
  assign n11391 = n11388 | n11389;
  assign n11392 = ~n11390 & n11391;
  assign n15241 = n11309 & n11392;
  assign n15242 = (n11392 & n15194) | (n11392 & n15241) | (n15194 & n15241);
  assign n15243 = n11309 | n11392;
  assign n15244 = n15194 | n15243;
  assign n11395 = ~n15242 & n15244;
  assign n11396 = x72 & x109;
  assign n11397 = n11395 & n11396;
  assign n11398 = n11395 | n11396;
  assign n11399 = ~n11397 & n11398;
  assign n15245 = n11316 & n11399;
  assign n15246 = (n11399 & n15198) | (n11399 & n15245) | (n15198 & n15245);
  assign n15247 = n11316 | n11399;
  assign n15248 = n15198 | n15247;
  assign n11402 = ~n15246 & n15248;
  assign n11403 = x71 & x110;
  assign n11404 = n11402 & n11403;
  assign n11405 = n11402 | n11403;
  assign n11406 = ~n11404 & n11405;
  assign n15249 = n11323 & n11406;
  assign n15250 = (n11406 & n15202) | (n11406 & n15249) | (n15202 & n15249);
  assign n15251 = n11323 | n11406;
  assign n15252 = n15202 | n15251;
  assign n11409 = ~n15250 & n15252;
  assign n11410 = x70 & x111;
  assign n11411 = n11409 & n11410;
  assign n11412 = n11409 | n11410;
  assign n11413 = ~n11411 & n11412;
  assign n15253 = n11330 & n11413;
  assign n15254 = (n11413 & n15206) | (n11413 & n15253) | (n15206 & n15253);
  assign n15255 = n11330 | n11413;
  assign n15256 = n15206 | n15255;
  assign n11416 = ~n15254 & n15256;
  assign n11427 = x79 & x103;
  assign n17470 = n11350 | n17462;
  assign n17471 = (n11267 & n17462) | (n11267 & n17470) | (n17462 & n17470);
  assign n15260 = n11427 & n17471;
  assign n66459 = n11427 & n17456;
  assign n66460 = n11427 & n17459;
  assign n66461 = (n17443 & n66459) | (n17443 & n66460) | (n66459 & n66460);
  assign n66462 = (n15163 & n66459) | (n15163 & n66460) | (n66459 & n66460);
  assign n50103 = (n17419 & n66461) | (n17419 & n66462) | (n66461 & n66462);
  assign n17473 = (n11350 & n11427) | (n11350 & n50103) | (n11427 & n50103);
  assign n15262 = (n17452 & n15260) | (n17452 & n17473) | (n15260 & n17473);
  assign n15263 = n11427 | n17471;
  assign n66463 = n11427 | n17456;
  assign n66464 = n11427 | n17459;
  assign n66465 = (n17443 & n66463) | (n17443 & n66464) | (n66463 & n66464);
  assign n66466 = (n15163 & n66463) | (n15163 & n66464) | (n66463 & n66464);
  assign n50106 = (n17419 & n66465) | (n17419 & n66466) | (n66465 & n66466);
  assign n17475 = n11350 | n50106;
  assign n15265 = (n17452 & n15263) | (n17452 & n17475) | (n15263 & n17475);
  assign n11430 = ~n15262 & n15265;
  assign n15266 = n11355 & n11430;
  assign n17476 = (n11430 & n15221) | (n11430 & n15266) | (n15221 & n15266);
  assign n17477 = (n11357 & n11430) | (n11357 & n15266) | (n11430 & n15266);
  assign n17478 = (n15174 & n17476) | (n15174 & n17477) | (n17476 & n17477);
  assign n15268 = n11355 | n11430;
  assign n17479 = n15221 | n15268;
  assign n17480 = n11357 | n15268;
  assign n17481 = (n15174 & n17479) | (n15174 & n17480) | (n17479 & n17480);
  assign n11433 = ~n17478 & n17481;
  assign n11434 = x78 & x104;
  assign n11435 = n11433 & n11434;
  assign n11436 = n11433 | n11434;
  assign n11437 = ~n11435 & n11436;
  assign n15270 = n11362 & n11437;
  assign n15271 = (n11437 & n15226) | (n11437 & n15270) | (n15226 & n15270);
  assign n15272 = n11362 | n11437;
  assign n15273 = n15226 | n15272;
  assign n11440 = ~n15271 & n15273;
  assign n11441 = x77 & x105;
  assign n11442 = n11440 & n11441;
  assign n11443 = n11440 | n11441;
  assign n11444 = ~n11442 & n11443;
  assign n15274 = n11369 & n11444;
  assign n15275 = (n11444 & n15230) | (n11444 & n15274) | (n15230 & n15274);
  assign n15276 = n11369 | n11444;
  assign n15277 = n15230 | n15276;
  assign n11447 = ~n15275 & n15277;
  assign n11448 = x76 & x106;
  assign n11449 = n11447 & n11448;
  assign n11450 = n11447 | n11448;
  assign n11451 = ~n11449 & n11450;
  assign n15278 = n11376 & n11451;
  assign n15279 = (n11451 & n15234) | (n11451 & n15278) | (n15234 & n15278);
  assign n15280 = n11376 | n11451;
  assign n15281 = n15234 | n15280;
  assign n11454 = ~n15279 & n15281;
  assign n11455 = x75 & x107;
  assign n11456 = n11454 & n11455;
  assign n11457 = n11454 | n11455;
  assign n11458 = ~n11456 & n11457;
  assign n15282 = n11383 & n11458;
  assign n15283 = (n11458 & n15238) | (n11458 & n15282) | (n15238 & n15282);
  assign n15284 = n11383 | n11458;
  assign n15285 = n15238 | n15284;
  assign n11461 = ~n15283 & n15285;
  assign n11462 = x74 & x108;
  assign n11463 = n11461 & n11462;
  assign n11464 = n11461 | n11462;
  assign n11465 = ~n11463 & n11464;
  assign n15286 = n11390 & n11465;
  assign n15287 = (n11465 & n15242) | (n11465 & n15286) | (n15242 & n15286);
  assign n15288 = n11390 | n11465;
  assign n15289 = n15242 | n15288;
  assign n11468 = ~n15287 & n15289;
  assign n11469 = x73 & x109;
  assign n11470 = n11468 & n11469;
  assign n11471 = n11468 | n11469;
  assign n11472 = ~n11470 & n11471;
  assign n15290 = n11397 & n11472;
  assign n15291 = (n11472 & n15246) | (n11472 & n15290) | (n15246 & n15290);
  assign n15292 = n11397 | n11472;
  assign n15293 = n15246 | n15292;
  assign n11475 = ~n15291 & n15293;
  assign n11476 = x72 & x110;
  assign n11477 = n11475 & n11476;
  assign n11478 = n11475 | n11476;
  assign n11479 = ~n11477 & n11478;
  assign n15294 = n11404 & n11479;
  assign n15295 = (n11479 & n15250) | (n11479 & n15294) | (n15250 & n15294);
  assign n15296 = n11404 | n11479;
  assign n15297 = n15250 | n15296;
  assign n11482 = ~n15295 & n15297;
  assign n11483 = x71 & x111;
  assign n11484 = n11482 & n11483;
  assign n11485 = n11482 | n11483;
  assign n11486 = ~n11484 & n11485;
  assign n15298 = n11411 & n11486;
  assign n15299 = (n11486 & n15254) | (n11486 & n15298) | (n15254 & n15298);
  assign n15300 = n11411 | n11486;
  assign n15301 = n15254 | n15300;
  assign n11489 = ~n15299 & n15301;
  assign n11499 = x79 & x104;
  assign n15303 = n11430 | n15262;
  assign n17482 = (n11355 & n15262) | (n11355 & n15303) | (n15262 & n15303);
  assign n15305 = n11499 & n17482;
  assign n66467 = n11427 & n11499;
  assign n66468 = n17471 & n66467;
  assign n66469 = n11499 & n50103;
  assign n66470 = (n11350 & n66467) | (n11350 & n66469) | (n66467 & n66469);
  assign n50109 = (n17452 & n66468) | (n17452 & n66470) | (n66468 & n66470);
  assign n17484 = (n11430 & n11499) | (n11430 & n50109) | (n11499 & n50109);
  assign n17485 = (n15221 & n15305) | (n15221 & n17484) | (n15305 & n17484);
  assign n17486 = (n11357 & n15305) | (n11357 & n17484) | (n15305 & n17484);
  assign n17487 = (n15174 & n17485) | (n15174 & n17486) | (n17485 & n17486);
  assign n15308 = n11499 | n17482;
  assign n66471 = n11427 | n11499;
  assign n66472 = (n11499 & n17471) | (n11499 & n66471) | (n17471 & n66471);
  assign n66473 = n11499 | n50103;
  assign n66474 = (n11350 & n66471) | (n11350 & n66473) | (n66471 & n66473);
  assign n50112 = (n17452 & n66472) | (n17452 & n66474) | (n66472 & n66474);
  assign n17489 = n11430 | n50112;
  assign n17490 = (n15221 & n15308) | (n15221 & n17489) | (n15308 & n17489);
  assign n17491 = (n11357 & n15308) | (n11357 & n17489) | (n15308 & n17489);
  assign n17492 = (n15174 & n17490) | (n15174 & n17491) | (n17490 & n17491);
  assign n11502 = ~n17487 & n17492;
  assign n15311 = n11435 & n11502;
  assign n17493 = (n11502 & n15270) | (n11502 & n15311) | (n15270 & n15311);
  assign n17494 = (n11437 & n11502) | (n11437 & n15311) | (n11502 & n15311);
  assign n17495 = (n15226 & n17493) | (n15226 & n17494) | (n17493 & n17494);
  assign n15313 = n11435 | n11502;
  assign n17496 = n15270 | n15313;
  assign n17497 = n11437 | n15313;
  assign n17498 = (n15226 & n17496) | (n15226 & n17497) | (n17496 & n17497);
  assign n11505 = ~n17495 & n17498;
  assign n11506 = x78 & x105;
  assign n11507 = n11505 & n11506;
  assign n11508 = n11505 | n11506;
  assign n11509 = ~n11507 & n11508;
  assign n15315 = n11442 & n11509;
  assign n15316 = (n11509 & n15275) | (n11509 & n15315) | (n15275 & n15315);
  assign n15317 = n11442 | n11509;
  assign n15318 = n15275 | n15317;
  assign n11512 = ~n15316 & n15318;
  assign n11513 = x77 & x106;
  assign n11514 = n11512 & n11513;
  assign n11515 = n11512 | n11513;
  assign n11516 = ~n11514 & n11515;
  assign n15319 = n11449 & n11516;
  assign n15320 = (n11516 & n15279) | (n11516 & n15319) | (n15279 & n15319);
  assign n15321 = n11449 | n11516;
  assign n15322 = n15279 | n15321;
  assign n11519 = ~n15320 & n15322;
  assign n11520 = x76 & x107;
  assign n11521 = n11519 & n11520;
  assign n11522 = n11519 | n11520;
  assign n11523 = ~n11521 & n11522;
  assign n15323 = n11456 & n11523;
  assign n15324 = (n11523 & n15283) | (n11523 & n15323) | (n15283 & n15323);
  assign n15325 = n11456 | n11523;
  assign n15326 = n15283 | n15325;
  assign n11526 = ~n15324 & n15326;
  assign n11527 = x75 & x108;
  assign n11528 = n11526 & n11527;
  assign n11529 = n11526 | n11527;
  assign n11530 = ~n11528 & n11529;
  assign n15327 = n11463 & n11530;
  assign n15328 = (n11530 & n15287) | (n11530 & n15327) | (n15287 & n15327);
  assign n15329 = n11463 | n11530;
  assign n15330 = n15287 | n15329;
  assign n11533 = ~n15328 & n15330;
  assign n11534 = x74 & x109;
  assign n11535 = n11533 & n11534;
  assign n11536 = n11533 | n11534;
  assign n11537 = ~n11535 & n11536;
  assign n15331 = n11470 & n11537;
  assign n15332 = (n11537 & n15291) | (n11537 & n15331) | (n15291 & n15331);
  assign n15333 = n11470 | n11537;
  assign n15334 = n15291 | n15333;
  assign n11540 = ~n15332 & n15334;
  assign n11541 = x73 & x110;
  assign n11542 = n11540 & n11541;
  assign n11543 = n11540 | n11541;
  assign n11544 = ~n11542 & n11543;
  assign n15335 = n11477 & n11544;
  assign n15336 = (n11544 & n15295) | (n11544 & n15335) | (n15295 & n15335);
  assign n15337 = n11477 | n11544;
  assign n15338 = n15295 | n15337;
  assign n11547 = ~n15336 & n15338;
  assign n11548 = x72 & x111;
  assign n11549 = n11547 & n11548;
  assign n11550 = n11547 | n11548;
  assign n11551 = ~n11549 & n11550;
  assign n15339 = n11484 & n11551;
  assign n15340 = (n11551 & n15299) | (n11551 & n15339) | (n15299 & n15339);
  assign n15341 = n11484 | n11551;
  assign n15342 = n15299 | n15341;
  assign n11554 = ~n15340 & n15342;
  assign n11563 = x79 & x105;
  assign n17499 = n11502 | n17487;
  assign n17500 = (n11435 & n17487) | (n11435 & n17499) | (n17487 & n17499);
  assign n15346 = n11563 & n17500;
  assign n17501 = n11563 & n17487;
  assign n17502 = (n11502 & n11563) | (n11502 & n17501) | (n11563 & n17501);
  assign n17503 = (n15270 & n15346) | (n15270 & n17502) | (n15346 & n17502);
  assign n17504 = (n11437 & n15346) | (n11437 & n17502) | (n15346 & n17502);
  assign n17505 = (n15226 & n17503) | (n15226 & n17504) | (n17503 & n17504);
  assign n15349 = n11563 | n17500;
  assign n17506 = n11563 | n17487;
  assign n17507 = n11502 | n17506;
  assign n17508 = (n15270 & n15349) | (n15270 & n17507) | (n15349 & n17507);
  assign n17509 = (n11437 & n15349) | (n11437 & n17507) | (n15349 & n17507);
  assign n17510 = (n15226 & n17508) | (n15226 & n17509) | (n17508 & n17509);
  assign n11566 = ~n17505 & n17510;
  assign n15352 = n11507 & n11566;
  assign n17511 = (n11566 & n15315) | (n11566 & n15352) | (n15315 & n15352);
  assign n17512 = (n11509 & n11566) | (n11509 & n15352) | (n11566 & n15352);
  assign n17513 = (n15275 & n17511) | (n15275 & n17512) | (n17511 & n17512);
  assign n15354 = n11507 | n11566;
  assign n17514 = n15315 | n15354;
  assign n17515 = n11509 | n15354;
  assign n17516 = (n15275 & n17514) | (n15275 & n17515) | (n17514 & n17515);
  assign n11569 = ~n17513 & n17516;
  assign n11570 = x78 & x106;
  assign n11571 = n11569 & n11570;
  assign n11572 = n11569 | n11570;
  assign n11573 = ~n11571 & n11572;
  assign n15356 = n11514 & n11573;
  assign n15357 = (n11573 & n15320) | (n11573 & n15356) | (n15320 & n15356);
  assign n15358 = n11514 | n11573;
  assign n15359 = n15320 | n15358;
  assign n11576 = ~n15357 & n15359;
  assign n11577 = x77 & x107;
  assign n11578 = n11576 & n11577;
  assign n11579 = n11576 | n11577;
  assign n11580 = ~n11578 & n11579;
  assign n15360 = n11521 & n11580;
  assign n15361 = (n11580 & n15324) | (n11580 & n15360) | (n15324 & n15360);
  assign n15362 = n11521 | n11580;
  assign n15363 = n15324 | n15362;
  assign n11583 = ~n15361 & n15363;
  assign n11584 = x76 & x108;
  assign n11585 = n11583 & n11584;
  assign n11586 = n11583 | n11584;
  assign n11587 = ~n11585 & n11586;
  assign n15364 = n11528 & n11587;
  assign n15365 = (n11587 & n15328) | (n11587 & n15364) | (n15328 & n15364);
  assign n15366 = n11528 | n11587;
  assign n15367 = n15328 | n15366;
  assign n11590 = ~n15365 & n15367;
  assign n11591 = x75 & x109;
  assign n11592 = n11590 & n11591;
  assign n11593 = n11590 | n11591;
  assign n11594 = ~n11592 & n11593;
  assign n15368 = n11535 & n11594;
  assign n15369 = (n11594 & n15332) | (n11594 & n15368) | (n15332 & n15368);
  assign n15370 = n11535 | n11594;
  assign n15371 = n15332 | n15370;
  assign n11597 = ~n15369 & n15371;
  assign n11598 = x74 & x110;
  assign n11599 = n11597 & n11598;
  assign n11600 = n11597 | n11598;
  assign n11601 = ~n11599 & n11600;
  assign n15372 = n11542 & n11601;
  assign n15373 = (n11601 & n15336) | (n11601 & n15372) | (n15336 & n15372);
  assign n15374 = n11542 | n11601;
  assign n15375 = n15336 | n15374;
  assign n11604 = ~n15373 & n15375;
  assign n11605 = x73 & x111;
  assign n11606 = n11604 & n11605;
  assign n11607 = n11604 | n11605;
  assign n11608 = ~n11606 & n11607;
  assign n15376 = n11549 & n11608;
  assign n15377 = (n11608 & n15340) | (n11608 & n15376) | (n15340 & n15376);
  assign n15378 = n11549 | n11608;
  assign n15379 = n15340 | n15378;
  assign n11611 = ~n15377 & n15379;
  assign n11619 = x79 & x106;
  assign n17517 = n11566 | n17505;
  assign n17518 = (n11507 & n17505) | (n11507 & n17517) | (n17505 & n17517);
  assign n15383 = n11619 & n17518;
  assign n17519 = n11619 & n17505;
  assign n17520 = (n11566 & n11619) | (n11566 & n17519) | (n11619 & n17519);
  assign n17521 = (n15315 & n15383) | (n15315 & n17520) | (n15383 & n17520);
  assign n17522 = (n11509 & n15383) | (n11509 & n17520) | (n15383 & n17520);
  assign n17523 = (n15275 & n17521) | (n15275 & n17522) | (n17521 & n17522);
  assign n15386 = n11619 | n17518;
  assign n17524 = n11619 | n17505;
  assign n17525 = n11566 | n17524;
  assign n17526 = (n15315 & n15386) | (n15315 & n17525) | (n15386 & n17525);
  assign n17527 = (n11509 & n15386) | (n11509 & n17525) | (n15386 & n17525);
  assign n17528 = (n15275 & n17526) | (n15275 & n17527) | (n17526 & n17527);
  assign n11622 = ~n17523 & n17528;
  assign n15389 = n11571 & n11622;
  assign n17529 = (n11622 & n15356) | (n11622 & n15389) | (n15356 & n15389);
  assign n17530 = (n11573 & n11622) | (n11573 & n15389) | (n11622 & n15389);
  assign n17531 = (n15320 & n17529) | (n15320 & n17530) | (n17529 & n17530);
  assign n15391 = n11571 | n11622;
  assign n17532 = n15356 | n15391;
  assign n17533 = n11573 | n15391;
  assign n17534 = (n15320 & n17532) | (n15320 & n17533) | (n17532 & n17533);
  assign n11625 = ~n17531 & n17534;
  assign n11626 = x78 & x107;
  assign n11627 = n11625 & n11626;
  assign n11628 = n11625 | n11626;
  assign n11629 = ~n11627 & n11628;
  assign n15393 = n11578 & n11629;
  assign n15394 = (n11629 & n15361) | (n11629 & n15393) | (n15361 & n15393);
  assign n15395 = n11578 | n11629;
  assign n15396 = n15361 | n15395;
  assign n11632 = ~n15394 & n15396;
  assign n11633 = x77 & x108;
  assign n11634 = n11632 & n11633;
  assign n11635 = n11632 | n11633;
  assign n11636 = ~n11634 & n11635;
  assign n15397 = n11585 & n11636;
  assign n15398 = (n11636 & n15365) | (n11636 & n15397) | (n15365 & n15397);
  assign n15399 = n11585 | n11636;
  assign n15400 = n15365 | n15399;
  assign n11639 = ~n15398 & n15400;
  assign n11640 = x76 & x109;
  assign n11641 = n11639 & n11640;
  assign n11642 = n11639 | n11640;
  assign n11643 = ~n11641 & n11642;
  assign n15401 = n11592 & n11643;
  assign n15402 = (n11643 & n15369) | (n11643 & n15401) | (n15369 & n15401);
  assign n15403 = n11592 | n11643;
  assign n15404 = n15369 | n15403;
  assign n11646 = ~n15402 & n15404;
  assign n11647 = x75 & x110;
  assign n11648 = n11646 & n11647;
  assign n11649 = n11646 | n11647;
  assign n11650 = ~n11648 & n11649;
  assign n15405 = n11599 & n11650;
  assign n15406 = (n11650 & n15373) | (n11650 & n15405) | (n15373 & n15405);
  assign n15407 = n11599 | n11650;
  assign n15408 = n15373 | n15407;
  assign n11653 = ~n15406 & n15408;
  assign n11654 = x74 & x111;
  assign n11655 = n11653 & n11654;
  assign n11656 = n11653 | n11654;
  assign n11657 = ~n11655 & n11656;
  assign n15409 = n11606 & n11657;
  assign n15410 = (n11657 & n15377) | (n11657 & n15409) | (n15377 & n15409);
  assign n15411 = n11606 | n11657;
  assign n15412 = n15377 | n15411;
  assign n11660 = ~n15410 & n15412;
  assign n11667 = x79 & x107;
  assign n17535 = n11622 | n17523;
  assign n17536 = (n11571 & n17523) | (n11571 & n17535) | (n17523 & n17535);
  assign n15416 = n11667 & n17536;
  assign n17537 = n11667 & n17523;
  assign n17538 = (n11622 & n11667) | (n11622 & n17537) | (n11667 & n17537);
  assign n17539 = (n15356 & n15416) | (n15356 & n17538) | (n15416 & n17538);
  assign n17540 = (n11573 & n15416) | (n11573 & n17538) | (n15416 & n17538);
  assign n17541 = (n15320 & n17539) | (n15320 & n17540) | (n17539 & n17540);
  assign n15419 = n11667 | n17536;
  assign n17542 = n11667 | n17523;
  assign n17543 = n11622 | n17542;
  assign n17544 = (n15356 & n15419) | (n15356 & n17543) | (n15419 & n17543);
  assign n17545 = (n11573 & n15419) | (n11573 & n17543) | (n15419 & n17543);
  assign n17546 = (n15320 & n17544) | (n15320 & n17545) | (n17544 & n17545);
  assign n11670 = ~n17541 & n17546;
  assign n15422 = n11627 & n11670;
  assign n17547 = (n11670 & n15393) | (n11670 & n15422) | (n15393 & n15422);
  assign n17548 = (n11629 & n11670) | (n11629 & n15422) | (n11670 & n15422);
  assign n17549 = (n15361 & n17547) | (n15361 & n17548) | (n17547 & n17548);
  assign n15424 = n11627 | n11670;
  assign n17550 = n15393 | n15424;
  assign n17551 = n11629 | n15424;
  assign n17552 = (n15361 & n17550) | (n15361 & n17551) | (n17550 & n17551);
  assign n11673 = ~n17549 & n17552;
  assign n11674 = x78 & x108;
  assign n11675 = n11673 & n11674;
  assign n11676 = n11673 | n11674;
  assign n11677 = ~n11675 & n11676;
  assign n15426 = n11634 & n11677;
  assign n15427 = (n11677 & n15398) | (n11677 & n15426) | (n15398 & n15426);
  assign n15428 = n11634 | n11677;
  assign n15429 = n15398 | n15428;
  assign n11680 = ~n15427 & n15429;
  assign n11681 = x77 & x109;
  assign n11682 = n11680 & n11681;
  assign n11683 = n11680 | n11681;
  assign n11684 = ~n11682 & n11683;
  assign n15430 = n11641 & n11684;
  assign n15431 = (n11684 & n15402) | (n11684 & n15430) | (n15402 & n15430);
  assign n15432 = n11641 | n11684;
  assign n15433 = n15402 | n15432;
  assign n11687 = ~n15431 & n15433;
  assign n11688 = x76 & x110;
  assign n11689 = n11687 & n11688;
  assign n11690 = n11687 | n11688;
  assign n11691 = ~n11689 & n11690;
  assign n15434 = n11648 & n11691;
  assign n15435 = (n11691 & n15406) | (n11691 & n15434) | (n15406 & n15434);
  assign n15436 = n11648 | n11691;
  assign n15437 = n15406 | n15436;
  assign n11694 = ~n15435 & n15437;
  assign n11695 = x75 & x111;
  assign n11696 = n11694 & n11695;
  assign n11697 = n11694 | n11695;
  assign n11698 = ~n11696 & n11697;
  assign n15438 = n11655 & n11698;
  assign n15439 = (n11698 & n15410) | (n11698 & n15438) | (n15410 & n15438);
  assign n15440 = n11655 | n11698;
  assign n15441 = n15410 | n15440;
  assign n11701 = ~n15439 & n15441;
  assign n11707 = x79 & x108;
  assign n17553 = n11670 | n17541;
  assign n17554 = (n11627 & n17541) | (n11627 & n17553) | (n17541 & n17553);
  assign n15445 = n11707 & n17554;
  assign n17555 = n11707 & n17541;
  assign n17556 = (n11670 & n11707) | (n11670 & n17555) | (n11707 & n17555);
  assign n17557 = (n15393 & n15445) | (n15393 & n17556) | (n15445 & n17556);
  assign n17558 = (n11629 & n15445) | (n11629 & n17556) | (n15445 & n17556);
  assign n17559 = (n15361 & n17557) | (n15361 & n17558) | (n17557 & n17558);
  assign n15448 = n11707 | n17554;
  assign n17560 = n11707 | n17541;
  assign n17561 = n11670 | n17560;
  assign n17562 = (n15393 & n15448) | (n15393 & n17561) | (n15448 & n17561);
  assign n17563 = (n11629 & n15448) | (n11629 & n17561) | (n15448 & n17561);
  assign n17564 = (n15361 & n17562) | (n15361 & n17563) | (n17562 & n17563);
  assign n11710 = ~n17559 & n17564;
  assign n15451 = n11675 & n11710;
  assign n17565 = (n11710 & n15426) | (n11710 & n15451) | (n15426 & n15451);
  assign n17566 = (n11677 & n11710) | (n11677 & n15451) | (n11710 & n15451);
  assign n17567 = (n15398 & n17565) | (n15398 & n17566) | (n17565 & n17566);
  assign n15453 = n11675 | n11710;
  assign n17568 = n15426 | n15453;
  assign n17569 = n11677 | n15453;
  assign n17570 = (n15398 & n17568) | (n15398 & n17569) | (n17568 & n17569);
  assign n11713 = ~n17567 & n17570;
  assign n11714 = x78 & x109;
  assign n11715 = n11713 & n11714;
  assign n11716 = n11713 | n11714;
  assign n11717 = ~n11715 & n11716;
  assign n15455 = n11682 & n11717;
  assign n15456 = (n11717 & n15431) | (n11717 & n15455) | (n15431 & n15455);
  assign n15457 = n11682 | n11717;
  assign n15458 = n15431 | n15457;
  assign n11720 = ~n15456 & n15458;
  assign n11721 = x77 & x110;
  assign n11722 = n11720 & n11721;
  assign n11723 = n11720 | n11721;
  assign n11724 = ~n11722 & n11723;
  assign n15459 = n11689 & n11724;
  assign n15460 = (n11724 & n15435) | (n11724 & n15459) | (n15435 & n15459);
  assign n15461 = n11689 | n11724;
  assign n15462 = n15435 | n15461;
  assign n11727 = ~n15460 & n15462;
  assign n11728 = x76 & x111;
  assign n11729 = n11727 & n11728;
  assign n11730 = n11727 | n11728;
  assign n11731 = ~n11729 & n11730;
  assign n15463 = n11696 & n11731;
  assign n15464 = (n11731 & n15439) | (n11731 & n15463) | (n15439 & n15463);
  assign n15465 = n11696 | n11731;
  assign n15466 = n15439 | n15465;
  assign n11734 = ~n15464 & n15466;
  assign n11739 = x79 & x109;
  assign n17571 = n11710 | n17559;
  assign n17572 = (n11675 & n17559) | (n11675 & n17571) | (n17559 & n17571);
  assign n15470 = n11739 & n17572;
  assign n17573 = n11739 & n17559;
  assign n17574 = (n11710 & n11739) | (n11710 & n17573) | (n11739 & n17573);
  assign n17575 = (n15426 & n15470) | (n15426 & n17574) | (n15470 & n17574);
  assign n17576 = (n11677 & n15470) | (n11677 & n17574) | (n15470 & n17574);
  assign n17577 = (n15398 & n17575) | (n15398 & n17576) | (n17575 & n17576);
  assign n15473 = n11739 | n17572;
  assign n17578 = n11739 | n17559;
  assign n17579 = n11710 | n17578;
  assign n17580 = (n15426 & n15473) | (n15426 & n17579) | (n15473 & n17579);
  assign n17581 = (n11677 & n15473) | (n11677 & n17579) | (n15473 & n17579);
  assign n17582 = (n15398 & n17580) | (n15398 & n17581) | (n17580 & n17581);
  assign n11742 = ~n17577 & n17582;
  assign n15476 = n11715 & n11742;
  assign n17583 = (n11742 & n15455) | (n11742 & n15476) | (n15455 & n15476);
  assign n17584 = (n11717 & n11742) | (n11717 & n15476) | (n11742 & n15476);
  assign n17585 = (n15431 & n17583) | (n15431 & n17584) | (n17583 & n17584);
  assign n15478 = n11715 | n11742;
  assign n17586 = n15455 | n15478;
  assign n17587 = n11717 | n15478;
  assign n17588 = (n15431 & n17586) | (n15431 & n17587) | (n17586 & n17587);
  assign n11745 = ~n17585 & n17588;
  assign n11746 = x78 & x110;
  assign n11747 = n11745 & n11746;
  assign n11748 = n11745 | n11746;
  assign n11749 = ~n11747 & n11748;
  assign n15480 = n11722 & n11749;
  assign n15481 = (n11749 & n15460) | (n11749 & n15480) | (n15460 & n15480);
  assign n15482 = n11722 | n11749;
  assign n15483 = n15460 | n15482;
  assign n11752 = ~n15481 & n15483;
  assign n11753 = x77 & x111;
  assign n11754 = n11752 & n11753;
  assign n11755 = n11752 | n11753;
  assign n11756 = ~n11754 & n11755;
  assign n15484 = n11729 & n11756;
  assign n15485 = (n11756 & n15464) | (n11756 & n15484) | (n15464 & n15484);
  assign n15486 = n11729 | n11756;
  assign n15487 = n15464 | n15486;
  assign n11759 = ~n15485 & n15487;
  assign n11763 = x79 & x110;
  assign n17589 = n11742 | n17577;
  assign n17590 = (n11715 & n17577) | (n11715 & n17589) | (n17577 & n17589);
  assign n15491 = n11763 & n17590;
  assign n17591 = n11763 & n17577;
  assign n17592 = (n11742 & n11763) | (n11742 & n17591) | (n11763 & n17591);
  assign n17593 = (n15455 & n15491) | (n15455 & n17592) | (n15491 & n17592);
  assign n17594 = (n11717 & n15491) | (n11717 & n17592) | (n15491 & n17592);
  assign n17595 = (n15431 & n17593) | (n15431 & n17594) | (n17593 & n17594);
  assign n15494 = n11763 | n17590;
  assign n17596 = n11763 | n17577;
  assign n17597 = n11742 | n17596;
  assign n17598 = (n15455 & n15494) | (n15455 & n17597) | (n15494 & n17597);
  assign n17599 = (n11717 & n15494) | (n11717 & n17597) | (n15494 & n17597);
  assign n17600 = (n15431 & n17598) | (n15431 & n17599) | (n17598 & n17599);
  assign n11766 = ~n17595 & n17600;
  assign n15497 = n11747 & n11766;
  assign n17601 = (n11766 & n15480) | (n11766 & n15497) | (n15480 & n15497);
  assign n17602 = (n11749 & n11766) | (n11749 & n15497) | (n11766 & n15497);
  assign n17603 = (n15460 & n17601) | (n15460 & n17602) | (n17601 & n17602);
  assign n15499 = n11747 | n11766;
  assign n17604 = n15480 | n15499;
  assign n17605 = n11749 | n15499;
  assign n17606 = (n15460 & n17604) | (n15460 & n17605) | (n17604 & n17605);
  assign n11769 = ~n17603 & n17606;
  assign n11770 = x78 & x111;
  assign n11771 = n11769 & n11770;
  assign n11772 = n11769 | n11770;
  assign n11773 = ~n11771 & n11772;
  assign n15501 = n11754 & n11773;
  assign n15502 = (n11773 & n15485) | (n11773 & n15501) | (n15485 & n15501);
  assign n15503 = n11754 | n11773;
  assign n15504 = n15485 | n15503;
  assign n11776 = ~n15502 & n15504;
  assign n11779 = x79 & x111;
  assign n17607 = n11766 | n17595;
  assign n17608 = (n11747 & n17595) | (n11747 & n17607) | (n17595 & n17607);
  assign n15508 = n11779 & n17608;
  assign n17609 = n11779 & n17595;
  assign n17610 = (n11766 & n11779) | (n11766 & n17609) | (n11779 & n17609);
  assign n17611 = (n15480 & n15508) | (n15480 & n17610) | (n15508 & n17610);
  assign n17612 = (n11749 & n15508) | (n11749 & n17610) | (n15508 & n17610);
  assign n17613 = (n15460 & n17611) | (n15460 & n17612) | (n17611 & n17612);
  assign n15511 = n11779 | n17608;
  assign n17614 = n11779 | n17595;
  assign n17615 = n11766 | n17614;
  assign n17616 = (n15480 & n15511) | (n15480 & n17615) | (n15511 & n17615);
  assign n17617 = (n11749 & n15511) | (n11749 & n17615) | (n15511 & n17615);
  assign n17618 = (n15460 & n17616) | (n15460 & n17617) | (n17616 & n17617);
  assign n11782 = ~n17613 & n17618;
  assign n15514 = n11771 & n11782;
  assign n17619 = (n11782 & n15501) | (n11782 & n15514) | (n15501 & n15514);
  assign n17620 = (n11773 & n11782) | (n11773 & n15514) | (n11782 & n15514);
  assign n17621 = (n15485 & n17619) | (n15485 & n17620) | (n17619 & n17620);
  assign n15516 = n11771 | n11782;
  assign n17622 = n15501 | n15516;
  assign n17623 = n11773 | n15516;
  assign n17624 = (n15485 & n17622) | (n15485 & n17623) | (n17622 & n17623);
  assign n11785 = ~n17621 & n17624;
  assign n15519 = n11782 | n17613;
  assign n17625 = n11782 | n17613;
  assign n17626 = (n11771 & n17613) | (n11771 & n17625) | (n17613 & n17625);
  assign n17627 = (n15501 & n15519) | (n15501 & n17626) | (n15519 & n17626);
  assign n17628 = (n11773 & n15519) | (n11773 & n17626) | (n15519 & n17626);
  assign n17629 = (n15485 & n17627) | (n15485 & n17628) | (n17627 & n17628);
  assign n17758 = x112 & x176;
  assign n17759 = x113 & x176;
  assign n17760 = x112 & x177;
  assign n17761 = n17759 & n17760;
  assign n17762 = n17759 | n17760;
  assign n17763 = ~n17761 & n17762;
  assign n17764 = x114 & x176;
  assign n17765 = x113 & x177;
  assign n17766 = n17764 & n17765;
  assign n17767 = n17764 | n17765;
  assign n17768 = ~n17766 & n17767;
  assign n17769 = n17761 & n17768;
  assign n17770 = n17761 | n17768;
  assign n17771 = ~n17769 & n17770;
  assign n17772 = x112 & x178;
  assign n17773 = n17771 & n17772;
  assign n17774 = n17771 | n17772;
  assign n17775 = ~n17773 & n17774;
  assign n50113 = n17761 | n17766;
  assign n50114 = (n17766 & n17768) | (n17766 & n50113) | (n17768 & n50113);
  assign n17777 = x115 & x176;
  assign n17778 = x114 & x177;
  assign n17779 = n17777 & n17778;
  assign n17780 = n17777 | n17778;
  assign n17781 = ~n17779 & n17780;
  assign n17782 = n50114 & n17781;
  assign n17783 = n50114 | n17781;
  assign n17784 = ~n17782 & n17783;
  assign n17785 = x113 & x178;
  assign n17786 = n17784 & n17785;
  assign n17787 = n17784 | n17785;
  assign n17788 = ~n17786 & n17787;
  assign n17789 = n17773 & n17788;
  assign n17790 = n17773 | n17788;
  assign n17791 = ~n17789 & n17790;
  assign n17792 = x112 & x179;
  assign n17793 = n17791 & n17792;
  assign n17794 = n17791 | n17792;
  assign n17795 = ~n17793 & n17794;
  assign n50115 = n17773 | n17786;
  assign n50116 = (n17786 & n17788) | (n17786 & n50115) | (n17788 & n50115);
  assign n50117 = n17779 | n17781;
  assign n50118 = (n17779 & n50114) | (n17779 & n50117) | (n50114 & n50117);
  assign n17798 = x116 & x176;
  assign n17799 = x115 & x177;
  assign n17800 = n17798 & n17799;
  assign n17801 = n17798 | n17799;
  assign n17802 = ~n17800 & n17801;
  assign n17803 = n50118 & n17802;
  assign n17804 = n50118 | n17802;
  assign n17805 = ~n17803 & n17804;
  assign n17806 = x114 & x178;
  assign n17807 = n17805 & n17806;
  assign n17808 = n17805 | n17806;
  assign n17809 = ~n17807 & n17808;
  assign n17810 = n50116 & n17809;
  assign n17811 = n50116 | n17809;
  assign n17812 = ~n17810 & n17811;
  assign n17813 = x113 & x179;
  assign n17814 = n17812 & n17813;
  assign n17815 = n17812 | n17813;
  assign n17816 = ~n17814 & n17815;
  assign n17817 = n17793 & n17816;
  assign n17818 = n17793 | n17816;
  assign n17819 = ~n17817 & n17818;
  assign n17820 = x112 & x180;
  assign n17821 = n17819 & n17820;
  assign n17822 = n17819 | n17820;
  assign n17823 = ~n17821 & n17822;
  assign n50119 = n17793 | n17814;
  assign n50120 = (n17814 & n17816) | (n17814 & n50119) | (n17816 & n50119);
  assign n17827 = x117 & x176;
  assign n17828 = x116 & x177;
  assign n17829 = n17827 & n17828;
  assign n17830 = n17827 | n17828;
  assign n17831 = ~n17829 & n17830;
  assign n50121 = n17800 | n17802;
  assign n50123 = n17831 & n50121;
  assign n50124 = n17800 & n17831;
  assign n50125 = (n50118 & n50123) | (n50118 & n50124) | (n50123 & n50124);
  assign n50126 = n17831 | n50121;
  assign n50127 = n17800 | n17831;
  assign n50128 = (n50118 & n50126) | (n50118 & n50127) | (n50126 & n50127);
  assign n17834 = ~n50125 & n50128;
  assign n17835 = x115 & x178;
  assign n17836 = n17834 & n17835;
  assign n17837 = n17834 | n17835;
  assign n17838 = ~n17836 & n17837;
  assign n50129 = n17807 & n17838;
  assign n50130 = (n17810 & n17838) | (n17810 & n50129) | (n17838 & n50129);
  assign n50131 = n17807 | n17838;
  assign n50132 = n17810 | n50131;
  assign n17841 = ~n50130 & n50132;
  assign n17842 = x114 & x179;
  assign n17843 = n17841 & n17842;
  assign n17844 = n17841 | n17842;
  assign n17845 = ~n17843 & n17844;
  assign n17846 = n50120 & n17845;
  assign n17847 = n50120 | n17845;
  assign n17848 = ~n17846 & n17847;
  assign n17849 = x113 & x180;
  assign n17850 = n17848 & n17849;
  assign n17851 = n17848 | n17849;
  assign n17852 = ~n17850 & n17851;
  assign n17853 = n17821 & n17852;
  assign n17854 = n17821 | n17852;
  assign n17855 = ~n17853 & n17854;
  assign n17856 = x112 & x181;
  assign n17857 = n17855 & n17856;
  assign n17858 = n17855 | n17856;
  assign n17859 = ~n17857 & n17858;
  assign n50133 = n17821 | n17850;
  assign n50134 = (n17850 & n17852) | (n17850 & n50133) | (n17852 & n50133);
  assign n17861 = n17843 | n17846;
  assign n17864 = x118 & x176;
  assign n17865 = x117 & x177;
  assign n17866 = n17864 & n17865;
  assign n17867 = n17864 | n17865;
  assign n17868 = ~n17866 & n17867;
  assign n50135 = n17829 & n17868;
  assign n50136 = (n17868 & n50125) | (n17868 & n50135) | (n50125 & n50135);
  assign n50137 = n17829 | n17868;
  assign n50138 = n50125 | n50137;
  assign n17871 = ~n50136 & n50138;
  assign n17872 = x116 & x178;
  assign n17873 = n17871 & n17872;
  assign n17874 = n17871 | n17872;
  assign n17875 = ~n17873 & n17874;
  assign n50139 = n17836 & n17875;
  assign n50140 = (n17875 & n50130) | (n17875 & n50139) | (n50130 & n50139);
  assign n50141 = n17836 | n17875;
  assign n50142 = n50130 | n50141;
  assign n17878 = ~n50140 & n50142;
  assign n17879 = x115 & x179;
  assign n17880 = n17878 & n17879;
  assign n17881 = n17878 | n17879;
  assign n17882 = ~n17880 & n17881;
  assign n17883 = n17861 & n17882;
  assign n17884 = n17861 | n17882;
  assign n17885 = ~n17883 & n17884;
  assign n17886 = x114 & x180;
  assign n17887 = n17885 & n17886;
  assign n17888 = n17885 | n17886;
  assign n17889 = ~n17887 & n17888;
  assign n17890 = n50134 & n17889;
  assign n17891 = n50134 | n17889;
  assign n17892 = ~n17890 & n17891;
  assign n17893 = x113 & x181;
  assign n17894 = n17892 & n17893;
  assign n17895 = n17892 | n17893;
  assign n17896 = ~n17894 & n17895;
  assign n17897 = n17857 & n17896;
  assign n17898 = n17857 | n17896;
  assign n17899 = ~n17897 & n17898;
  assign n17900 = x112 & x182;
  assign n17901 = n17899 & n17900;
  assign n17902 = n17899 | n17900;
  assign n17903 = ~n17901 & n17902;
  assign n66475 = n17857 | n17893;
  assign n66476 = (n17857 & n17892) | (n17857 & n66475) | (n17892 & n66475);
  assign n50144 = (n17894 & n17896) | (n17894 & n66476) | (n17896 & n66476);
  assign n50145 = n17887 | n50134;
  assign n50146 = (n17887 & n17889) | (n17887 & n50145) | (n17889 & n50145);
  assign n50147 = n17880 | n17882;
  assign n50148 = (n17861 & n17880) | (n17861 & n50147) | (n17880 & n50147);
  assign n17909 = x119 & x176;
  assign n17910 = x118 & x177;
  assign n17911 = n17909 & n17910;
  assign n17912 = n17909 | n17910;
  assign n17913 = ~n17911 & n17912;
  assign n66477 = n17829 | n17866;
  assign n66478 = (n17866 & n17868) | (n17866 & n66477) | (n17868 & n66477);
  assign n50152 = n17913 & n66478;
  assign n50150 = n17866 | n17868;
  assign n50153 = n17913 & n50150;
  assign n50154 = (n50125 & n50152) | (n50125 & n50153) | (n50152 & n50153);
  assign n50155 = n17913 | n66478;
  assign n50156 = n17913 | n50150;
  assign n50157 = (n50125 & n50155) | (n50125 & n50156) | (n50155 & n50156);
  assign n17916 = ~n50154 & n50157;
  assign n17917 = x117 & x178;
  assign n17918 = n17916 & n17917;
  assign n17919 = n17916 | n17917;
  assign n17920 = ~n17918 & n17919;
  assign n50158 = n17873 & n17920;
  assign n50159 = (n17920 & n50140) | (n17920 & n50158) | (n50140 & n50158);
  assign n50160 = n17873 | n17920;
  assign n50161 = n50140 | n50160;
  assign n17923 = ~n50159 & n50161;
  assign n17924 = x116 & x179;
  assign n17925 = n17923 & n17924;
  assign n17926 = n17923 | n17924;
  assign n17927 = ~n17925 & n17926;
  assign n17928 = n50148 & n17927;
  assign n17929 = n50148 | n17927;
  assign n17930 = ~n17928 & n17929;
  assign n17931 = x115 & x180;
  assign n17932 = n17930 & n17931;
  assign n17933 = n17930 | n17931;
  assign n17934 = ~n17932 & n17933;
  assign n17935 = n50146 & n17934;
  assign n17936 = n50146 | n17934;
  assign n17937 = ~n17935 & n17936;
  assign n17938 = x114 & x181;
  assign n17939 = n17937 & n17938;
  assign n17940 = n17937 | n17938;
  assign n17941 = ~n17939 & n17940;
  assign n17942 = n50144 & n17941;
  assign n17943 = n50144 | n17941;
  assign n17944 = ~n17942 & n17943;
  assign n17945 = x113 & x182;
  assign n17946 = n17944 & n17945;
  assign n17947 = n17944 | n17945;
  assign n17948 = ~n17946 & n17947;
  assign n17949 = n17901 & n17948;
  assign n17950 = n17901 | n17948;
  assign n17951 = ~n17949 & n17950;
  assign n17952 = x112 & x183;
  assign n17953 = n17951 & n17952;
  assign n17954 = n17951 | n17952;
  assign n17955 = ~n17953 & n17954;
  assign n50162 = n17901 | n17946;
  assign n50163 = (n17946 & n17948) | (n17946 & n50162) | (n17948 & n50162);
  assign n17957 = n17939 | n17942;
  assign n17958 = n17932 | n17935;
  assign n50164 = n17925 | n17927;
  assign n50165 = (n17925 & n50148) | (n17925 & n50164) | (n50148 & n50164);
  assign n17962 = x120 & x176;
  assign n17963 = x119 & x177;
  assign n17964 = n17962 & n17963;
  assign n17965 = n17962 | n17963;
  assign n17966 = ~n17964 & n17965;
  assign n50169 = n17911 & n17966;
  assign n66481 = (n17966 & n50153) | (n17966 & n50169) | (n50153 & n50169);
  assign n66482 = (n17966 & n50152) | (n17966 & n50169) | (n50152 & n50169);
  assign n66483 = (n50125 & n66481) | (n50125 & n66482) | (n66481 & n66482);
  assign n50171 = n17911 | n17966;
  assign n66484 = n50153 | n50171;
  assign n66485 = n50152 | n50171;
  assign n66486 = (n50125 & n66484) | (n50125 & n66485) | (n66484 & n66485);
  assign n17969 = ~n66483 & n66486;
  assign n17970 = x118 & x178;
  assign n17971 = n17969 & n17970;
  assign n17972 = n17969 | n17970;
  assign n17973 = ~n17971 & n17972;
  assign n50167 = n17918 | n17920;
  assign n66487 = n17973 & n50167;
  assign n66479 = n17873 | n17918;
  assign n66480 = (n17918 & n17920) | (n17918 & n66479) | (n17920 & n66479);
  assign n66488 = n17973 & n66480;
  assign n66489 = (n50140 & n66487) | (n50140 & n66488) | (n66487 & n66488);
  assign n66490 = n17973 | n50167;
  assign n66491 = n17973 | n66480;
  assign n66492 = (n50140 & n66490) | (n50140 & n66491) | (n66490 & n66491);
  assign n17976 = ~n66489 & n66492;
  assign n17977 = x117 & x179;
  assign n17978 = n17976 & n17977;
  assign n17979 = n17976 | n17977;
  assign n17980 = ~n17978 & n17979;
  assign n17981 = n50165 & n17980;
  assign n17982 = n50165 | n17980;
  assign n17983 = ~n17981 & n17982;
  assign n17984 = x116 & x180;
  assign n17985 = n17983 & n17984;
  assign n17986 = n17983 | n17984;
  assign n17987 = ~n17985 & n17986;
  assign n17988 = n17958 & n17987;
  assign n17989 = n17958 | n17987;
  assign n17990 = ~n17988 & n17989;
  assign n17991 = x115 & x181;
  assign n17992 = n17990 & n17991;
  assign n17993 = n17990 | n17991;
  assign n17994 = ~n17992 & n17993;
  assign n17995 = n17957 & n17994;
  assign n17996 = n17957 | n17994;
  assign n17997 = ~n17995 & n17996;
  assign n17998 = x114 & x182;
  assign n17999 = n17997 & n17998;
  assign n18000 = n17997 | n17998;
  assign n18001 = ~n17999 & n18000;
  assign n18002 = n50163 & n18001;
  assign n18003 = n50163 | n18001;
  assign n18004 = ~n18002 & n18003;
  assign n18005 = x113 & x183;
  assign n18006 = n18004 & n18005;
  assign n18007 = n18004 | n18005;
  assign n18008 = ~n18006 & n18007;
  assign n18009 = n17953 & n18008;
  assign n18010 = n17953 | n18008;
  assign n18011 = ~n18009 & n18010;
  assign n18012 = x112 & x184;
  assign n18013 = n18011 & n18012;
  assign n18014 = n18011 | n18012;
  assign n18015 = ~n18013 & n18014;
  assign n66493 = n17953 | n18005;
  assign n66494 = (n17953 & n18004) | (n17953 & n66493) | (n18004 & n66493);
  assign n50174 = (n18006 & n18008) | (n18006 & n66494) | (n18008 & n66494);
  assign n50175 = n17999 | n50163;
  assign n50176 = (n17999 & n18001) | (n17999 & n50175) | (n18001 & n50175);
  assign n18018 = n17992 | n17995;
  assign n50177 = n17985 | n17987;
  assign n50178 = (n17958 & n17985) | (n17958 & n50177) | (n17985 & n50177);
  assign n50168 = (n50140 & n66480) | (n50140 & n50167) | (n66480 & n50167);
  assign n18023 = x121 & x176;
  assign n18024 = x120 & x177;
  assign n18025 = n18023 & n18024;
  assign n18026 = n18023 | n18024;
  assign n18027 = ~n18025 & n18026;
  assign n66495 = n17911 | n17964;
  assign n66496 = (n17964 & n17966) | (n17964 & n66495) | (n17966 & n66495);
  assign n50186 = n18027 & n66496;
  assign n50184 = n17964 | n17966;
  assign n50187 = n18027 & n50184;
  assign n66497 = (n50153 & n50186) | (n50153 & n50187) | (n50186 & n50187);
  assign n66498 = (n50152 & n50186) | (n50152 & n50187) | (n50186 & n50187);
  assign n66499 = (n50125 & n66497) | (n50125 & n66498) | (n66497 & n66498);
  assign n50189 = n18027 | n66496;
  assign n50190 = n18027 | n50184;
  assign n66500 = (n50153 & n50189) | (n50153 & n50190) | (n50189 & n50190);
  assign n66501 = (n50152 & n50189) | (n50152 & n50190) | (n50189 & n50190);
  assign n66502 = (n50125 & n66500) | (n50125 & n66501) | (n66500 & n66501);
  assign n18030 = ~n66499 & n66502;
  assign n18031 = x119 & x178;
  assign n18032 = n18030 & n18031;
  assign n18033 = n18030 | n18031;
  assign n18034 = ~n18032 & n18033;
  assign n50181 = n17971 | n17973;
  assign n50192 = n18034 & n50181;
  assign n50193 = n17971 & n18034;
  assign n50194 = (n50168 & n50192) | (n50168 & n50193) | (n50192 & n50193);
  assign n50195 = n18034 | n50181;
  assign n50196 = n17971 | n18034;
  assign n50197 = (n50168 & n50195) | (n50168 & n50196) | (n50195 & n50196);
  assign n18037 = ~n50194 & n50197;
  assign n18038 = x118 & x179;
  assign n18039 = n18037 & n18038;
  assign n18040 = n18037 | n18038;
  assign n18041 = ~n18039 & n18040;
  assign n50179 = n17978 | n17980;
  assign n66503 = n18041 & n50179;
  assign n66504 = n17978 & n18041;
  assign n66505 = (n50165 & n66503) | (n50165 & n66504) | (n66503 & n66504);
  assign n66506 = n18041 | n50179;
  assign n66507 = n17978 | n18041;
  assign n66508 = (n50165 & n66506) | (n50165 & n66507) | (n66506 & n66507);
  assign n18044 = ~n66505 & n66508;
  assign n18045 = x117 & x180;
  assign n18046 = n18044 & n18045;
  assign n18047 = n18044 | n18045;
  assign n18048 = ~n18046 & n18047;
  assign n18049 = n50178 & n18048;
  assign n18050 = n50178 | n18048;
  assign n18051 = ~n18049 & n18050;
  assign n18052 = x116 & x181;
  assign n18053 = n18051 & n18052;
  assign n18054 = n18051 | n18052;
  assign n18055 = ~n18053 & n18054;
  assign n18056 = n18018 & n18055;
  assign n18057 = n18018 | n18055;
  assign n18058 = ~n18056 & n18057;
  assign n18059 = x115 & x182;
  assign n18060 = n18058 & n18059;
  assign n18061 = n18058 | n18059;
  assign n18062 = ~n18060 & n18061;
  assign n18063 = n50176 & n18062;
  assign n18064 = n50176 | n18062;
  assign n18065 = ~n18063 & n18064;
  assign n18066 = x114 & x183;
  assign n18067 = n18065 & n18066;
  assign n18068 = n18065 | n18066;
  assign n18069 = ~n18067 & n18068;
  assign n18070 = n50174 & n18069;
  assign n18071 = n50174 | n18069;
  assign n18072 = ~n18070 & n18071;
  assign n18073 = x113 & x184;
  assign n18074 = n18072 & n18073;
  assign n18075 = n18072 | n18073;
  assign n18076 = ~n18074 & n18075;
  assign n18077 = n18013 & n18076;
  assign n18078 = n18013 | n18076;
  assign n18079 = ~n18077 & n18078;
  assign n18080 = x112 & x185;
  assign n18081 = n18079 & n18080;
  assign n18082 = n18079 | n18080;
  assign n18083 = ~n18081 & n18082;
  assign n66509 = n18013 | n18073;
  assign n66510 = (n18013 & n18072) | (n18013 & n66509) | (n18072 & n66509);
  assign n50199 = (n18074 & n18076) | (n18074 & n66510) | (n18076 & n66510);
  assign n50200 = n18067 | n50174;
  assign n50201 = (n18067 & n18069) | (n18067 & n50200) | (n18069 & n50200);
  assign n50202 = n18060 | n50176;
  assign n50203 = (n18060 & n18062) | (n18060 & n50202) | (n18062 & n50202);
  assign n50204 = n18053 | n18055;
  assign n50205 = (n18018 & n18053) | (n18018 & n50204) | (n18053 & n50204);
  assign n50180 = (n17978 & n50165) | (n17978 & n50179) | (n50165 & n50179);
  assign n66511 = n18025 | n18027;
  assign n66512 = (n18025 & n66496) | (n18025 & n66511) | (n66496 & n66511);
  assign n66513 = (n18025 & n50184) | (n18025 & n66511) | (n50184 & n66511);
  assign n66514 = (n50153 & n66512) | (n50153 & n66513) | (n66512 & n66513);
  assign n66515 = (n50152 & n66512) | (n50152 & n66513) | (n66512 & n66513);
  assign n66516 = (n50125 & n66514) | (n50125 & n66515) | (n66514 & n66515);
  assign n18092 = x122 & x176;
  assign n18093 = x121 & x177;
  assign n18094 = n18092 & n18093;
  assign n18095 = n18092 | n18093;
  assign n18096 = ~n18094 & n18095;
  assign n18097 = n66516 & n18096;
  assign n18098 = n66516 | n18096;
  assign n18099 = ~n18097 & n18098;
  assign n18100 = x120 & x178;
  assign n18101 = n18099 & n18100;
  assign n18102 = n18099 | n18100;
  assign n18103 = ~n18101 & n18102;
  assign n50213 = n18032 & n18103;
  assign n66517 = (n18103 & n50192) | (n18103 & n50213) | (n50192 & n50213);
  assign n66518 = (n18103 & n50193) | (n18103 & n50213) | (n50193 & n50213);
  assign n66519 = (n50168 & n66517) | (n50168 & n66518) | (n66517 & n66518);
  assign n50215 = n18032 | n18103;
  assign n66520 = n50192 | n50215;
  assign n66521 = n50193 | n50215;
  assign n66522 = (n50168 & n66520) | (n50168 & n66521) | (n66520 & n66521);
  assign n18106 = ~n66519 & n66522;
  assign n18107 = x119 & x179;
  assign n18108 = n18106 & n18107;
  assign n18109 = n18106 | n18107;
  assign n18110 = ~n18108 & n18109;
  assign n50208 = n18039 | n18041;
  assign n50217 = n18110 & n50208;
  assign n50218 = n18039 & n18110;
  assign n50219 = (n50180 & n50217) | (n50180 & n50218) | (n50217 & n50218);
  assign n50220 = n18110 | n50208;
  assign n50221 = n18039 | n18110;
  assign n50222 = (n50180 & n50220) | (n50180 & n50221) | (n50220 & n50221);
  assign n18113 = ~n50219 & n50222;
  assign n18114 = x118 & x180;
  assign n18115 = n18113 & n18114;
  assign n18116 = n18113 | n18114;
  assign n18117 = ~n18115 & n18116;
  assign n50206 = n18046 | n18048;
  assign n66523 = n18117 & n50206;
  assign n66524 = n18046 & n18117;
  assign n66525 = (n50178 & n66523) | (n50178 & n66524) | (n66523 & n66524);
  assign n66526 = n18117 | n50206;
  assign n66527 = n18046 | n18117;
  assign n66528 = (n50178 & n66526) | (n50178 & n66527) | (n66526 & n66527);
  assign n18120 = ~n66525 & n66528;
  assign n18121 = x117 & x181;
  assign n18122 = n18120 & n18121;
  assign n18123 = n18120 | n18121;
  assign n18124 = ~n18122 & n18123;
  assign n18125 = n50205 & n18124;
  assign n18126 = n50205 | n18124;
  assign n18127 = ~n18125 & n18126;
  assign n18128 = x116 & x182;
  assign n18129 = n18127 & n18128;
  assign n18130 = n18127 | n18128;
  assign n18131 = ~n18129 & n18130;
  assign n18132 = n50203 & n18131;
  assign n18133 = n50203 | n18131;
  assign n18134 = ~n18132 & n18133;
  assign n18135 = x115 & x183;
  assign n18136 = n18134 & n18135;
  assign n18137 = n18134 | n18135;
  assign n18138 = ~n18136 & n18137;
  assign n18139 = n50201 & n18138;
  assign n18140 = n50201 | n18138;
  assign n18141 = ~n18139 & n18140;
  assign n18142 = x114 & x184;
  assign n18143 = n18141 & n18142;
  assign n18144 = n18141 | n18142;
  assign n18145 = ~n18143 & n18144;
  assign n18146 = n50199 & n18145;
  assign n18147 = n50199 | n18145;
  assign n18148 = ~n18146 & n18147;
  assign n18149 = x113 & x185;
  assign n18150 = n18148 & n18149;
  assign n18151 = n18148 | n18149;
  assign n18152 = ~n18150 & n18151;
  assign n18153 = n18081 & n18152;
  assign n18154 = n18081 | n18152;
  assign n18155 = ~n18153 & n18154;
  assign n18156 = x112 & x186;
  assign n18157 = n18155 & n18156;
  assign n18158 = n18155 | n18156;
  assign n18159 = ~n18157 & n18158;
  assign n50223 = n18081 | n18150;
  assign n50224 = (n18150 & n18152) | (n18150 & n50223) | (n18152 & n50223);
  assign n18161 = n18143 | n18146;
  assign n18162 = n18136 | n18139;
  assign n50207 = (n18046 & n50178) | (n18046 & n50206) | (n50178 & n50206);
  assign n50230 = n18101 | n18103;
  assign n66529 = n18032 | n18101;
  assign n66530 = (n18101 & n18103) | (n18101 & n66529) | (n18103 & n66529);
  assign n66531 = (n50192 & n50230) | (n50192 & n66530) | (n50230 & n66530);
  assign n66532 = (n50193 & n50230) | (n50193 & n66530) | (n50230 & n66530);
  assign n66533 = (n50168 & n66531) | (n50168 & n66532) | (n66531 & n66532);
  assign n18169 = x123 & x176;
  assign n18170 = x122 & x177;
  assign n18171 = n18169 & n18170;
  assign n18172 = n18169 | n18170;
  assign n18173 = ~n18171 & n18172;
  assign n50232 = n18094 | n18096;
  assign n50234 = n18173 & n50232;
  assign n50235 = n18094 & n18173;
  assign n50236 = (n66516 & n50234) | (n66516 & n50235) | (n50234 & n50235);
  assign n50237 = n18173 | n50232;
  assign n50238 = n18094 | n18173;
  assign n50239 = (n66516 & n50237) | (n66516 & n50238) | (n50237 & n50238);
  assign n18176 = ~n50236 & n50239;
  assign n18177 = x121 & x178;
  assign n18178 = n18176 & n18177;
  assign n18179 = n18176 | n18177;
  assign n18180 = ~n18178 & n18179;
  assign n18181 = n66533 & n18180;
  assign n18182 = n66533 | n18180;
  assign n18183 = ~n18181 & n18182;
  assign n18184 = x120 & x179;
  assign n18185 = n18183 & n18184;
  assign n18186 = n18183 | n18184;
  assign n18187 = ~n18185 & n18186;
  assign n50240 = n18108 & n18187;
  assign n50241 = (n18187 & n50219) | (n18187 & n50240) | (n50219 & n50240);
  assign n50242 = n18108 | n18187;
  assign n50243 = n50219 | n50242;
  assign n18190 = ~n50241 & n50243;
  assign n18191 = x119 & x180;
  assign n18192 = n18190 & n18191;
  assign n18193 = n18190 | n18191;
  assign n18194 = ~n18192 & n18193;
  assign n50227 = n18115 | n18117;
  assign n50244 = n18194 & n50227;
  assign n50245 = n18115 & n18194;
  assign n50246 = (n50207 & n50244) | (n50207 & n50245) | (n50244 & n50245);
  assign n50247 = n18194 | n50227;
  assign n50248 = n18115 | n18194;
  assign n50249 = (n50207 & n50247) | (n50207 & n50248) | (n50247 & n50248);
  assign n18197 = ~n50246 & n50249;
  assign n18198 = x118 & x181;
  assign n18199 = n18197 & n18198;
  assign n18200 = n18197 | n18198;
  assign n18201 = ~n18199 & n18200;
  assign n50225 = n18122 | n18124;
  assign n66534 = n18201 & n50225;
  assign n66535 = n18122 & n18201;
  assign n66536 = (n50205 & n66534) | (n50205 & n66535) | (n66534 & n66535);
  assign n66537 = n18201 | n50225;
  assign n66538 = n18122 | n18201;
  assign n66539 = (n50205 & n66537) | (n50205 & n66538) | (n66537 & n66538);
  assign n18204 = ~n66536 & n66539;
  assign n18205 = x117 & x182;
  assign n18206 = n18204 & n18205;
  assign n18207 = n18204 | n18205;
  assign n18208 = ~n18206 & n18207;
  assign n66540 = n18129 & n18208;
  assign n66541 = (n18132 & n18208) | (n18132 & n66540) | (n18208 & n66540);
  assign n66542 = n18129 | n18208;
  assign n66543 = n18132 | n66542;
  assign n18211 = ~n66541 & n66543;
  assign n18212 = x116 & x183;
  assign n18213 = n18211 & n18212;
  assign n18214 = n18211 | n18212;
  assign n18215 = ~n18213 & n18214;
  assign n18216 = n18162 & n18215;
  assign n18217 = n18162 | n18215;
  assign n18218 = ~n18216 & n18217;
  assign n18219 = x115 & x184;
  assign n18220 = n18218 & n18219;
  assign n18221 = n18218 | n18219;
  assign n18222 = ~n18220 & n18221;
  assign n18223 = n18161 & n18222;
  assign n18224 = n18161 | n18222;
  assign n18225 = ~n18223 & n18224;
  assign n18226 = x114 & x185;
  assign n18227 = n18225 & n18226;
  assign n18228 = n18225 | n18226;
  assign n18229 = ~n18227 & n18228;
  assign n18230 = n50224 & n18229;
  assign n18231 = n50224 | n18229;
  assign n18232 = ~n18230 & n18231;
  assign n18233 = x113 & x186;
  assign n18234 = n18232 & n18233;
  assign n18235 = n18232 | n18233;
  assign n18236 = ~n18234 & n18235;
  assign n18237 = n18157 & n18236;
  assign n18238 = n18157 | n18236;
  assign n18239 = ~n18237 & n18238;
  assign n18240 = x112 & x187;
  assign n18241 = n18239 & n18240;
  assign n18242 = n18239 | n18240;
  assign n18243 = ~n18241 & n18242;
  assign n66544 = n18157 | n18233;
  assign n66545 = (n18157 & n18232) | (n18157 & n66544) | (n18232 & n66544);
  assign n50251 = (n18234 & n18236) | (n18234 & n66545) | (n18236 & n66545);
  assign n50252 = n18227 | n50224;
  assign n50253 = (n18227 & n18229) | (n18227 & n50252) | (n18229 & n50252);
  assign n18246 = n18220 | n18223;
  assign n66546 = n18213 | n18215;
  assign n66547 = (n18162 & n18213) | (n18162 & n66546) | (n18213 & n66546);
  assign n18163 = n18129 | n18132;
  assign n50226 = (n18122 & n50205) | (n18122 & n50225) | (n50205 & n50225);
  assign n18254 = x124 & x176;
  assign n18255 = x123 & x177;
  assign n18256 = n18254 & n18255;
  assign n18257 = n18254 | n18255;
  assign n18258 = ~n18256 & n18257;
  assign n66548 = n18171 | n18173;
  assign n66549 = (n18171 & n50232) | (n18171 & n66548) | (n50232 & n66548);
  assign n50263 = n18258 & n66549;
  assign n66550 = n18094 | n18171;
  assign n66551 = (n18171 & n18173) | (n18171 & n66550) | (n18173 & n66550);
  assign n50264 = n18258 & n66551;
  assign n50265 = (n66516 & n50263) | (n66516 & n50264) | (n50263 & n50264);
  assign n50266 = n18258 | n66549;
  assign n50267 = n18258 | n66551;
  assign n50268 = (n66516 & n50266) | (n66516 & n50267) | (n50266 & n50267);
  assign n18261 = ~n50265 & n50268;
  assign n18262 = x122 & x178;
  assign n18263 = n18261 & n18262;
  assign n18264 = n18261 | n18262;
  assign n18265 = ~n18263 & n18264;
  assign n50258 = n18178 | n18180;
  assign n50269 = n18265 & n50258;
  assign n50270 = n18178 & n18265;
  assign n50271 = (n66533 & n50269) | (n66533 & n50270) | (n50269 & n50270);
  assign n50272 = n18265 | n50258;
  assign n50273 = n18178 | n18265;
  assign n50274 = (n66533 & n50272) | (n66533 & n50273) | (n50272 & n50273);
  assign n18268 = ~n50271 & n50274;
  assign n18269 = x121 & x179;
  assign n18270 = n18268 & n18269;
  assign n18271 = n18268 | n18269;
  assign n18272 = ~n18270 & n18271;
  assign n50275 = n18185 & n18272;
  assign n66552 = (n18272 & n50240) | (n18272 & n50275) | (n50240 & n50275);
  assign n66553 = (n18187 & n18272) | (n18187 & n50275) | (n18272 & n50275);
  assign n66554 = (n50219 & n66552) | (n50219 & n66553) | (n66552 & n66553);
  assign n50277 = n18185 | n18272;
  assign n66555 = n50240 | n50277;
  assign n66556 = n18187 | n50277;
  assign n66557 = (n50219 & n66555) | (n50219 & n66556) | (n66555 & n66556);
  assign n18275 = ~n66554 & n66557;
  assign n18276 = x120 & x180;
  assign n18277 = n18275 & n18276;
  assign n18278 = n18275 | n18276;
  assign n18279 = ~n18277 & n18278;
  assign n50279 = n18192 & n18279;
  assign n50280 = (n18279 & n50246) | (n18279 & n50279) | (n50246 & n50279);
  assign n50281 = n18192 | n18279;
  assign n50282 = n50246 | n50281;
  assign n18282 = ~n50280 & n50282;
  assign n18283 = x119 & x181;
  assign n18284 = n18282 & n18283;
  assign n18285 = n18282 | n18283;
  assign n18286 = ~n18284 & n18285;
  assign n50256 = n18199 | n18201;
  assign n50283 = n18286 & n50256;
  assign n50284 = n18199 & n18286;
  assign n50285 = (n50226 & n50283) | (n50226 & n50284) | (n50283 & n50284);
  assign n50286 = n18286 | n50256;
  assign n50287 = n18199 | n18286;
  assign n50288 = (n50226 & n50286) | (n50226 & n50287) | (n50286 & n50287);
  assign n18289 = ~n50285 & n50288;
  assign n18290 = x118 & x182;
  assign n18291 = n18289 & n18290;
  assign n18292 = n18289 | n18290;
  assign n18293 = ~n18291 & n18292;
  assign n50254 = n18206 | n18208;
  assign n66558 = n18293 & n50254;
  assign n66559 = n18206 & n18293;
  assign n66560 = (n18163 & n66558) | (n18163 & n66559) | (n66558 & n66559);
  assign n66561 = n18293 | n50254;
  assign n66562 = n18206 | n18293;
  assign n66563 = (n18163 & n66561) | (n18163 & n66562) | (n66561 & n66562);
  assign n18296 = ~n66560 & n66563;
  assign n18297 = x117 & x183;
  assign n18298 = n18296 & n18297;
  assign n18299 = n18296 | n18297;
  assign n18300 = ~n18298 & n18299;
  assign n18301 = n66547 & n18300;
  assign n18302 = n66547 | n18300;
  assign n18303 = ~n18301 & n18302;
  assign n18304 = x116 & x184;
  assign n18305 = n18303 & n18304;
  assign n18306 = n18303 | n18304;
  assign n18307 = ~n18305 & n18306;
  assign n18308 = n18246 & n18307;
  assign n18309 = n18246 | n18307;
  assign n18310 = ~n18308 & n18309;
  assign n18311 = x115 & x185;
  assign n18312 = n18310 & n18311;
  assign n18313 = n18310 | n18311;
  assign n18314 = ~n18312 & n18313;
  assign n18315 = n50253 & n18314;
  assign n18316 = n50253 | n18314;
  assign n18317 = ~n18315 & n18316;
  assign n18318 = x114 & x186;
  assign n18319 = n18317 & n18318;
  assign n18320 = n18317 | n18318;
  assign n18321 = ~n18319 & n18320;
  assign n18322 = n50251 & n18321;
  assign n18323 = n50251 | n18321;
  assign n18324 = ~n18322 & n18323;
  assign n18325 = x113 & x187;
  assign n18326 = n18324 & n18325;
  assign n18327 = n18324 | n18325;
  assign n18328 = ~n18326 & n18327;
  assign n18329 = n18241 & n18328;
  assign n18330 = n18241 | n18328;
  assign n18331 = ~n18329 & n18330;
  assign n18332 = x112 & x188;
  assign n18333 = n18331 & n18332;
  assign n18334 = n18331 | n18332;
  assign n18335 = ~n18333 & n18334;
  assign n66564 = n18241 | n18325;
  assign n66565 = (n18241 & n18324) | (n18241 & n66564) | (n18324 & n66564);
  assign n50290 = (n18326 & n18328) | (n18326 & n66565) | (n18328 & n66565);
  assign n50291 = n18319 | n50251;
  assign n50292 = (n18319 & n18321) | (n18319 & n50291) | (n18321 & n50291);
  assign n50293 = n18312 | n50253;
  assign n50294 = (n18312 & n18314) | (n18312 & n50293) | (n18314 & n50293);
  assign n66566 = n18305 | n18307;
  assign n66567 = (n18246 & n18305) | (n18246 & n66566) | (n18305 & n66566);
  assign n50295 = n18298 | n18300;
  assign n50296 = (n66547 & n18298) | (n66547 & n50295) | (n18298 & n50295);
  assign n50255 = (n18163 & n18206) | (n18163 & n50254) | (n18206 & n50254);
  assign n50300 = n18270 | n18272;
  assign n66568 = n18185 | n18270;
  assign n66569 = (n18270 & n18272) | (n18270 & n66568) | (n18272 & n66568);
  assign n66570 = (n50240 & n50300) | (n50240 & n66569) | (n50300 & n66569);
  assign n66571 = (n18187 & n50300) | (n18187 & n66569) | (n50300 & n66569);
  assign n66572 = (n50219 & n66570) | (n50219 & n66571) | (n66570 & n66571);
  assign n18347 = x125 & x176;
  assign n18348 = x124 & x177;
  assign n18349 = n18347 & n18348;
  assign n18350 = n18347 | n18348;
  assign n18351 = ~n18349 & n18350;
  assign n66577 = n18256 | n18258;
  assign n66578 = (n18256 & n66549) | (n18256 & n66577) | (n66549 & n66577);
  assign n66580 = n18351 & n66578;
  assign n66579 = (n18256 & n66551) | (n18256 & n66577) | (n66551 & n66577);
  assign n66581 = n18351 & n66579;
  assign n66582 = (n66516 & n66580) | (n66516 & n66581) | (n66580 & n66581);
  assign n66583 = n18351 | n66578;
  assign n66584 = n18351 | n66579;
  assign n66585 = (n66516 & n66583) | (n66516 & n66584) | (n66583 & n66584);
  assign n18354 = ~n66582 & n66585;
  assign n18355 = x123 & x178;
  assign n18356 = n18354 & n18355;
  assign n18357 = n18354 | n18355;
  assign n18358 = ~n18356 & n18357;
  assign n66573 = n18263 | n18265;
  assign n66574 = (n18263 & n50258) | (n18263 & n66573) | (n50258 & n66573);
  assign n66586 = n18358 & n66574;
  assign n66575 = n18178 | n18263;
  assign n66576 = (n18263 & n18265) | (n18263 & n66575) | (n18265 & n66575);
  assign n66587 = n18358 & n66576;
  assign n66588 = (n66533 & n66586) | (n66533 & n66587) | (n66586 & n66587);
  assign n66589 = n18358 | n66574;
  assign n66590 = n18358 | n66576;
  assign n66591 = (n66533 & n66589) | (n66533 & n66590) | (n66589 & n66590);
  assign n18361 = ~n66588 & n66591;
  assign n18362 = x122 & x179;
  assign n18363 = n18361 & n18362;
  assign n18364 = n18361 | n18362;
  assign n18365 = ~n18363 & n18364;
  assign n18366 = n66572 & n18365;
  assign n18367 = n66572 | n18365;
  assign n18368 = ~n18366 & n18367;
  assign n18369 = x121 & x180;
  assign n18370 = n18368 & n18369;
  assign n18371 = n18368 | n18369;
  assign n18372 = ~n18370 & n18371;
  assign n50308 = n18277 & n18372;
  assign n50309 = (n18372 & n50280) | (n18372 & n50308) | (n50280 & n50308);
  assign n50310 = n18277 | n18372;
  assign n50311 = n50280 | n50310;
  assign n18375 = ~n50309 & n50311;
  assign n18376 = x120 & x181;
  assign n18377 = n18375 & n18376;
  assign n18378 = n18375 | n18376;
  assign n18379 = ~n18377 & n18378;
  assign n50312 = n18284 & n18379;
  assign n50313 = (n18379 & n50285) | (n18379 & n50312) | (n50285 & n50312);
  assign n50314 = n18284 | n18379;
  assign n50315 = n50285 | n50314;
  assign n18382 = ~n50313 & n50315;
  assign n18383 = x119 & x182;
  assign n18384 = n18382 & n18383;
  assign n18385 = n18382 | n18383;
  assign n18386 = ~n18384 & n18385;
  assign n50297 = n18291 | n18293;
  assign n50316 = n18386 & n50297;
  assign n50317 = n18291 & n18386;
  assign n50318 = (n50255 & n50316) | (n50255 & n50317) | (n50316 & n50317);
  assign n50319 = n18386 | n50297;
  assign n50320 = n18291 | n18386;
  assign n50321 = (n50255 & n50319) | (n50255 & n50320) | (n50319 & n50320);
  assign n18389 = ~n50318 & n50321;
  assign n18390 = x118 & x183;
  assign n18391 = n18389 & n18390;
  assign n18392 = n18389 | n18390;
  assign n18393 = ~n18391 & n18392;
  assign n18394 = n50296 & n18393;
  assign n18395 = n50296 | n18393;
  assign n18396 = ~n18394 & n18395;
  assign n18397 = x117 & x184;
  assign n18398 = n18396 & n18397;
  assign n18399 = n18396 | n18397;
  assign n18400 = ~n18398 & n18399;
  assign n18401 = n66567 & n18400;
  assign n18402 = n66567 | n18400;
  assign n18403 = ~n18401 & n18402;
  assign n18404 = x116 & x185;
  assign n18405 = n18403 & n18404;
  assign n18406 = n18403 | n18404;
  assign n18407 = ~n18405 & n18406;
  assign n18408 = n50294 & n18407;
  assign n18409 = n50294 | n18407;
  assign n18410 = ~n18408 & n18409;
  assign n18411 = x115 & x186;
  assign n18412 = n18410 & n18411;
  assign n18413 = n18410 | n18411;
  assign n18414 = ~n18412 & n18413;
  assign n18415 = n50292 & n18414;
  assign n18416 = n50292 | n18414;
  assign n18417 = ~n18415 & n18416;
  assign n18418 = x114 & x187;
  assign n18419 = n18417 & n18418;
  assign n18420 = n18417 | n18418;
  assign n18421 = ~n18419 & n18420;
  assign n18422 = n50290 & n18421;
  assign n18423 = n50290 | n18421;
  assign n18424 = ~n18422 & n18423;
  assign n18425 = x113 & x188;
  assign n18426 = n18424 & n18425;
  assign n18427 = n18424 | n18425;
  assign n18428 = ~n18426 & n18427;
  assign n18429 = n18333 & n18428;
  assign n18430 = n18333 | n18428;
  assign n18431 = ~n18429 & n18430;
  assign n18432 = x112 & x189;
  assign n18433 = n18431 & n18432;
  assign n18434 = n18431 | n18432;
  assign n18435 = ~n18433 & n18434;
  assign n50322 = n18333 | n18426;
  assign n50323 = (n18426 & n18428) | (n18426 & n50322) | (n18428 & n50322);
  assign n50324 = n18419 | n50290;
  assign n50325 = (n18419 & n18421) | (n18419 & n50324) | (n18421 & n50324);
  assign n50326 = n18412 | n50292;
  assign n50327 = (n18412 & n18414) | (n18412 & n50326) | (n18414 & n50326);
  assign n50328 = n18405 | n50294;
  assign n50329 = (n18405 & n18407) | (n18405 & n50328) | (n18407 & n50328);
  assign n50330 = n18398 | n18400;
  assign n50331 = (n66567 & n18398) | (n66567 & n50330) | (n18398 & n50330);
  assign n18448 = x126 & x176;
  assign n18449 = x125 & x177;
  assign n18450 = n18448 & n18449;
  assign n18451 = n18448 | n18449;
  assign n18452 = ~n18450 & n18451;
  assign n50338 = n18349 | n18351;
  assign n50340 = n18452 & n50338;
  assign n50341 = n18349 & n18452;
  assign n66592 = (n50340 & n50341) | (n50340 & n66578) | (n50341 & n66578);
  assign n66593 = (n50340 & n50341) | (n50340 & n66579) | (n50341 & n66579);
  assign n66594 = (n66516 & n66592) | (n66516 & n66593) | (n66592 & n66593);
  assign n50343 = n18452 | n50338;
  assign n50344 = n18349 | n18452;
  assign n66595 = (n50343 & n50344) | (n50343 & n66578) | (n50344 & n66578);
  assign n66596 = (n50343 & n50344) | (n50343 & n66579) | (n50344 & n66579);
  assign n66597 = (n66516 & n66595) | (n66516 & n66596) | (n66595 & n66596);
  assign n18455 = ~n66594 & n66597;
  assign n18456 = x124 & x178;
  assign n18457 = n18455 & n18456;
  assign n18458 = n18455 | n18456;
  assign n18459 = ~n18457 & n18458;
  assign n50336 = n18356 | n18358;
  assign n50346 = n18459 & n50336;
  assign n50347 = n18356 & n18459;
  assign n66598 = (n50346 & n50347) | (n50346 & n66574) | (n50347 & n66574);
  assign n66599 = (n50346 & n50347) | (n50346 & n66576) | (n50347 & n66576);
  assign n66600 = (n66533 & n66598) | (n66533 & n66599) | (n66598 & n66599);
  assign n50349 = n18459 | n50336;
  assign n50350 = n18356 | n18459;
  assign n66601 = (n50349 & n50350) | (n50349 & n66574) | (n50350 & n66574);
  assign n66602 = (n50349 & n50350) | (n50349 & n66576) | (n50350 & n66576);
  assign n66603 = (n66533 & n66601) | (n66533 & n66602) | (n66601 & n66602);
  assign n18462 = ~n66600 & n66603;
  assign n18463 = x123 & x179;
  assign n18464 = n18462 & n18463;
  assign n18465 = n18462 | n18463;
  assign n18466 = ~n18464 & n18465;
  assign n50334 = n18363 | n18365;
  assign n50352 = n18466 & n50334;
  assign n50353 = n18363 & n18466;
  assign n50354 = (n66572 & n50352) | (n66572 & n50353) | (n50352 & n50353);
  assign n50355 = n18466 | n50334;
  assign n50356 = n18363 | n18466;
  assign n50357 = (n66572 & n50355) | (n66572 & n50356) | (n50355 & n50356);
  assign n18469 = ~n50354 & n50357;
  assign n18470 = x122 & x180;
  assign n18471 = n18469 & n18470;
  assign n18472 = n18469 | n18470;
  assign n18473 = ~n18471 & n18472;
  assign n50358 = n18370 & n18473;
  assign n66604 = (n18473 & n50308) | (n18473 & n50358) | (n50308 & n50358);
  assign n66605 = (n18372 & n18473) | (n18372 & n50358) | (n18473 & n50358);
  assign n66606 = (n50280 & n66604) | (n50280 & n66605) | (n66604 & n66605);
  assign n50360 = n18370 | n18473;
  assign n66607 = n50308 | n50360;
  assign n66608 = n18372 | n50360;
  assign n66609 = (n50280 & n66607) | (n50280 & n66608) | (n66607 & n66608);
  assign n18476 = ~n66606 & n66609;
  assign n18477 = x121 & x181;
  assign n18478 = n18476 & n18477;
  assign n18479 = n18476 | n18477;
  assign n18480 = ~n18478 & n18479;
  assign n50362 = n18377 & n18480;
  assign n50363 = (n18480 & n50313) | (n18480 & n50362) | (n50313 & n50362);
  assign n50364 = n18377 | n18480;
  assign n50365 = n50313 | n50364;
  assign n18483 = ~n50363 & n50365;
  assign n18484 = x120 & x182;
  assign n18485 = n18483 & n18484;
  assign n18486 = n18483 | n18484;
  assign n18487 = ~n18485 & n18486;
  assign n50366 = n18384 & n18487;
  assign n50367 = (n18487 & n50318) | (n18487 & n50366) | (n50318 & n50366);
  assign n50368 = n18384 | n18487;
  assign n50369 = n50318 | n50368;
  assign n18490 = ~n50367 & n50369;
  assign n18491 = x119 & x183;
  assign n18492 = n18490 & n18491;
  assign n18493 = n18490 | n18491;
  assign n18494 = ~n18492 & n18493;
  assign n50332 = n18391 | n18393;
  assign n50370 = n18494 & n50332;
  assign n50371 = n18391 & n18494;
  assign n50372 = (n50296 & n50370) | (n50296 & n50371) | (n50370 & n50371);
  assign n50373 = n18494 | n50332;
  assign n50374 = n18391 | n18494;
  assign n50375 = (n50296 & n50373) | (n50296 & n50374) | (n50373 & n50374);
  assign n18497 = ~n50372 & n50375;
  assign n18498 = x118 & x184;
  assign n18499 = n18497 & n18498;
  assign n18500 = n18497 | n18498;
  assign n18501 = ~n18499 & n18500;
  assign n18502 = n50331 & n18501;
  assign n18503 = n50331 | n18501;
  assign n18504 = ~n18502 & n18503;
  assign n18505 = x117 & x185;
  assign n18506 = n18504 & n18505;
  assign n18507 = n18504 | n18505;
  assign n18508 = ~n18506 & n18507;
  assign n18509 = n50329 & n18508;
  assign n18510 = n50329 | n18508;
  assign n18511 = ~n18509 & n18510;
  assign n18512 = x116 & x186;
  assign n18513 = n18511 & n18512;
  assign n18514 = n18511 | n18512;
  assign n18515 = ~n18513 & n18514;
  assign n18516 = n50327 & n18515;
  assign n18517 = n50327 | n18515;
  assign n18518 = ~n18516 & n18517;
  assign n18519 = x115 & x187;
  assign n18520 = n18518 & n18519;
  assign n18521 = n18518 | n18519;
  assign n18522 = ~n18520 & n18521;
  assign n18523 = n50325 & n18522;
  assign n18524 = n50325 | n18522;
  assign n18525 = ~n18523 & n18524;
  assign n18526 = x114 & x188;
  assign n18527 = n18525 & n18526;
  assign n18528 = n18525 | n18526;
  assign n18529 = ~n18527 & n18528;
  assign n18530 = n50323 & n18529;
  assign n18531 = n50323 | n18529;
  assign n18532 = ~n18530 & n18531;
  assign n18533 = x113 & x189;
  assign n18534 = n18532 & n18533;
  assign n18535 = n18532 | n18533;
  assign n18536 = ~n18534 & n18535;
  assign n18537 = n18433 & n18536;
  assign n18538 = n18433 | n18536;
  assign n18539 = ~n18537 & n18538;
  assign n18540 = x112 & x190;
  assign n18541 = n18539 & n18540;
  assign n18542 = n18539 | n18540;
  assign n18543 = ~n18541 & n18542;
  assign n66610 = n18433 | n18533;
  assign n66611 = (n18433 & n18532) | (n18433 & n66610) | (n18532 & n66610);
  assign n50377 = (n18534 & n18536) | (n18534 & n66611) | (n18536 & n66611);
  assign n66612 = n18527 | n50323;
  assign n66613 = (n18527 & n18529) | (n18527 & n66612) | (n18529 & n66612);
  assign n18546 = n18520 | n18523;
  assign n18547 = n18513 | n18516;
  assign n50381 = n18471 | n18473;
  assign n66614 = n18370 | n18471;
  assign n66615 = (n18471 & n18473) | (n18471 & n66614) | (n18473 & n66614);
  assign n66616 = (n50308 & n50381) | (n50308 & n66615) | (n50381 & n66615);
  assign n66617 = (n18372 & n50381) | (n18372 & n66615) | (n50381 & n66615);
  assign n66618 = (n50280 & n66616) | (n50280 & n66617) | (n66616 & n66617);
  assign n66619 = n18457 | n18459;
  assign n66620 = (n18457 & n50336) | (n18457 & n66619) | (n50336 & n66619);
  assign n66621 = n18356 | n18457;
  assign n66622 = (n18457 & n18459) | (n18457 & n66621) | (n18459 & n66621);
  assign n66623 = (n66574 & n66620) | (n66574 & n66622) | (n66620 & n66622);
  assign n66624 = (n66576 & n66620) | (n66576 & n66622) | (n66620 & n66622);
  assign n66625 = (n66533 & n66623) | (n66533 & n66624) | (n66623 & n66624);
  assign n18557 = x127 & x176;
  assign n18558 = x126 & x177;
  assign n18559 = n18557 & n18558;
  assign n18560 = n18557 | n18558;
  assign n18561 = ~n18559 & n18560;
  assign n66626 = n18450 | n18452;
  assign n66627 = (n18450 & n50338) | (n18450 & n66626) | (n50338 & n66626);
  assign n50389 = n18561 & n66627;
  assign n66628 = n18349 | n18450;
  assign n66629 = (n18450 & n18452) | (n18450 & n66628) | (n18452 & n66628);
  assign n50390 = n18561 & n66629;
  assign n66630 = (n50389 & n50390) | (n50389 & n66578) | (n50390 & n66578);
  assign n66631 = (n50389 & n50390) | (n50389 & n66579) | (n50390 & n66579);
  assign n66632 = (n66516 & n66630) | (n66516 & n66631) | (n66630 & n66631);
  assign n50392 = n18561 | n66627;
  assign n50393 = n18561 | n66629;
  assign n66633 = (n50392 & n50393) | (n50392 & n66578) | (n50393 & n66578);
  assign n66634 = (n50392 & n50393) | (n50392 & n66579) | (n50393 & n66579);
  assign n66635 = (n66516 & n66633) | (n66516 & n66634) | (n66633 & n66634);
  assign n18564 = ~n66632 & n66635;
  assign n18565 = x125 & x178;
  assign n18566 = n18564 & n18565;
  assign n18567 = n18564 | n18565;
  assign n18568 = ~n18566 & n18567;
  assign n18569 = n66625 & n18568;
  assign n18570 = n66625 | n18568;
  assign n18571 = ~n18569 & n18570;
  assign n18572 = x124 & x179;
  assign n18573 = n18571 & n18572;
  assign n18574 = n18571 | n18572;
  assign n18575 = ~n18573 & n18574;
  assign n50395 = n18464 & n18575;
  assign n66636 = (n18575 & n50352) | (n18575 & n50395) | (n50352 & n50395);
  assign n66637 = (n18575 & n50353) | (n18575 & n50395) | (n50353 & n50395);
  assign n66638 = (n66572 & n66636) | (n66572 & n66637) | (n66636 & n66637);
  assign n50397 = n18464 | n18575;
  assign n66639 = n50352 | n50397;
  assign n66640 = n50353 | n50397;
  assign n66641 = (n66572 & n66639) | (n66572 & n66640) | (n66639 & n66640);
  assign n18578 = ~n66638 & n66641;
  assign n18579 = x123 & x180;
  assign n18580 = n18578 & n18579;
  assign n18581 = n18578 | n18579;
  assign n18582 = ~n18580 & n18581;
  assign n18583 = n66618 & n18582;
  assign n18584 = n66618 | n18582;
  assign n18585 = ~n18583 & n18584;
  assign n18586 = x122 & x181;
  assign n18587 = n18585 & n18586;
  assign n18588 = n18585 | n18586;
  assign n18589 = ~n18587 & n18588;
  assign n50399 = n18478 & n18589;
  assign n50400 = (n18589 & n50363) | (n18589 & n50399) | (n50363 & n50399);
  assign n50401 = n18478 | n18589;
  assign n50402 = n50363 | n50401;
  assign n18592 = ~n50400 & n50402;
  assign n18593 = x121 & x182;
  assign n18594 = n18592 & n18593;
  assign n18595 = n18592 | n18593;
  assign n18596 = ~n18594 & n18595;
  assign n50403 = n18485 & n18596;
  assign n50404 = (n18596 & n50367) | (n18596 & n50403) | (n50367 & n50403);
  assign n50405 = n18485 | n18596;
  assign n50406 = n50367 | n50405;
  assign n18599 = ~n50404 & n50406;
  assign n18600 = x120 & x183;
  assign n18601 = n18599 & n18600;
  assign n18602 = n18599 | n18600;
  assign n18603 = ~n18601 & n18602;
  assign n50407 = n18492 & n18603;
  assign n50408 = (n18603 & n50372) | (n18603 & n50407) | (n50372 & n50407);
  assign n50409 = n18492 | n18603;
  assign n50410 = n50372 | n50409;
  assign n18606 = ~n50408 & n50410;
  assign n18607 = x119 & x184;
  assign n18608 = n18606 & n18607;
  assign n18609 = n18606 | n18607;
  assign n18610 = ~n18608 & n18609;
  assign n50378 = n18499 | n18501;
  assign n50411 = n18610 & n50378;
  assign n50412 = n18499 & n18610;
  assign n50413 = (n50331 & n50411) | (n50331 & n50412) | (n50411 & n50412);
  assign n50414 = n18610 | n50378;
  assign n50415 = n18499 | n18610;
  assign n50416 = (n50331 & n50414) | (n50331 & n50415) | (n50414 & n50415);
  assign n18613 = ~n50413 & n50416;
  assign n18614 = x118 & x185;
  assign n18615 = n18613 & n18614;
  assign n18616 = n18613 | n18614;
  assign n18617 = ~n18615 & n18616;
  assign n50417 = n18506 & n18617;
  assign n50418 = (n18509 & n18617) | (n18509 & n50417) | (n18617 & n50417);
  assign n50419 = n18506 | n18617;
  assign n50420 = n18509 | n50419;
  assign n18620 = ~n50418 & n50420;
  assign n18621 = x117 & x186;
  assign n18622 = n18620 & n18621;
  assign n18623 = n18620 | n18621;
  assign n18624 = ~n18622 & n18623;
  assign n18625 = n18547 & n18624;
  assign n18626 = n18547 | n18624;
  assign n18627 = ~n18625 & n18626;
  assign n18628 = x116 & x187;
  assign n18629 = n18627 & n18628;
  assign n18630 = n18627 | n18628;
  assign n18631 = ~n18629 & n18630;
  assign n18632 = n18546 & n18631;
  assign n18633 = n18546 | n18631;
  assign n18634 = ~n18632 & n18633;
  assign n18635 = x115 & x188;
  assign n18636 = n18634 & n18635;
  assign n18637 = n18634 | n18635;
  assign n18638 = ~n18636 & n18637;
  assign n18639 = n66613 & n18638;
  assign n18640 = n66613 | n18638;
  assign n18641 = ~n18639 & n18640;
  assign n18642 = x114 & x189;
  assign n18643 = n18641 & n18642;
  assign n18644 = n18641 | n18642;
  assign n18645 = ~n18643 & n18644;
  assign n18646 = n50377 & n18645;
  assign n18647 = n50377 | n18645;
  assign n18648 = ~n18646 & n18647;
  assign n18649 = x113 & x190;
  assign n18650 = n18648 & n18649;
  assign n18651 = n18648 | n18649;
  assign n18652 = ~n18650 & n18651;
  assign n18653 = n18541 & n18652;
  assign n18654 = n18541 | n18652;
  assign n18655 = ~n18653 & n18654;
  assign n18656 = x112 & x191;
  assign n18657 = n18655 & n18656;
  assign n18658 = n18655 | n18656;
  assign n18659 = ~n18657 & n18658;
  assign n66642 = n18541 | n18649;
  assign n66643 = (n18541 & n18648) | (n18541 & n66642) | (n18648 & n66642);
  assign n50422 = (n18650 & n18652) | (n18650 & n66643) | (n18652 & n66643);
  assign n50423 = n18643 | n50377;
  assign n50424 = (n18643 & n18645) | (n18643 & n50423) | (n18645 & n50423);
  assign n66644 = n18636 | n66613;
  assign n66645 = (n18636 & n18638) | (n18636 & n66644) | (n18638 & n66644);
  assign n18663 = n18629 | n18632;
  assign n50425 = n18622 | n18624;
  assign n50426 = (n18547 & n18622) | (n18547 & n50425) | (n18622 & n50425);
  assign n50430 = n18573 | n18575;
  assign n66646 = n18464 | n18573;
  assign n66647 = (n18573 & n18575) | (n18573 & n66646) | (n18575 & n66646);
  assign n66648 = (n50352 & n50430) | (n50352 & n66647) | (n50430 & n66647);
  assign n66649 = (n50353 & n50430) | (n50353 & n66647) | (n50430 & n66647);
  assign n66650 = (n66572 & n66648) | (n66572 & n66649) | (n66648 & n66649);
  assign n18674 = x128 & x176;
  assign n18675 = x127 & x177;
  assign n18676 = n18674 & n18675;
  assign n18677 = n18674 | n18675;
  assign n18678 = ~n18676 & n18677;
  assign n66651 = n18559 | n18561;
  assign n66656 = (n18559 & n66629) | (n18559 & n66651) | (n66629 & n66651);
  assign n50438 = n18678 & n66656;
  assign n66653 = n18678 & n66651;
  assign n66654 = n18559 & n18678;
  assign n66655 = (n66627 & n66653) | (n66627 & n66654) | (n66653 & n66654);
  assign n66657 = (n50438 & n66578) | (n50438 & n66655) | (n66578 & n66655);
  assign n66658 = (n50438 & n66579) | (n50438 & n66655) | (n66579 & n66655);
  assign n66659 = (n66516 & n66657) | (n66516 & n66658) | (n66657 & n66658);
  assign n50441 = n18678 | n66656;
  assign n66660 = n18678 | n66651;
  assign n66661 = n18559 | n18678;
  assign n66662 = (n66627 & n66660) | (n66627 & n66661) | (n66660 & n66661);
  assign n66663 = (n50441 & n66578) | (n50441 & n66662) | (n66578 & n66662);
  assign n66664 = (n50441 & n66579) | (n50441 & n66662) | (n66579 & n66662);
  assign n66665 = (n66516 & n66663) | (n66516 & n66664) | (n66663 & n66664);
  assign n18681 = ~n66659 & n66665;
  assign n18682 = x126 & x178;
  assign n18683 = n18681 & n18682;
  assign n18684 = n18681 | n18682;
  assign n18685 = ~n18683 & n18684;
  assign n50432 = n18566 | n18568;
  assign n50443 = n18685 & n50432;
  assign n50444 = n18566 & n18685;
  assign n50445 = (n66625 & n50443) | (n66625 & n50444) | (n50443 & n50444);
  assign n50446 = n18685 | n50432;
  assign n50447 = n18566 | n18685;
  assign n50448 = (n66625 & n50446) | (n66625 & n50447) | (n50446 & n50447);
  assign n18688 = ~n50445 & n50448;
  assign n18689 = x125 & x179;
  assign n18690 = n18688 & n18689;
  assign n18691 = n18688 | n18689;
  assign n18692 = ~n18690 & n18691;
  assign n18693 = n66650 & n18692;
  assign n18694 = n66650 | n18692;
  assign n18695 = ~n18693 & n18694;
  assign n18696 = x124 & x180;
  assign n18697 = n18695 & n18696;
  assign n18698 = n18695 | n18696;
  assign n18699 = ~n18697 & n18698;
  assign n50427 = n18580 | n18582;
  assign n50449 = n18699 & n50427;
  assign n50450 = n18580 & n18699;
  assign n50451 = (n66618 & n50449) | (n66618 & n50450) | (n50449 & n50450);
  assign n50452 = n18699 | n50427;
  assign n50453 = n18580 | n18699;
  assign n50454 = (n66618 & n50452) | (n66618 & n50453) | (n50452 & n50453);
  assign n18702 = ~n50451 & n50454;
  assign n18703 = x123 & x181;
  assign n18704 = n18702 & n18703;
  assign n18705 = n18702 | n18703;
  assign n18706 = ~n18704 & n18705;
  assign n50455 = n18587 & n18706;
  assign n66666 = (n18706 & n50399) | (n18706 & n50455) | (n50399 & n50455);
  assign n66667 = (n18589 & n18706) | (n18589 & n50455) | (n18706 & n50455);
  assign n66668 = (n50363 & n66666) | (n50363 & n66667) | (n66666 & n66667);
  assign n50457 = n18587 | n18706;
  assign n66669 = n50399 | n50457;
  assign n66670 = n18589 | n50457;
  assign n66671 = (n50363 & n66669) | (n50363 & n66670) | (n66669 & n66670);
  assign n18709 = ~n66668 & n66671;
  assign n18710 = x122 & x182;
  assign n18711 = n18709 & n18710;
  assign n18712 = n18709 | n18710;
  assign n18713 = ~n18711 & n18712;
  assign n50459 = n18594 & n18713;
  assign n50460 = (n18713 & n50404) | (n18713 & n50459) | (n50404 & n50459);
  assign n50461 = n18594 | n18713;
  assign n50462 = n50404 | n50461;
  assign n18716 = ~n50460 & n50462;
  assign n18717 = x121 & x183;
  assign n18718 = n18716 & n18717;
  assign n18719 = n18716 | n18717;
  assign n18720 = ~n18718 & n18719;
  assign n50463 = n18601 & n18720;
  assign n50464 = (n18720 & n50408) | (n18720 & n50463) | (n50408 & n50463);
  assign n50465 = n18601 | n18720;
  assign n50466 = n50408 | n50465;
  assign n18723 = ~n50464 & n50466;
  assign n18724 = x120 & x184;
  assign n18725 = n18723 & n18724;
  assign n18726 = n18723 | n18724;
  assign n18727 = ~n18725 & n18726;
  assign n50467 = n18608 & n18727;
  assign n50468 = (n18727 & n50413) | (n18727 & n50467) | (n50413 & n50467);
  assign n50469 = n18608 | n18727;
  assign n50470 = n50413 | n50469;
  assign n18730 = ~n50468 & n50470;
  assign n18731 = x119 & x185;
  assign n18732 = n18730 & n18731;
  assign n18733 = n18730 | n18731;
  assign n18734 = ~n18732 & n18733;
  assign n50471 = n18615 & n18734;
  assign n50472 = (n18734 & n50418) | (n18734 & n50471) | (n50418 & n50471);
  assign n50473 = n18615 | n18734;
  assign n50474 = n50418 | n50473;
  assign n18737 = ~n50472 & n50474;
  assign n18738 = x118 & x186;
  assign n18739 = n18737 & n18738;
  assign n18740 = n18737 | n18738;
  assign n18741 = ~n18739 & n18740;
  assign n18742 = n50426 & n18741;
  assign n18743 = n50426 | n18741;
  assign n18744 = ~n18742 & n18743;
  assign n18745 = x117 & x187;
  assign n18746 = n18744 & n18745;
  assign n18747 = n18744 | n18745;
  assign n18748 = ~n18746 & n18747;
  assign n18749 = n18663 & n18748;
  assign n18750 = n18663 | n18748;
  assign n18751 = ~n18749 & n18750;
  assign n18752 = x116 & x188;
  assign n18753 = n18751 & n18752;
  assign n18754 = n18751 | n18752;
  assign n18755 = ~n18753 & n18754;
  assign n18756 = n66645 & n18755;
  assign n18757 = n66645 | n18755;
  assign n18758 = ~n18756 & n18757;
  assign n18759 = x115 & x189;
  assign n18760 = n18758 & n18759;
  assign n18761 = n18758 | n18759;
  assign n18762 = ~n18760 & n18761;
  assign n18763 = n50424 & n18762;
  assign n18764 = n50424 | n18762;
  assign n18765 = ~n18763 & n18764;
  assign n18766 = x114 & x190;
  assign n18767 = n18765 & n18766;
  assign n18768 = n18765 | n18766;
  assign n18769 = ~n18767 & n18768;
  assign n18770 = n50422 & n18769;
  assign n18771 = n50422 | n18769;
  assign n18772 = ~n18770 & n18771;
  assign n18773 = x113 & x191;
  assign n18774 = n18772 & n18773;
  assign n18775 = n18772 | n18773;
  assign n18776 = ~n18774 & n18775;
  assign n18777 = n18657 & n18776;
  assign n18778 = n18657 | n18776;
  assign n18779 = ~n18777 & n18778;
  assign n18780 = x112 & x192;
  assign n18781 = n18779 & n18780;
  assign n18782 = n18779 | n18780;
  assign n18783 = ~n18781 & n18782;
  assign n66672 = n18657 | n18773;
  assign n66673 = (n18657 & n18772) | (n18657 & n66672) | (n18772 & n66672);
  assign n50476 = (n18774 & n18776) | (n18774 & n66673) | (n18776 & n66673);
  assign n50477 = n18767 | n50422;
  assign n50478 = (n18767 & n18769) | (n18767 & n50477) | (n18769 & n50477);
  assign n50479 = n18760 | n50424;
  assign n50480 = (n18760 & n18762) | (n18760 & n50479) | (n18762 & n50479);
  assign n66674 = n18753 | n66645;
  assign n66675 = (n18753 & n18755) | (n18753 & n66674) | (n18755 & n66674);
  assign n50481 = n18746 | n18748;
  assign n50482 = (n18663 & n18746) | (n18663 & n50481) | (n18746 & n50481);
  assign n50483 = n18739 | n18741;
  assign n50484 = (n18739 & n50426) | (n18739 & n50483) | (n50426 & n50483);
  assign n50486 = n18704 | n18706;
  assign n66676 = n18587 | n18704;
  assign n66677 = (n18704 & n18706) | (n18704 & n66676) | (n18706 & n66676);
  assign n66678 = (n50399 & n50486) | (n50399 & n66677) | (n50486 & n66677);
  assign n66679 = (n18589 & n50486) | (n18589 & n66677) | (n50486 & n66677);
  assign n66680 = (n50363 & n66678) | (n50363 & n66679) | (n66678 & n66679);
  assign n18799 = x129 & x176;
  assign n18800 = x128 & x177;
  assign n18801 = n18799 & n18800;
  assign n18802 = n18799 | n18800;
  assign n18803 = ~n18801 & n18802;
  assign n50493 = n18676 & n18803;
  assign n50494 = (n18803 & n66659) | (n18803 & n50493) | (n66659 & n50493);
  assign n50495 = n18676 | n18803;
  assign n50496 = n66659 | n50495;
  assign n18806 = ~n50494 & n50496;
  assign n18807 = x127 & x178;
  assign n18808 = n18806 & n18807;
  assign n18809 = n18806 | n18807;
  assign n18810 = ~n18808 & n18809;
  assign n66681 = n18683 | n18685;
  assign n66682 = (n18683 & n50432) | (n18683 & n66681) | (n50432 & n66681);
  assign n50497 = n18810 & n66682;
  assign n66683 = n18566 | n18683;
  assign n66684 = (n18683 & n18685) | (n18683 & n66683) | (n18685 & n66683);
  assign n50498 = n18810 & n66684;
  assign n50499 = (n66625 & n50497) | (n66625 & n50498) | (n50497 & n50498);
  assign n50500 = n18810 | n66682;
  assign n50501 = n18810 | n66684;
  assign n50502 = (n66625 & n50500) | (n66625 & n50501) | (n50500 & n50501);
  assign n18813 = ~n50499 & n50502;
  assign n18814 = x126 & x179;
  assign n18815 = n18813 & n18814;
  assign n18816 = n18813 | n18814;
  assign n18817 = ~n18815 & n18816;
  assign n50488 = n18690 | n18692;
  assign n50503 = n18817 & n50488;
  assign n50504 = n18690 & n18817;
  assign n50505 = (n66650 & n50503) | (n66650 & n50504) | (n50503 & n50504);
  assign n50506 = n18817 | n50488;
  assign n50507 = n18690 | n18817;
  assign n50508 = (n66650 & n50506) | (n66650 & n50507) | (n50506 & n50507);
  assign n18820 = ~n50505 & n50508;
  assign n18821 = x125 & x180;
  assign n18822 = n18820 & n18821;
  assign n18823 = n18820 | n18821;
  assign n18824 = ~n18822 & n18823;
  assign n50509 = n18697 & n18824;
  assign n66685 = (n18824 & n50450) | (n18824 & n50509) | (n50450 & n50509);
  assign n66686 = (n18824 & n50449) | (n18824 & n50509) | (n50449 & n50509);
  assign n66687 = (n66618 & n66685) | (n66618 & n66686) | (n66685 & n66686);
  assign n50511 = n18697 | n18824;
  assign n66688 = n50450 | n50511;
  assign n66689 = n50449 | n50511;
  assign n66690 = (n66618 & n66688) | (n66618 & n66689) | (n66688 & n66689);
  assign n18827 = ~n66687 & n66690;
  assign n18828 = x124 & x181;
  assign n18829 = n18827 & n18828;
  assign n18830 = n18827 | n18828;
  assign n18831 = ~n18829 & n18830;
  assign n18832 = n66680 & n18831;
  assign n18833 = n66680 | n18831;
  assign n18834 = ~n18832 & n18833;
  assign n18835 = x123 & x182;
  assign n18836 = n18834 & n18835;
  assign n18837 = n18834 | n18835;
  assign n18838 = ~n18836 & n18837;
  assign n50513 = n18711 & n18838;
  assign n50514 = (n18838 & n50460) | (n18838 & n50513) | (n50460 & n50513);
  assign n50515 = n18711 | n18838;
  assign n50516 = n50460 | n50515;
  assign n18841 = ~n50514 & n50516;
  assign n18842 = x122 & x183;
  assign n18843 = n18841 & n18842;
  assign n18844 = n18841 | n18842;
  assign n18845 = ~n18843 & n18844;
  assign n50517 = n18718 & n18845;
  assign n50518 = (n18845 & n50464) | (n18845 & n50517) | (n50464 & n50517);
  assign n50519 = n18718 | n18845;
  assign n50520 = n50464 | n50519;
  assign n18848 = ~n50518 & n50520;
  assign n18849 = x121 & x184;
  assign n18850 = n18848 & n18849;
  assign n18851 = n18848 | n18849;
  assign n18852 = ~n18850 & n18851;
  assign n50521 = n18725 & n18852;
  assign n50522 = (n18852 & n50468) | (n18852 & n50521) | (n50468 & n50521);
  assign n50523 = n18725 | n18852;
  assign n50524 = n50468 | n50523;
  assign n18855 = ~n50522 & n50524;
  assign n18856 = x120 & x185;
  assign n18857 = n18855 & n18856;
  assign n18858 = n18855 | n18856;
  assign n18859 = ~n18857 & n18858;
  assign n50525 = n18732 & n18859;
  assign n50526 = (n18859 & n50472) | (n18859 & n50525) | (n50472 & n50525);
  assign n50527 = n18732 | n18859;
  assign n50528 = n50472 | n50527;
  assign n18862 = ~n50526 & n50528;
  assign n18863 = x119 & x186;
  assign n18864 = n18862 & n18863;
  assign n18865 = n18862 | n18863;
  assign n18866 = ~n18864 & n18865;
  assign n18867 = n50484 & n18866;
  assign n18868 = n50484 | n18866;
  assign n18869 = ~n18867 & n18868;
  assign n18870 = x118 & x187;
  assign n18871 = n18869 & n18870;
  assign n18872 = n18869 | n18870;
  assign n18873 = ~n18871 & n18872;
  assign n18874 = n50482 & n18873;
  assign n18875 = n50482 | n18873;
  assign n18876 = ~n18874 & n18875;
  assign n18877 = x117 & x188;
  assign n18878 = n18876 & n18877;
  assign n18879 = n18876 | n18877;
  assign n18880 = ~n18878 & n18879;
  assign n18881 = n66675 & n18880;
  assign n18882 = n66675 | n18880;
  assign n18883 = ~n18881 & n18882;
  assign n18884 = x116 & x189;
  assign n18885 = n18883 & n18884;
  assign n18886 = n18883 | n18884;
  assign n18887 = ~n18885 & n18886;
  assign n18888 = n50480 & n18887;
  assign n18889 = n50480 | n18887;
  assign n18890 = ~n18888 & n18889;
  assign n18891 = x115 & x190;
  assign n18892 = n18890 & n18891;
  assign n18893 = n18890 | n18891;
  assign n18894 = ~n18892 & n18893;
  assign n18895 = n50478 & n18894;
  assign n18896 = n50478 | n18894;
  assign n18897 = ~n18895 & n18896;
  assign n18898 = x114 & x191;
  assign n18899 = n18897 & n18898;
  assign n18900 = n18897 | n18898;
  assign n18901 = ~n18899 & n18900;
  assign n18902 = n50476 & n18901;
  assign n18903 = n50476 | n18901;
  assign n18904 = ~n18902 & n18903;
  assign n18905 = x113 & x192;
  assign n18906 = n18904 & n18905;
  assign n18907 = n18904 | n18905;
  assign n18908 = ~n18906 & n18907;
  assign n18909 = n18781 & n18908;
  assign n18910 = n18781 | n18908;
  assign n18911 = ~n18909 & n18910;
  assign n18912 = x112 & x193;
  assign n18913 = n18911 & n18912;
  assign n18914 = n18911 | n18912;
  assign n18915 = ~n18913 & n18914;
  assign n50529 = n18781 | n18906;
  assign n50530 = (n18906 & n18908) | (n18906 & n50529) | (n18908 & n50529);
  assign n50531 = n18899 | n50476;
  assign n50532 = (n18899 & n18901) | (n18899 & n50531) | (n18901 & n50531);
  assign n50533 = n18892 | n50478;
  assign n50534 = (n18892 & n18894) | (n18892 & n50533) | (n18894 & n50533);
  assign n50535 = n18885 | n50480;
  assign n50536 = (n18885 & n18887) | (n18885 & n50535) | (n18887 & n50535);
  assign n50537 = n18878 | n18880;
  assign n50538 = (n66675 & n18878) | (n66675 & n50537) | (n18878 & n50537);
  assign n50539 = n18871 | n18873;
  assign n50540 = (n18871 & n50482) | (n18871 & n50539) | (n50482 & n50539);
  assign n50541 = n18864 | n18866;
  assign n50542 = (n18864 & n50484) | (n18864 & n50541) | (n50484 & n50541);
  assign n50546 = n18822 | n18824;
  assign n66691 = n18697 | n18822;
  assign n66692 = (n18822 & n18824) | (n18822 & n66691) | (n18824 & n66691);
  assign n66693 = (n50450 & n50546) | (n50450 & n66692) | (n50546 & n66692);
  assign n66694 = (n50449 & n50546) | (n50449 & n66692) | (n50546 & n66692);
  assign n66695 = (n66618 & n66693) | (n66618 & n66694) | (n66693 & n66694);
  assign n18932 = x130 & x176;
  assign n18933 = x129 & x177;
  assign n18934 = n18932 & n18933;
  assign n18935 = n18932 | n18933;
  assign n18936 = ~n18934 & n18935;
  assign n66700 = n18676 | n18801;
  assign n66701 = (n18801 & n18803) | (n18801 & n66700) | (n18803 & n66700);
  assign n50554 = n18936 & n66701;
  assign n50552 = n18801 | n18803;
  assign n50555 = n18936 & n50552;
  assign n50556 = (n66659 & n50554) | (n66659 & n50555) | (n50554 & n50555);
  assign n50557 = n18936 | n66701;
  assign n50558 = n18936 | n50552;
  assign n50559 = (n66659 & n50557) | (n66659 & n50558) | (n50557 & n50558);
  assign n18939 = ~n50556 & n50559;
  assign n18940 = x128 & x178;
  assign n18941 = n18939 & n18940;
  assign n18942 = n18939 | n18940;
  assign n18943 = ~n18941 & n18942;
  assign n50560 = n18808 & n18943;
  assign n66702 = (n18943 & n50497) | (n18943 & n50560) | (n50497 & n50560);
  assign n66703 = (n18943 & n50498) | (n18943 & n50560) | (n50498 & n50560);
  assign n66704 = (n66625 & n66702) | (n66625 & n66703) | (n66702 & n66703);
  assign n50562 = n18808 | n18943;
  assign n66705 = n50497 | n50562;
  assign n66706 = n50498 | n50562;
  assign n66707 = (n66625 & n66705) | (n66625 & n66706) | (n66705 & n66706);
  assign n18946 = ~n66704 & n66707;
  assign n18947 = x127 & x179;
  assign n18948 = n18946 & n18947;
  assign n18949 = n18946 | n18947;
  assign n18950 = ~n18948 & n18949;
  assign n66696 = n18815 | n18817;
  assign n66697 = (n18815 & n50488) | (n18815 & n66696) | (n50488 & n66696);
  assign n66708 = n18950 & n66697;
  assign n66698 = n18690 | n18815;
  assign n66699 = (n18815 & n18817) | (n18815 & n66698) | (n18817 & n66698);
  assign n66709 = n18950 & n66699;
  assign n66710 = (n66650 & n66708) | (n66650 & n66709) | (n66708 & n66709);
  assign n66711 = n18950 | n66697;
  assign n66712 = n18950 | n66699;
  assign n66713 = (n66650 & n66711) | (n66650 & n66712) | (n66711 & n66712);
  assign n18953 = ~n66710 & n66713;
  assign n18954 = x126 & x180;
  assign n18955 = n18953 & n18954;
  assign n18956 = n18953 | n18954;
  assign n18957 = ~n18955 & n18956;
  assign n18958 = n66695 & n18957;
  assign n18959 = n66695 | n18957;
  assign n18960 = ~n18958 & n18959;
  assign n18961 = x125 & x181;
  assign n18962 = n18960 & n18961;
  assign n18963 = n18960 | n18961;
  assign n18964 = ~n18962 & n18963;
  assign n50543 = n18829 | n18831;
  assign n50564 = n18964 & n50543;
  assign n50565 = n18829 & n18964;
  assign n50566 = (n66680 & n50564) | (n66680 & n50565) | (n50564 & n50565);
  assign n50567 = n18964 | n50543;
  assign n50568 = n18829 | n18964;
  assign n50569 = (n66680 & n50567) | (n66680 & n50568) | (n50567 & n50568);
  assign n18967 = ~n50566 & n50569;
  assign n18968 = x124 & x182;
  assign n18969 = n18967 & n18968;
  assign n18970 = n18967 | n18968;
  assign n18971 = ~n18969 & n18970;
  assign n50570 = n18836 & n18971;
  assign n66714 = (n18971 & n50513) | (n18971 & n50570) | (n50513 & n50570);
  assign n66715 = (n18838 & n18971) | (n18838 & n50570) | (n18971 & n50570);
  assign n66716 = (n50460 & n66714) | (n50460 & n66715) | (n66714 & n66715);
  assign n50572 = n18836 | n18971;
  assign n66717 = n50513 | n50572;
  assign n66718 = n18838 | n50572;
  assign n66719 = (n50460 & n66717) | (n50460 & n66718) | (n66717 & n66718);
  assign n18974 = ~n66716 & n66719;
  assign n18975 = x123 & x183;
  assign n18976 = n18974 & n18975;
  assign n18977 = n18974 | n18975;
  assign n18978 = ~n18976 & n18977;
  assign n50574 = n18843 & n18978;
  assign n50575 = (n18978 & n50518) | (n18978 & n50574) | (n50518 & n50574);
  assign n50576 = n18843 | n18978;
  assign n50577 = n50518 | n50576;
  assign n18981 = ~n50575 & n50577;
  assign n18982 = x122 & x184;
  assign n18983 = n18981 & n18982;
  assign n18984 = n18981 | n18982;
  assign n18985 = ~n18983 & n18984;
  assign n50578 = n18850 & n18985;
  assign n50579 = (n18985 & n50522) | (n18985 & n50578) | (n50522 & n50578);
  assign n50580 = n18850 | n18985;
  assign n50581 = n50522 | n50580;
  assign n18988 = ~n50579 & n50581;
  assign n18989 = x121 & x185;
  assign n18990 = n18988 & n18989;
  assign n18991 = n18988 | n18989;
  assign n18992 = ~n18990 & n18991;
  assign n50582 = n18857 & n18992;
  assign n50583 = (n18992 & n50526) | (n18992 & n50582) | (n50526 & n50582);
  assign n50584 = n18857 | n18992;
  assign n50585 = n50526 | n50584;
  assign n18995 = ~n50583 & n50585;
  assign n18996 = x120 & x186;
  assign n18997 = n18995 & n18996;
  assign n18998 = n18995 | n18996;
  assign n18999 = ~n18997 & n18998;
  assign n19000 = n50542 & n18999;
  assign n19001 = n50542 | n18999;
  assign n19002 = ~n19000 & n19001;
  assign n19003 = x119 & x187;
  assign n19004 = n19002 & n19003;
  assign n19005 = n19002 | n19003;
  assign n19006 = ~n19004 & n19005;
  assign n19007 = n50540 & n19006;
  assign n19008 = n50540 | n19006;
  assign n19009 = ~n19007 & n19008;
  assign n19010 = x118 & x188;
  assign n19011 = n19009 & n19010;
  assign n19012 = n19009 | n19010;
  assign n19013 = ~n19011 & n19012;
  assign n19014 = n50538 & n19013;
  assign n19015 = n50538 | n19013;
  assign n19016 = ~n19014 & n19015;
  assign n19017 = x117 & x189;
  assign n19018 = n19016 & n19017;
  assign n19019 = n19016 | n19017;
  assign n19020 = ~n19018 & n19019;
  assign n19021 = n50536 & n19020;
  assign n19022 = n50536 | n19020;
  assign n19023 = ~n19021 & n19022;
  assign n19024 = x116 & x190;
  assign n19025 = n19023 & n19024;
  assign n19026 = n19023 | n19024;
  assign n19027 = ~n19025 & n19026;
  assign n19028 = n50534 & n19027;
  assign n19029 = n50534 | n19027;
  assign n19030 = ~n19028 & n19029;
  assign n19031 = x115 & x191;
  assign n19032 = n19030 & n19031;
  assign n19033 = n19030 | n19031;
  assign n19034 = ~n19032 & n19033;
  assign n19035 = n50532 & n19034;
  assign n19036 = n50532 | n19034;
  assign n19037 = ~n19035 & n19036;
  assign n19038 = x114 & x192;
  assign n19039 = n19037 & n19038;
  assign n19040 = n19037 | n19038;
  assign n19041 = ~n19039 & n19040;
  assign n19042 = n50530 & n19041;
  assign n19043 = n50530 | n19041;
  assign n19044 = ~n19042 & n19043;
  assign n19045 = x113 & x193;
  assign n19046 = n19044 & n19045;
  assign n19047 = n19044 | n19045;
  assign n19048 = ~n19046 & n19047;
  assign n19049 = n18913 & n19048;
  assign n19050 = n18913 | n19048;
  assign n19051 = ~n19049 & n19050;
  assign n19052 = x112 & x194;
  assign n19053 = n19051 & n19052;
  assign n19054 = n19051 | n19052;
  assign n19055 = ~n19053 & n19054;
  assign n66720 = n18913 | n19045;
  assign n66721 = (n18913 & n19044) | (n18913 & n66720) | (n19044 & n66720);
  assign n50587 = (n19046 & n19048) | (n19046 & n66721) | (n19048 & n66721);
  assign n66722 = n19039 | n50530;
  assign n66723 = (n19039 & n19041) | (n19039 & n66722) | (n19041 & n66722);
  assign n19058 = n19032 | n19035;
  assign n19059 = n19025 | n19028;
  assign n19060 = n19018 | n19021;
  assign n50588 = n19011 | n19013;
  assign n50589 = (n19011 & n50538) | (n19011 & n50588) | (n50538 & n50588);
  assign n50590 = n19004 | n19006;
  assign n50591 = (n19004 & n50540) | (n19004 & n50590) | (n50540 & n50590);
  assign n50592 = n18997 | n18999;
  assign n50593 = (n18997 & n50542) | (n18997 & n50592) | (n50542 & n50592);
  assign n50595 = n18969 | n18971;
  assign n66724 = n18836 | n18969;
  assign n66725 = (n18969 & n18971) | (n18969 & n66724) | (n18971 & n66724);
  assign n66726 = (n50513 & n50595) | (n50513 & n66725) | (n50595 & n66725);
  assign n66727 = (n18838 & n50595) | (n18838 & n66725) | (n50595 & n66725);
  assign n66728 = (n50460 & n66726) | (n50460 & n66727) | (n66726 & n66727);
  assign n19073 = x131 & x176;
  assign n19074 = x130 & x177;
  assign n19075 = n19073 & n19074;
  assign n19076 = n19073 | n19074;
  assign n19077 = ~n19075 & n19076;
  assign n66729 = n18934 | n18936;
  assign n66730 = (n18934 & n66701) | (n18934 & n66729) | (n66701 & n66729);
  assign n50607 = n19077 & n66730;
  assign n66731 = (n18934 & n50552) | (n18934 & n66729) | (n50552 & n66729);
  assign n50608 = n19077 & n66731;
  assign n50609 = (n66659 & n50607) | (n66659 & n50608) | (n50607 & n50608);
  assign n50610 = n19077 | n66730;
  assign n50611 = n19077 | n66731;
  assign n50612 = (n66659 & n50610) | (n66659 & n50611) | (n50610 & n50611);
  assign n19080 = ~n50609 & n50612;
  assign n19081 = x129 & x178;
  assign n19082 = n19080 & n19081;
  assign n19083 = n19080 | n19081;
  assign n19084 = ~n19082 & n19083;
  assign n66732 = n18808 | n18941;
  assign n66733 = (n18941 & n18943) | (n18941 & n66732) | (n18943 & n66732);
  assign n50613 = n19084 & n66733;
  assign n50602 = n18941 | n18943;
  assign n50614 = n19084 & n50602;
  assign n66734 = (n50497 & n50613) | (n50497 & n50614) | (n50613 & n50614);
  assign n66735 = (n50498 & n50613) | (n50498 & n50614) | (n50613 & n50614);
  assign n66736 = (n66625 & n66734) | (n66625 & n66735) | (n66734 & n66735);
  assign n50616 = n19084 | n66733;
  assign n50617 = n19084 | n50602;
  assign n66737 = (n50497 & n50616) | (n50497 & n50617) | (n50616 & n50617);
  assign n66738 = (n50498 & n50616) | (n50498 & n50617) | (n50616 & n50617);
  assign n66739 = (n66625 & n66737) | (n66625 & n66738) | (n66737 & n66738);
  assign n19087 = ~n66736 & n66739;
  assign n19088 = x128 & x179;
  assign n19089 = n19087 & n19088;
  assign n19090 = n19087 | n19088;
  assign n19091 = ~n19089 & n19090;
  assign n50599 = n18948 | n18950;
  assign n50619 = n19091 & n50599;
  assign n50620 = n18948 & n19091;
  assign n66740 = (n50619 & n50620) | (n50619 & n66697) | (n50620 & n66697);
  assign n66741 = (n50619 & n50620) | (n50619 & n66699) | (n50620 & n66699);
  assign n66742 = (n66650 & n66740) | (n66650 & n66741) | (n66740 & n66741);
  assign n50622 = n19091 | n50599;
  assign n50623 = n18948 | n19091;
  assign n66743 = (n50622 & n50623) | (n50622 & n66697) | (n50623 & n66697);
  assign n66744 = (n50622 & n50623) | (n50622 & n66699) | (n50623 & n66699);
  assign n66745 = (n66650 & n66743) | (n66650 & n66744) | (n66743 & n66744);
  assign n19094 = ~n66742 & n66745;
  assign n19095 = x127 & x180;
  assign n19096 = n19094 & n19095;
  assign n19097 = n19094 | n19095;
  assign n19098 = ~n19096 & n19097;
  assign n50597 = n18955 | n18957;
  assign n50625 = n19098 & n50597;
  assign n50626 = n18955 & n19098;
  assign n50627 = (n66695 & n50625) | (n66695 & n50626) | (n50625 & n50626);
  assign n50628 = n19098 | n50597;
  assign n50629 = n18955 | n19098;
  assign n50630 = (n66695 & n50628) | (n66695 & n50629) | (n50628 & n50629);
  assign n19101 = ~n50627 & n50630;
  assign n19102 = x126 & x181;
  assign n19103 = n19101 & n19102;
  assign n19104 = n19101 | n19102;
  assign n19105 = ~n19103 & n19104;
  assign n50631 = n18962 & n19105;
  assign n66746 = (n19105 & n50565) | (n19105 & n50631) | (n50565 & n50631);
  assign n66747 = (n19105 & n50564) | (n19105 & n50631) | (n50564 & n50631);
  assign n66748 = (n66680 & n66746) | (n66680 & n66747) | (n66746 & n66747);
  assign n50633 = n18962 | n19105;
  assign n66749 = n50565 | n50633;
  assign n66750 = n50564 | n50633;
  assign n66751 = (n66680 & n66749) | (n66680 & n66750) | (n66749 & n66750);
  assign n19108 = ~n66748 & n66751;
  assign n19109 = x125 & x182;
  assign n19110 = n19108 & n19109;
  assign n19111 = n19108 | n19109;
  assign n19112 = ~n19110 & n19111;
  assign n19113 = n66728 & n19112;
  assign n19114 = n66728 | n19112;
  assign n19115 = ~n19113 & n19114;
  assign n19116 = x124 & x183;
  assign n19117 = n19115 & n19116;
  assign n19118 = n19115 | n19116;
  assign n19119 = ~n19117 & n19118;
  assign n50635 = n18976 & n19119;
  assign n50636 = (n19119 & n50575) | (n19119 & n50635) | (n50575 & n50635);
  assign n50637 = n18976 | n19119;
  assign n50638 = n50575 | n50637;
  assign n19122 = ~n50636 & n50638;
  assign n19123 = x123 & x184;
  assign n19124 = n19122 & n19123;
  assign n19125 = n19122 | n19123;
  assign n19126 = ~n19124 & n19125;
  assign n50639 = n18983 & n19126;
  assign n50640 = (n19126 & n50579) | (n19126 & n50639) | (n50579 & n50639);
  assign n50641 = n18983 | n19126;
  assign n50642 = n50579 | n50641;
  assign n19129 = ~n50640 & n50642;
  assign n19130 = x122 & x185;
  assign n19131 = n19129 & n19130;
  assign n19132 = n19129 | n19130;
  assign n19133 = ~n19131 & n19132;
  assign n50643 = n18990 & n19133;
  assign n50644 = (n19133 & n50583) | (n19133 & n50643) | (n50583 & n50643);
  assign n50645 = n18990 | n19133;
  assign n50646 = n50583 | n50645;
  assign n19136 = ~n50644 & n50646;
  assign n19137 = x121 & x186;
  assign n19138 = n19136 & n19137;
  assign n19139 = n19136 | n19137;
  assign n19140 = ~n19138 & n19139;
  assign n19141 = n50593 & n19140;
  assign n19142 = n50593 | n19140;
  assign n19143 = ~n19141 & n19142;
  assign n19144 = x120 & x187;
  assign n19145 = n19143 & n19144;
  assign n19146 = n19143 | n19144;
  assign n19147 = ~n19145 & n19146;
  assign n19148 = n50591 & n19147;
  assign n19149 = n50591 | n19147;
  assign n19150 = ~n19148 & n19149;
  assign n19151 = x119 & x188;
  assign n19152 = n19150 & n19151;
  assign n19153 = n19150 | n19151;
  assign n19154 = ~n19152 & n19153;
  assign n19155 = n50589 & n19154;
  assign n19156 = n50589 | n19154;
  assign n19157 = ~n19155 & n19156;
  assign n19158 = x118 & x189;
  assign n19159 = n19157 & n19158;
  assign n19160 = n19157 | n19158;
  assign n19161 = ~n19159 & n19160;
  assign n19162 = n19060 & n19161;
  assign n19163 = n19060 | n19161;
  assign n19164 = ~n19162 & n19163;
  assign n19165 = x117 & x190;
  assign n19166 = n19164 & n19165;
  assign n19167 = n19164 | n19165;
  assign n19168 = ~n19166 & n19167;
  assign n19169 = n19059 & n19168;
  assign n19170 = n19059 | n19168;
  assign n19171 = ~n19169 & n19170;
  assign n19172 = x116 & x191;
  assign n19173 = n19171 & n19172;
  assign n19174 = n19171 | n19172;
  assign n19175 = ~n19173 & n19174;
  assign n19176 = n19058 & n19175;
  assign n19177 = n19058 | n19175;
  assign n19178 = ~n19176 & n19177;
  assign n19179 = x115 & x192;
  assign n19180 = n19178 & n19179;
  assign n19181 = n19178 | n19179;
  assign n19182 = ~n19180 & n19181;
  assign n19183 = n66723 & n19182;
  assign n19184 = n66723 | n19182;
  assign n19185 = ~n19183 & n19184;
  assign n19186 = x114 & x193;
  assign n19187 = n19185 & n19186;
  assign n19188 = n19185 | n19186;
  assign n19189 = ~n19187 & n19188;
  assign n19190 = n50587 & n19189;
  assign n19191 = n50587 | n19189;
  assign n19192 = ~n19190 & n19191;
  assign n19193 = x113 & x194;
  assign n19194 = n19192 & n19193;
  assign n19195 = n19192 | n19193;
  assign n19196 = ~n19194 & n19195;
  assign n19197 = n19053 & n19196;
  assign n19198 = n19053 | n19196;
  assign n19199 = ~n19197 & n19198;
  assign n19200 = x112 & x195;
  assign n19201 = n19199 & n19200;
  assign n19202 = n19199 | n19200;
  assign n19203 = ~n19201 & n19202;
  assign n66752 = n19053 | n19193;
  assign n66753 = (n19053 & n19192) | (n19053 & n66752) | (n19192 & n66752);
  assign n50648 = (n19194 & n19196) | (n19194 & n66753) | (n19196 & n66753);
  assign n50649 = n19187 | n50587;
  assign n50650 = (n19187 & n19189) | (n19187 & n50649) | (n19189 & n50649);
  assign n66754 = n19180 | n66723;
  assign n66755 = (n19180 & n19182) | (n19180 & n66754) | (n19182 & n66754);
  assign n19207 = n19173 | n19176;
  assign n19208 = n19166 | n19169;
  assign n50651 = n19159 | n19161;
  assign n50652 = (n19060 & n19159) | (n19060 & n50651) | (n19159 & n50651);
  assign n50653 = n19152 | n19154;
  assign n50654 = (n19152 & n50589) | (n19152 & n50653) | (n50589 & n50653);
  assign n50655 = n19145 | n19147;
  assign n50656 = (n19145 & n50591) | (n19145 & n50655) | (n50591 & n50655);
  assign n50657 = n19138 | n19140;
  assign n50658 = (n19138 & n50593) | (n19138 & n50657) | (n50593 & n50657);
  assign n50662 = n19103 | n19105;
  assign n66756 = n18962 | n19103;
  assign n66757 = (n19103 & n19105) | (n19103 & n66756) | (n19105 & n66756);
  assign n66758 = (n50565 & n50662) | (n50565 & n66757) | (n50662 & n66757);
  assign n66759 = (n50564 & n50662) | (n50564 & n66757) | (n50662 & n66757);
  assign n66760 = (n66680 & n66758) | (n66680 & n66759) | (n66758 & n66759);
  assign n66761 = n19089 | n19091;
  assign n66762 = (n19089 & n50599) | (n19089 & n66761) | (n50599 & n66761);
  assign n66763 = n18948 | n19089;
  assign n66764 = (n19089 & n19091) | (n19089 & n66763) | (n19091 & n66763);
  assign n66765 = (n66697 & n66762) | (n66697 & n66764) | (n66762 & n66764);
  assign n66766 = (n66699 & n66762) | (n66699 & n66764) | (n66762 & n66764);
  assign n66767 = (n66650 & n66765) | (n66650 & n66766) | (n66765 & n66766);
  assign n66768 = n19082 | n19084;
  assign n66769 = (n19082 & n66733) | (n19082 & n66768) | (n66733 & n66768);
  assign n66770 = (n19082 & n50602) | (n19082 & n66768) | (n50602 & n66768);
  assign n66771 = (n50497 & n66769) | (n50497 & n66770) | (n66769 & n66770);
  assign n66772 = (n50498 & n66769) | (n50498 & n66770) | (n66769 & n66770);
  assign n66773 = (n66625 & n66771) | (n66625 & n66772) | (n66771 & n66772);
  assign n19222 = x132 & x176;
  assign n19223 = x131 & x177;
  assign n19224 = n19222 & n19223;
  assign n19225 = n19222 | n19223;
  assign n19226 = ~n19224 & n19225;
  assign n66774 = n19075 | n19077;
  assign n66776 = n19226 & n66774;
  assign n66777 = n19075 & n19226;
  assign n66778 = (n66730 & n66776) | (n66730 & n66777) | (n66776 & n66777);
  assign n66780 = (n66731 & n66776) | (n66731 & n66777) | (n66776 & n66777);
  assign n50675 = (n66659 & n66778) | (n66659 & n66780) | (n66778 & n66780);
  assign n66781 = n19226 | n66774;
  assign n66782 = n19075 | n19226;
  assign n66783 = (n66730 & n66781) | (n66730 & n66782) | (n66781 & n66782);
  assign n66784 = (n66731 & n66781) | (n66731 & n66782) | (n66781 & n66782);
  assign n50678 = (n66659 & n66783) | (n66659 & n66784) | (n66783 & n66784);
  assign n19229 = ~n50675 & n50678;
  assign n19230 = x130 & x178;
  assign n19231 = n19229 & n19230;
  assign n19232 = n19229 | n19230;
  assign n19233 = ~n19231 & n19232;
  assign n19234 = n66773 & n19233;
  assign n19235 = n66773 | n19233;
  assign n19236 = ~n19234 & n19235;
  assign n19237 = x129 & x179;
  assign n19238 = n19236 & n19237;
  assign n19239 = n19236 | n19237;
  assign n19240 = ~n19238 & n19239;
  assign n19241 = n66767 & n19240;
  assign n19242 = n66767 | n19240;
  assign n19243 = ~n19241 & n19242;
  assign n19244 = x128 & x180;
  assign n19245 = n19243 & n19244;
  assign n19246 = n19243 | n19244;
  assign n19247 = ~n19245 & n19246;
  assign n50679 = n19096 & n19247;
  assign n66785 = (n19247 & n50625) | (n19247 & n50679) | (n50625 & n50679);
  assign n66786 = (n19247 & n50626) | (n19247 & n50679) | (n50626 & n50679);
  assign n66787 = (n66695 & n66785) | (n66695 & n66786) | (n66785 & n66786);
  assign n50681 = n19096 | n19247;
  assign n66788 = n50625 | n50681;
  assign n66789 = n50626 | n50681;
  assign n66790 = (n66695 & n66788) | (n66695 & n66789) | (n66788 & n66789);
  assign n19250 = ~n66787 & n66790;
  assign n19251 = x127 & x181;
  assign n19252 = n19250 & n19251;
  assign n19253 = n19250 | n19251;
  assign n19254 = ~n19252 & n19253;
  assign n19255 = n66760 & n19254;
  assign n19256 = n66760 | n19254;
  assign n19257 = ~n19255 & n19256;
  assign n19258 = x126 & x182;
  assign n19259 = n19257 & n19258;
  assign n19260 = n19257 | n19258;
  assign n19261 = ~n19259 & n19260;
  assign n50659 = n19110 | n19112;
  assign n50683 = n19261 & n50659;
  assign n50684 = n19110 & n19261;
  assign n50685 = (n66728 & n50683) | (n66728 & n50684) | (n50683 & n50684);
  assign n50686 = n19261 | n50659;
  assign n50687 = n19110 | n19261;
  assign n50688 = (n66728 & n50686) | (n66728 & n50687) | (n50686 & n50687);
  assign n19264 = ~n50685 & n50688;
  assign n19265 = x125 & x183;
  assign n19266 = n19264 & n19265;
  assign n19267 = n19264 | n19265;
  assign n19268 = ~n19266 & n19267;
  assign n50689 = n19117 & n19268;
  assign n66791 = (n19268 & n50635) | (n19268 & n50689) | (n50635 & n50689);
  assign n66792 = (n19119 & n19268) | (n19119 & n50689) | (n19268 & n50689);
  assign n66793 = (n50575 & n66791) | (n50575 & n66792) | (n66791 & n66792);
  assign n50691 = n19117 | n19268;
  assign n66794 = n50635 | n50691;
  assign n66795 = n19119 | n50691;
  assign n66796 = (n50575 & n66794) | (n50575 & n66795) | (n66794 & n66795);
  assign n19271 = ~n66793 & n66796;
  assign n19272 = x124 & x184;
  assign n19273 = n19271 & n19272;
  assign n19274 = n19271 | n19272;
  assign n19275 = ~n19273 & n19274;
  assign n50693 = n19124 & n19275;
  assign n50694 = (n19275 & n50640) | (n19275 & n50693) | (n50640 & n50693);
  assign n50695 = n19124 | n19275;
  assign n50696 = n50640 | n50695;
  assign n19278 = ~n50694 & n50696;
  assign n19279 = x123 & x185;
  assign n19280 = n19278 & n19279;
  assign n19281 = n19278 | n19279;
  assign n19282 = ~n19280 & n19281;
  assign n50697 = n19131 & n19282;
  assign n50698 = (n19282 & n50644) | (n19282 & n50697) | (n50644 & n50697);
  assign n50699 = n19131 | n19282;
  assign n50700 = n50644 | n50699;
  assign n19285 = ~n50698 & n50700;
  assign n19286 = x122 & x186;
  assign n19287 = n19285 & n19286;
  assign n19288 = n19285 | n19286;
  assign n19289 = ~n19287 & n19288;
  assign n19290 = n50658 & n19289;
  assign n19291 = n50658 | n19289;
  assign n19292 = ~n19290 & n19291;
  assign n19293 = x121 & x187;
  assign n19294 = n19292 & n19293;
  assign n19295 = n19292 | n19293;
  assign n19296 = ~n19294 & n19295;
  assign n19297 = n50656 & n19296;
  assign n19298 = n50656 | n19296;
  assign n19299 = ~n19297 & n19298;
  assign n19300 = x120 & x188;
  assign n19301 = n19299 & n19300;
  assign n19302 = n19299 | n19300;
  assign n19303 = ~n19301 & n19302;
  assign n19304 = n50654 & n19303;
  assign n19305 = n50654 | n19303;
  assign n19306 = ~n19304 & n19305;
  assign n19307 = x119 & x189;
  assign n19308 = n19306 & n19307;
  assign n19309 = n19306 | n19307;
  assign n19310 = ~n19308 & n19309;
  assign n19311 = n50652 & n19310;
  assign n19312 = n50652 | n19310;
  assign n19313 = ~n19311 & n19312;
  assign n19314 = x118 & x190;
  assign n19315 = n19313 & n19314;
  assign n19316 = n19313 | n19314;
  assign n19317 = ~n19315 & n19316;
  assign n19318 = n19208 & n19317;
  assign n19319 = n19208 | n19317;
  assign n19320 = ~n19318 & n19319;
  assign n19321 = x117 & x191;
  assign n19322 = n19320 & n19321;
  assign n19323 = n19320 | n19321;
  assign n19324 = ~n19322 & n19323;
  assign n19325 = n19207 & n19324;
  assign n19326 = n19207 | n19324;
  assign n19327 = ~n19325 & n19326;
  assign n19328 = x116 & x192;
  assign n19329 = n19327 & n19328;
  assign n19330 = n19327 | n19328;
  assign n19331 = ~n19329 & n19330;
  assign n19332 = n66755 & n19331;
  assign n19333 = n66755 | n19331;
  assign n19334 = ~n19332 & n19333;
  assign n19335 = x115 & x193;
  assign n19336 = n19334 & n19335;
  assign n19337 = n19334 | n19335;
  assign n19338 = ~n19336 & n19337;
  assign n19339 = n50650 & n19338;
  assign n19340 = n50650 | n19338;
  assign n19341 = ~n19339 & n19340;
  assign n19342 = x114 & x194;
  assign n19343 = n19341 & n19342;
  assign n19344 = n19341 | n19342;
  assign n19345 = ~n19343 & n19344;
  assign n19346 = n50648 & n19345;
  assign n19347 = n50648 | n19345;
  assign n19348 = ~n19346 & n19347;
  assign n19349 = x113 & x195;
  assign n19350 = n19348 & n19349;
  assign n19351 = n19348 | n19349;
  assign n19352 = ~n19350 & n19351;
  assign n19353 = n19201 & n19352;
  assign n19354 = n19201 | n19352;
  assign n19355 = ~n19353 & n19354;
  assign n19356 = x112 & x196;
  assign n19357 = n19355 & n19356;
  assign n19358 = n19355 | n19356;
  assign n19359 = ~n19357 & n19358;
  assign n66797 = n19201 | n19349;
  assign n66798 = (n19201 & n19348) | (n19201 & n66797) | (n19348 & n66797);
  assign n50702 = (n19350 & n19352) | (n19350 & n66798) | (n19352 & n66798);
  assign n50703 = n19343 | n50648;
  assign n50704 = (n19343 & n19345) | (n19343 & n50703) | (n19345 & n50703);
  assign n50705 = n19336 | n50650;
  assign n50706 = (n19336 & n19338) | (n19336 & n50705) | (n19338 & n50705);
  assign n66799 = n19329 | n66755;
  assign n66800 = (n19329 & n19331) | (n19329 & n66799) | (n19331 & n66799);
  assign n19364 = n19322 | n19325;
  assign n50707 = n19315 | n19317;
  assign n50708 = (n19208 & n19315) | (n19208 & n50707) | (n19315 & n50707);
  assign n50709 = n19308 | n19310;
  assign n50710 = (n19308 & n50652) | (n19308 & n50709) | (n50652 & n50709);
  assign n50711 = n19301 | n19303;
  assign n50712 = (n19301 & n50654) | (n19301 & n50711) | (n50654 & n50711);
  assign n50713 = n19294 | n19296;
  assign n50714 = (n19294 & n50656) | (n19294 & n50713) | (n50656 & n50713);
  assign n50715 = n19287 | n19289;
  assign n50716 = (n19287 & n50658) | (n19287 & n50715) | (n50658 & n50715);
  assign n50718 = n19266 | n19268;
  assign n66801 = n19117 | n19266;
  assign n66802 = (n19266 & n19268) | (n19266 & n66801) | (n19268 & n66801);
  assign n66803 = (n50635 & n50718) | (n50635 & n66802) | (n50718 & n66802);
  assign n66804 = (n19119 & n50718) | (n19119 & n66802) | (n50718 & n66802);
  assign n66805 = (n50575 & n66803) | (n50575 & n66804) | (n66803 & n66804);
  assign n50723 = n19245 | n19247;
  assign n66806 = n19096 | n19245;
  assign n66807 = (n19245 & n19247) | (n19245 & n66806) | (n19247 & n66806);
  assign n66808 = (n50625 & n50723) | (n50625 & n66807) | (n50723 & n66807);
  assign n66809 = (n50626 & n50723) | (n50626 & n66807) | (n50723 & n66807);
  assign n66810 = (n66695 & n66808) | (n66695 & n66809) | (n66808 & n66809);
  assign n19379 = x133 & x176;
  assign n19380 = x132 & x177;
  assign n19381 = n19379 & n19380;
  assign n19382 = n19379 | n19380;
  assign n19383 = ~n19381 & n19382;
  assign n50729 = n19224 & n19383;
  assign n66811 = (n19383 & n50729) | (n19383 & n66780) | (n50729 & n66780);
  assign n66812 = (n19383 & n50729) | (n19383 & n66778) | (n50729 & n66778);
  assign n66813 = (n66659 & n66811) | (n66659 & n66812) | (n66811 & n66812);
  assign n50731 = n19224 | n19383;
  assign n66814 = n50731 | n66780;
  assign n66815 = n50731 | n66778;
  assign n66816 = (n66659 & n66814) | (n66659 & n66815) | (n66814 & n66815);
  assign n19386 = ~n66813 & n66816;
  assign n19387 = x131 & x178;
  assign n19388 = n19386 & n19387;
  assign n19389 = n19386 | n19387;
  assign n19390 = ~n19388 & n19389;
  assign n50727 = n19231 | n19233;
  assign n50733 = n19390 & n50727;
  assign n50734 = n19231 & n19390;
  assign n50735 = (n66773 & n50733) | (n66773 & n50734) | (n50733 & n50734);
  assign n50736 = n19390 | n50727;
  assign n50737 = n19231 | n19390;
  assign n50738 = (n66773 & n50736) | (n66773 & n50737) | (n50736 & n50737);
  assign n19393 = ~n50735 & n50738;
  assign n19394 = x130 & x179;
  assign n19395 = n19393 & n19394;
  assign n19396 = n19393 | n19394;
  assign n19397 = ~n19395 & n19396;
  assign n50725 = n19238 | n19240;
  assign n50739 = n19397 & n50725;
  assign n50740 = n19238 & n19397;
  assign n50741 = (n66767 & n50739) | (n66767 & n50740) | (n50739 & n50740);
  assign n50742 = n19397 | n50725;
  assign n50743 = n19238 | n19397;
  assign n50744 = (n66767 & n50742) | (n66767 & n50743) | (n50742 & n50743);
  assign n19400 = ~n50741 & n50744;
  assign n19401 = x129 & x180;
  assign n19402 = n19400 & n19401;
  assign n19403 = n19400 | n19401;
  assign n19404 = ~n19402 & n19403;
  assign n19405 = n66810 & n19404;
  assign n19406 = n66810 | n19404;
  assign n19407 = ~n19405 & n19406;
  assign n19408 = x128 & x181;
  assign n19409 = n19407 & n19408;
  assign n19410 = n19407 | n19408;
  assign n19411 = ~n19409 & n19410;
  assign n50720 = n19252 | n19254;
  assign n50745 = n19411 & n50720;
  assign n50746 = n19252 & n19411;
  assign n50747 = (n66760 & n50745) | (n66760 & n50746) | (n50745 & n50746);
  assign n50748 = n19411 | n50720;
  assign n50749 = n19252 | n19411;
  assign n50750 = (n66760 & n50748) | (n66760 & n50749) | (n50748 & n50749);
  assign n19414 = ~n50747 & n50750;
  assign n19415 = x127 & x182;
  assign n19416 = n19414 & n19415;
  assign n19417 = n19414 | n19415;
  assign n19418 = ~n19416 & n19417;
  assign n50751 = n19259 & n19418;
  assign n66817 = (n19418 & n50684) | (n19418 & n50751) | (n50684 & n50751);
  assign n66818 = (n19418 & n50683) | (n19418 & n50751) | (n50683 & n50751);
  assign n66819 = (n66728 & n66817) | (n66728 & n66818) | (n66817 & n66818);
  assign n50753 = n19259 | n19418;
  assign n66820 = n50684 | n50753;
  assign n66821 = n50683 | n50753;
  assign n66822 = (n66728 & n66820) | (n66728 & n66821) | (n66820 & n66821);
  assign n19421 = ~n66819 & n66822;
  assign n19422 = x126 & x183;
  assign n19423 = n19421 & n19422;
  assign n19424 = n19421 | n19422;
  assign n19425 = ~n19423 & n19424;
  assign n19426 = n66805 & n19425;
  assign n19427 = n66805 | n19425;
  assign n19428 = ~n19426 & n19427;
  assign n19429 = x125 & x184;
  assign n19430 = n19428 & n19429;
  assign n19431 = n19428 | n19429;
  assign n19432 = ~n19430 & n19431;
  assign n50755 = n19273 & n19432;
  assign n50756 = (n19432 & n50694) | (n19432 & n50755) | (n50694 & n50755);
  assign n50757 = n19273 | n19432;
  assign n50758 = n50694 | n50757;
  assign n19435 = ~n50756 & n50758;
  assign n19436 = x124 & x185;
  assign n19437 = n19435 & n19436;
  assign n19438 = n19435 | n19436;
  assign n19439 = ~n19437 & n19438;
  assign n50759 = n19280 & n19439;
  assign n50760 = (n19439 & n50698) | (n19439 & n50759) | (n50698 & n50759);
  assign n50761 = n19280 | n19439;
  assign n50762 = n50698 | n50761;
  assign n19442 = ~n50760 & n50762;
  assign n19443 = x123 & x186;
  assign n19444 = n19442 & n19443;
  assign n19445 = n19442 | n19443;
  assign n19446 = ~n19444 & n19445;
  assign n19447 = n50716 & n19446;
  assign n19448 = n50716 | n19446;
  assign n19449 = ~n19447 & n19448;
  assign n19450 = x122 & x187;
  assign n19451 = n19449 & n19450;
  assign n19452 = n19449 | n19450;
  assign n19453 = ~n19451 & n19452;
  assign n19454 = n50714 & n19453;
  assign n19455 = n50714 | n19453;
  assign n19456 = ~n19454 & n19455;
  assign n19457 = x121 & x188;
  assign n19458 = n19456 & n19457;
  assign n19459 = n19456 | n19457;
  assign n19460 = ~n19458 & n19459;
  assign n19461 = n50712 & n19460;
  assign n19462 = n50712 | n19460;
  assign n19463 = ~n19461 & n19462;
  assign n19464 = x120 & x189;
  assign n19465 = n19463 & n19464;
  assign n19466 = n19463 | n19464;
  assign n19467 = ~n19465 & n19466;
  assign n19468 = n50710 & n19467;
  assign n19469 = n50710 | n19467;
  assign n19470 = ~n19468 & n19469;
  assign n19471 = x119 & x190;
  assign n19472 = n19470 & n19471;
  assign n19473 = n19470 | n19471;
  assign n19474 = ~n19472 & n19473;
  assign n19475 = n50708 & n19474;
  assign n19476 = n50708 | n19474;
  assign n19477 = ~n19475 & n19476;
  assign n19478 = x118 & x191;
  assign n19479 = n19477 & n19478;
  assign n19480 = n19477 | n19478;
  assign n19481 = ~n19479 & n19480;
  assign n19482 = n19364 & n19481;
  assign n19483 = n19364 | n19481;
  assign n19484 = ~n19482 & n19483;
  assign n19485 = x117 & x192;
  assign n19486 = n19484 & n19485;
  assign n19487 = n19484 | n19485;
  assign n19488 = ~n19486 & n19487;
  assign n19489 = n66800 & n19488;
  assign n19490 = n66800 | n19488;
  assign n19491 = ~n19489 & n19490;
  assign n19492 = x116 & x193;
  assign n19493 = n19491 & n19492;
  assign n19494 = n19491 | n19492;
  assign n19495 = ~n19493 & n19494;
  assign n19496 = n50706 & n19495;
  assign n19497 = n50706 | n19495;
  assign n19498 = ~n19496 & n19497;
  assign n19499 = x115 & x194;
  assign n19500 = n19498 & n19499;
  assign n19501 = n19498 | n19499;
  assign n19502 = ~n19500 & n19501;
  assign n19503 = n50704 & n19502;
  assign n19504 = n50704 | n19502;
  assign n19505 = ~n19503 & n19504;
  assign n19506 = x114 & x195;
  assign n19507 = n19505 & n19506;
  assign n19508 = n19505 | n19506;
  assign n19509 = ~n19507 & n19508;
  assign n19510 = n50702 & n19509;
  assign n19511 = n50702 | n19509;
  assign n19512 = ~n19510 & n19511;
  assign n19513 = x113 & x196;
  assign n19514 = n19512 & n19513;
  assign n19515 = n19512 | n19513;
  assign n19516 = ~n19514 & n19515;
  assign n19517 = n19357 & n19516;
  assign n19518 = n19357 | n19516;
  assign n19519 = ~n19517 & n19518;
  assign n19520 = x112 & x197;
  assign n19521 = n19519 & n19520;
  assign n19522 = n19519 | n19520;
  assign n19523 = ~n19521 & n19522;
  assign n66823 = n19357 | n19513;
  assign n66824 = (n19357 & n19512) | (n19357 & n66823) | (n19512 & n66823);
  assign n50764 = (n19514 & n19516) | (n19514 & n66824) | (n19516 & n66824);
  assign n50765 = n19507 | n50702;
  assign n50766 = (n19507 & n19509) | (n19507 & n50765) | (n19509 & n50765);
  assign n50767 = n19500 | n50704;
  assign n50768 = (n19500 & n19502) | (n19500 & n50767) | (n19502 & n50767);
  assign n50769 = n19493 | n50706;
  assign n50770 = (n19493 & n19495) | (n19493 & n50769) | (n19495 & n50769);
  assign n66825 = n19486 | n66800;
  assign n66826 = (n19486 & n19488) | (n19486 & n66825) | (n19488 & n66825);
  assign n50771 = n19479 | n19481;
  assign n50772 = (n19364 & n19479) | (n19364 & n50771) | (n19479 & n50771);
  assign n50773 = n19472 | n19474;
  assign n50774 = (n19472 & n50708) | (n19472 & n50773) | (n50708 & n50773);
  assign n50775 = n19465 | n19467;
  assign n50776 = (n19465 & n50710) | (n19465 & n50775) | (n50710 & n50775);
  assign n50777 = n19458 | n19460;
  assign n50778 = (n19458 & n50712) | (n19458 & n50777) | (n50712 & n50777);
  assign n50779 = n19451 | n19453;
  assign n50780 = (n19451 & n50714) | (n19451 & n50779) | (n50714 & n50779);
  assign n50781 = n19444 | n19446;
  assign n50782 = (n19444 & n50716) | (n19444 & n50781) | (n50716 & n50781);
  assign n50786 = n19416 | n19418;
  assign n66827 = n19259 | n19416;
  assign n66828 = (n19416 & n19418) | (n19416 & n66827) | (n19418 & n66827);
  assign n66829 = (n50684 & n50786) | (n50684 & n66828) | (n50786 & n66828);
  assign n66830 = (n50683 & n50786) | (n50683 & n66828) | (n50786 & n66828);
  assign n66831 = (n66728 & n66829) | (n66728 & n66830) | (n66829 & n66830);
  assign n19544 = x134 & x176;
  assign n19545 = x133 & x177;
  assign n19546 = n19544 & n19545;
  assign n19547 = n19544 | n19545;
  assign n19548 = ~n19546 & n19547;
  assign n66836 = n19224 | n19381;
  assign n66837 = (n19381 & n19383) | (n19381 & n66836) | (n19383 & n66836);
  assign n50799 = n19548 & n66837;
  assign n50797 = n19381 | n19383;
  assign n50800 = n19548 & n50797;
  assign n66838 = (n50799 & n50800) | (n50799 & n66780) | (n50800 & n66780);
  assign n66839 = (n50799 & n50800) | (n50799 & n66778) | (n50800 & n66778);
  assign n66840 = (n66659 & n66838) | (n66659 & n66839) | (n66838 & n66839);
  assign n50802 = n19548 | n66837;
  assign n50803 = n19548 | n50797;
  assign n66841 = (n50802 & n50803) | (n50802 & n66780) | (n50803 & n66780);
  assign n66842 = (n50802 & n50803) | (n50802 & n66778) | (n50803 & n66778);
  assign n66843 = (n66659 & n66841) | (n66659 & n66842) | (n66841 & n66842);
  assign n19551 = ~n66840 & n66843;
  assign n19552 = x132 & x178;
  assign n19553 = n19551 & n19552;
  assign n19554 = n19551 | n19552;
  assign n19555 = ~n19553 & n19554;
  assign n66844 = n19388 | n19390;
  assign n66845 = (n19388 & n50727) | (n19388 & n66844) | (n50727 & n66844);
  assign n50805 = n19555 & n66845;
  assign n66846 = n19231 | n19388;
  assign n66847 = (n19388 & n19390) | (n19388 & n66846) | (n19390 & n66846);
  assign n50806 = n19555 & n66847;
  assign n50807 = (n66773 & n50805) | (n66773 & n50806) | (n50805 & n50806);
  assign n50808 = n19555 | n66845;
  assign n50809 = n19555 | n66847;
  assign n50810 = (n66773 & n50808) | (n66773 & n50809) | (n50808 & n50809);
  assign n19558 = ~n50807 & n50810;
  assign n19559 = x131 & x179;
  assign n19560 = n19558 & n19559;
  assign n19561 = n19558 | n19559;
  assign n19562 = ~n19560 & n19561;
  assign n66832 = n19395 | n19397;
  assign n66833 = (n19395 & n50725) | (n19395 & n66832) | (n50725 & n66832);
  assign n66848 = n19562 & n66833;
  assign n66834 = n19238 | n19395;
  assign n66835 = (n19395 & n19397) | (n19395 & n66834) | (n19397 & n66834);
  assign n66849 = n19562 & n66835;
  assign n66850 = (n66767 & n66848) | (n66767 & n66849) | (n66848 & n66849);
  assign n66851 = n19562 | n66833;
  assign n66852 = n19562 | n66835;
  assign n66853 = (n66767 & n66851) | (n66767 & n66852) | (n66851 & n66852);
  assign n19565 = ~n66850 & n66853;
  assign n19566 = x130 & x180;
  assign n19567 = n19565 & n19566;
  assign n19568 = n19565 | n19566;
  assign n19569 = ~n19567 & n19568;
  assign n50788 = n19402 | n19404;
  assign n50811 = n19569 & n50788;
  assign n50812 = n19402 & n19569;
  assign n50813 = (n66810 & n50811) | (n66810 & n50812) | (n50811 & n50812);
  assign n50814 = n19569 | n50788;
  assign n50815 = n19402 | n19569;
  assign n50816 = (n66810 & n50814) | (n66810 & n50815) | (n50814 & n50815);
  assign n19572 = ~n50813 & n50816;
  assign n19573 = x129 & x181;
  assign n19574 = n19572 & n19573;
  assign n19575 = n19572 | n19573;
  assign n19576 = ~n19574 & n19575;
  assign n50817 = n19409 & n19576;
  assign n66854 = (n19576 & n50746) | (n19576 & n50817) | (n50746 & n50817);
  assign n66855 = (n19576 & n50745) | (n19576 & n50817) | (n50745 & n50817);
  assign n66856 = (n66760 & n66854) | (n66760 & n66855) | (n66854 & n66855);
  assign n50819 = n19409 | n19576;
  assign n66857 = n50746 | n50819;
  assign n66858 = n50745 | n50819;
  assign n66859 = (n66760 & n66857) | (n66760 & n66858) | (n66857 & n66858);
  assign n19579 = ~n66856 & n66859;
  assign n19580 = x128 & x182;
  assign n19581 = n19579 & n19580;
  assign n19582 = n19579 | n19580;
  assign n19583 = ~n19581 & n19582;
  assign n19584 = n66831 & n19583;
  assign n19585 = n66831 | n19583;
  assign n19586 = ~n19584 & n19585;
  assign n19587 = x127 & x183;
  assign n19588 = n19586 & n19587;
  assign n19589 = n19586 | n19587;
  assign n19590 = ~n19588 & n19589;
  assign n50783 = n19423 | n19425;
  assign n50821 = n19590 & n50783;
  assign n50822 = n19423 & n19590;
  assign n50823 = (n66805 & n50821) | (n66805 & n50822) | (n50821 & n50822);
  assign n50824 = n19590 | n50783;
  assign n50825 = n19423 | n19590;
  assign n50826 = (n66805 & n50824) | (n66805 & n50825) | (n50824 & n50825);
  assign n19593 = ~n50823 & n50826;
  assign n19594 = x126 & x184;
  assign n19595 = n19593 & n19594;
  assign n19596 = n19593 | n19594;
  assign n19597 = ~n19595 & n19596;
  assign n50827 = n19430 & n19597;
  assign n66860 = (n19597 & n50755) | (n19597 & n50827) | (n50755 & n50827);
  assign n66861 = (n19432 & n19597) | (n19432 & n50827) | (n19597 & n50827);
  assign n66862 = (n50694 & n66860) | (n50694 & n66861) | (n66860 & n66861);
  assign n50829 = n19430 | n19597;
  assign n66863 = n50755 | n50829;
  assign n66864 = n19432 | n50829;
  assign n66865 = (n50694 & n66863) | (n50694 & n66864) | (n66863 & n66864);
  assign n19600 = ~n66862 & n66865;
  assign n19601 = x125 & x185;
  assign n19602 = n19600 & n19601;
  assign n19603 = n19600 | n19601;
  assign n19604 = ~n19602 & n19603;
  assign n50831 = n19437 & n19604;
  assign n50832 = (n19604 & n50760) | (n19604 & n50831) | (n50760 & n50831);
  assign n50833 = n19437 | n19604;
  assign n50834 = n50760 | n50833;
  assign n19607 = ~n50832 & n50834;
  assign n19608 = x124 & x186;
  assign n19609 = n19607 & n19608;
  assign n19610 = n19607 | n19608;
  assign n19611 = ~n19609 & n19610;
  assign n19612 = n50782 & n19611;
  assign n19613 = n50782 | n19611;
  assign n19614 = ~n19612 & n19613;
  assign n19615 = x123 & x187;
  assign n19616 = n19614 & n19615;
  assign n19617 = n19614 | n19615;
  assign n19618 = ~n19616 & n19617;
  assign n19619 = n50780 & n19618;
  assign n19620 = n50780 | n19618;
  assign n19621 = ~n19619 & n19620;
  assign n19622 = x122 & x188;
  assign n19623 = n19621 & n19622;
  assign n19624 = n19621 | n19622;
  assign n19625 = ~n19623 & n19624;
  assign n19626 = n50778 & n19625;
  assign n19627 = n50778 | n19625;
  assign n19628 = ~n19626 & n19627;
  assign n19629 = x121 & x189;
  assign n19630 = n19628 & n19629;
  assign n19631 = n19628 | n19629;
  assign n19632 = ~n19630 & n19631;
  assign n19633 = n50776 & n19632;
  assign n19634 = n50776 | n19632;
  assign n19635 = ~n19633 & n19634;
  assign n19636 = x120 & x190;
  assign n19637 = n19635 & n19636;
  assign n19638 = n19635 | n19636;
  assign n19639 = ~n19637 & n19638;
  assign n19640 = n50774 & n19639;
  assign n19641 = n50774 | n19639;
  assign n19642 = ~n19640 & n19641;
  assign n19643 = x119 & x191;
  assign n19644 = n19642 & n19643;
  assign n19645 = n19642 | n19643;
  assign n19646 = ~n19644 & n19645;
  assign n19647 = n50772 & n19646;
  assign n19648 = n50772 | n19646;
  assign n19649 = ~n19647 & n19648;
  assign n19650 = x118 & x192;
  assign n19651 = n19649 & n19650;
  assign n19652 = n19649 | n19650;
  assign n19653 = ~n19651 & n19652;
  assign n19654 = n66826 & n19653;
  assign n19655 = n66826 | n19653;
  assign n19656 = ~n19654 & n19655;
  assign n19657 = x117 & x193;
  assign n19658 = n19656 & n19657;
  assign n19659 = n19656 | n19657;
  assign n19660 = ~n19658 & n19659;
  assign n19661 = n50770 & n19660;
  assign n19662 = n50770 | n19660;
  assign n19663 = ~n19661 & n19662;
  assign n19664 = x116 & x194;
  assign n19665 = n19663 & n19664;
  assign n19666 = n19663 | n19664;
  assign n19667 = ~n19665 & n19666;
  assign n19668 = n50768 & n19667;
  assign n19669 = n50768 | n19667;
  assign n19670 = ~n19668 & n19669;
  assign n19671 = x115 & x195;
  assign n19672 = n19670 & n19671;
  assign n19673 = n19670 | n19671;
  assign n19674 = ~n19672 & n19673;
  assign n19675 = n50766 & n19674;
  assign n19676 = n50766 | n19674;
  assign n19677 = ~n19675 & n19676;
  assign n19678 = x114 & x196;
  assign n19679 = n19677 & n19678;
  assign n19680 = n19677 | n19678;
  assign n19681 = ~n19679 & n19680;
  assign n19682 = n50764 & n19681;
  assign n19683 = n50764 | n19681;
  assign n19684 = ~n19682 & n19683;
  assign n19685 = x113 & x197;
  assign n19686 = n19684 & n19685;
  assign n19687 = n19684 | n19685;
  assign n19688 = ~n19686 & n19687;
  assign n19689 = n19521 & n19688;
  assign n19690 = n19521 | n19688;
  assign n19691 = ~n19689 & n19690;
  assign n19692 = x112 & x198;
  assign n19693 = n19691 & n19692;
  assign n19694 = n19691 | n19692;
  assign n19695 = ~n19693 & n19694;
  assign n50835 = n19521 | n19686;
  assign n50836 = (n19686 & n19688) | (n19686 & n50835) | (n19688 & n50835);
  assign n50837 = n19679 | n50764;
  assign n50838 = (n19679 & n19681) | (n19679 & n50837) | (n19681 & n50837);
  assign n50839 = n19672 | n50766;
  assign n50840 = (n19672 & n19674) | (n19672 & n50839) | (n19674 & n50839);
  assign n50841 = n19665 | n50768;
  assign n50842 = (n19665 & n19667) | (n19665 & n50841) | (n19667 & n50841);
  assign n50843 = n19658 | n50770;
  assign n50844 = (n19658 & n19660) | (n19658 & n50843) | (n19660 & n50843);
  assign n50845 = n19651 | n19653;
  assign n50846 = (n66826 & n19651) | (n66826 & n50845) | (n19651 & n50845);
  assign n50847 = n19644 | n19646;
  assign n50848 = (n19644 & n50772) | (n19644 & n50847) | (n50772 & n50847);
  assign n50849 = n19637 | n19639;
  assign n50850 = (n19637 & n50774) | (n19637 & n50849) | (n50774 & n50849);
  assign n50851 = n19630 | n19632;
  assign n50852 = (n19630 & n50776) | (n19630 & n50851) | (n50776 & n50851);
  assign n50853 = n19623 | n19625;
  assign n50854 = (n19623 & n50778) | (n19623 & n50853) | (n50778 & n50853);
  assign n50855 = n19616 | n19618;
  assign n50856 = (n19616 & n50780) | (n19616 & n50855) | (n50780 & n50855);
  assign n50857 = n19609 | n19611;
  assign n50858 = (n19609 & n50782) | (n19609 & n50857) | (n50782 & n50857);
  assign n50860 = n19595 | n19597;
  assign n66866 = n19430 | n19595;
  assign n66867 = (n19595 & n19597) | (n19595 & n66866) | (n19597 & n66866);
  assign n66868 = (n50755 & n50860) | (n50755 & n66867) | (n50860 & n66867);
  assign n66869 = (n19432 & n50860) | (n19432 & n66867) | (n50860 & n66867);
  assign n66870 = (n50694 & n66868) | (n50694 & n66869) | (n66868 & n66869);
  assign n50865 = n19574 | n19576;
  assign n66871 = n19409 | n19574;
  assign n66872 = (n19574 & n19576) | (n19574 & n66871) | (n19576 & n66871);
  assign n66873 = (n50746 & n50865) | (n50746 & n66872) | (n50865 & n66872);
  assign n66874 = (n50745 & n50865) | (n50745 & n66872) | (n50865 & n66872);
  assign n66875 = (n66760 & n66873) | (n66760 & n66874) | (n66873 & n66874);
  assign n19717 = x135 & x176;
  assign n19718 = x134 & x177;
  assign n19719 = n19717 & n19718;
  assign n19720 = n19717 | n19718;
  assign n19721 = ~n19719 & n19720;
  assign n66883 = n19546 | n19548;
  assign n66884 = (n19546 & n66837) | (n19546 & n66883) | (n66837 & n66883);
  assign n50878 = n19721 & n66884;
  assign n66885 = (n19546 & n50797) | (n19546 & n66883) | (n50797 & n66883);
  assign n50879 = n19721 & n66885;
  assign n66886 = (n50878 & n50879) | (n50878 & n66780) | (n50879 & n66780);
  assign n66887 = (n50878 & n50879) | (n50878 & n66778) | (n50879 & n66778);
  assign n66888 = (n66659 & n66886) | (n66659 & n66887) | (n66886 & n66887);
  assign n50881 = n19721 | n66884;
  assign n50882 = n19721 | n66885;
  assign n66889 = (n50881 & n50882) | (n50881 & n66780) | (n50882 & n66780);
  assign n66890 = (n50881 & n50882) | (n50881 & n66778) | (n50882 & n66778);
  assign n66891 = (n66659 & n66889) | (n66659 & n66890) | (n66889 & n66890);
  assign n19724 = ~n66888 & n66891;
  assign n19725 = x133 & x178;
  assign n19726 = n19724 & n19725;
  assign n19727 = n19724 | n19725;
  assign n19728 = ~n19726 & n19727;
  assign n66880 = n19553 | n19555;
  assign n66882 = (n19553 & n66845) | (n19553 & n66880) | (n66845 & n66880);
  assign n66892 = n19728 & n66882;
  assign n66881 = (n19553 & n66847) | (n19553 & n66880) | (n66847 & n66880);
  assign n66893 = n19728 & n66881;
  assign n66894 = (n66773 & n66892) | (n66773 & n66893) | (n66892 & n66893);
  assign n66895 = n19728 | n66882;
  assign n66896 = n19728 | n66881;
  assign n66897 = (n66773 & n66895) | (n66773 & n66896) | (n66895 & n66896);
  assign n19731 = ~n66894 & n66897;
  assign n19732 = x132 & x179;
  assign n19733 = n19731 & n19732;
  assign n19734 = n19731 | n19732;
  assign n19735 = ~n19733 & n19734;
  assign n50870 = n19560 | n19562;
  assign n50884 = n19735 & n50870;
  assign n50885 = n19560 & n19735;
  assign n66898 = (n50884 & n50885) | (n50884 & n66833) | (n50885 & n66833);
  assign n66899 = (n50884 & n50885) | (n50884 & n66835) | (n50885 & n66835);
  assign n66900 = (n66767 & n66898) | (n66767 & n66899) | (n66898 & n66899);
  assign n50887 = n19735 | n50870;
  assign n50888 = n19560 | n19735;
  assign n66901 = (n50887 & n50888) | (n50887 & n66833) | (n50888 & n66833);
  assign n66902 = (n50887 & n50888) | (n50887 & n66835) | (n50888 & n66835);
  assign n66903 = (n66767 & n66901) | (n66767 & n66902) | (n66901 & n66902);
  assign n19738 = ~n66900 & n66903;
  assign n19739 = x131 & x180;
  assign n19740 = n19738 & n19739;
  assign n19741 = n19738 | n19739;
  assign n19742 = ~n19740 & n19741;
  assign n66878 = n19567 | n19569;
  assign n66879 = (n19567 & n50788) | (n19567 & n66878) | (n50788 & n66878);
  assign n66904 = n19742 & n66879;
  assign n66876 = n19402 | n19567;
  assign n66877 = (n19567 & n19569) | (n19567 & n66876) | (n19569 & n66876);
  assign n66905 = n19742 & n66877;
  assign n66906 = (n66810 & n66904) | (n66810 & n66905) | (n66904 & n66905);
  assign n66907 = n19742 | n66879;
  assign n66908 = n19742 | n66877;
  assign n66909 = (n66810 & n66907) | (n66810 & n66908) | (n66907 & n66908);
  assign n19745 = ~n66906 & n66909;
  assign n19746 = x130 & x181;
  assign n19747 = n19745 & n19746;
  assign n19748 = n19745 | n19746;
  assign n19749 = ~n19747 & n19748;
  assign n19750 = n66875 & n19749;
  assign n19751 = n66875 | n19749;
  assign n19752 = ~n19750 & n19751;
  assign n19753 = x129 & x182;
  assign n19754 = n19752 & n19753;
  assign n19755 = n19752 | n19753;
  assign n19756 = ~n19754 & n19755;
  assign n50862 = n19581 | n19583;
  assign n50890 = n19756 & n50862;
  assign n50891 = n19581 & n19756;
  assign n50892 = (n66831 & n50890) | (n66831 & n50891) | (n50890 & n50891);
  assign n50893 = n19756 | n50862;
  assign n50894 = n19581 | n19756;
  assign n50895 = (n66831 & n50893) | (n66831 & n50894) | (n50893 & n50894);
  assign n19759 = ~n50892 & n50895;
  assign n19760 = x128 & x183;
  assign n19761 = n19759 & n19760;
  assign n19762 = n19759 | n19760;
  assign n19763 = ~n19761 & n19762;
  assign n50896 = n19588 & n19763;
  assign n66910 = (n19763 & n50822) | (n19763 & n50896) | (n50822 & n50896);
  assign n66911 = (n19763 & n50821) | (n19763 & n50896) | (n50821 & n50896);
  assign n66912 = (n66805 & n66910) | (n66805 & n66911) | (n66910 & n66911);
  assign n50898 = n19588 | n19763;
  assign n66913 = n50822 | n50898;
  assign n66914 = n50821 | n50898;
  assign n66915 = (n66805 & n66913) | (n66805 & n66914) | (n66913 & n66914);
  assign n19766 = ~n66912 & n66915;
  assign n19767 = x127 & x184;
  assign n19768 = n19766 & n19767;
  assign n19769 = n19766 | n19767;
  assign n19770 = ~n19768 & n19769;
  assign n19771 = n66870 & n19770;
  assign n19772 = n66870 | n19770;
  assign n19773 = ~n19771 & n19772;
  assign n19774 = x126 & x185;
  assign n19775 = n19773 & n19774;
  assign n19776 = n19773 | n19774;
  assign n19777 = ~n19775 & n19776;
  assign n50900 = n19602 & n19777;
  assign n50901 = (n19777 & n50832) | (n19777 & n50900) | (n50832 & n50900);
  assign n50902 = n19602 | n19777;
  assign n50903 = n50832 | n50902;
  assign n19780 = ~n50901 & n50903;
  assign n19781 = x125 & x186;
  assign n19782 = n19780 & n19781;
  assign n19783 = n19780 | n19781;
  assign n19784 = ~n19782 & n19783;
  assign n19785 = n50858 & n19784;
  assign n19786 = n50858 | n19784;
  assign n19787 = ~n19785 & n19786;
  assign n19788 = x124 & x187;
  assign n19789 = n19787 & n19788;
  assign n19790 = n19787 | n19788;
  assign n19791 = ~n19789 & n19790;
  assign n19792 = n50856 & n19791;
  assign n19793 = n50856 | n19791;
  assign n19794 = ~n19792 & n19793;
  assign n19795 = x123 & x188;
  assign n19796 = n19794 & n19795;
  assign n19797 = n19794 | n19795;
  assign n19798 = ~n19796 & n19797;
  assign n19799 = n50854 & n19798;
  assign n19800 = n50854 | n19798;
  assign n19801 = ~n19799 & n19800;
  assign n19802 = x122 & x189;
  assign n19803 = n19801 & n19802;
  assign n19804 = n19801 | n19802;
  assign n19805 = ~n19803 & n19804;
  assign n19806 = n50852 & n19805;
  assign n19807 = n50852 | n19805;
  assign n19808 = ~n19806 & n19807;
  assign n19809 = x121 & x190;
  assign n19810 = n19808 & n19809;
  assign n19811 = n19808 | n19809;
  assign n19812 = ~n19810 & n19811;
  assign n19813 = n50850 & n19812;
  assign n19814 = n50850 | n19812;
  assign n19815 = ~n19813 & n19814;
  assign n19816 = x120 & x191;
  assign n19817 = n19815 & n19816;
  assign n19818 = n19815 | n19816;
  assign n19819 = ~n19817 & n19818;
  assign n19820 = n50848 & n19819;
  assign n19821 = n50848 | n19819;
  assign n19822 = ~n19820 & n19821;
  assign n19823 = x119 & x192;
  assign n19824 = n19822 & n19823;
  assign n19825 = n19822 | n19823;
  assign n19826 = ~n19824 & n19825;
  assign n19827 = n50846 & n19826;
  assign n19828 = n50846 | n19826;
  assign n19829 = ~n19827 & n19828;
  assign n19830 = x118 & x193;
  assign n19831 = n19829 & n19830;
  assign n19832 = n19829 | n19830;
  assign n19833 = ~n19831 & n19832;
  assign n19834 = n50844 & n19833;
  assign n19835 = n50844 | n19833;
  assign n19836 = ~n19834 & n19835;
  assign n19837 = x117 & x194;
  assign n19838 = n19836 & n19837;
  assign n19839 = n19836 | n19837;
  assign n19840 = ~n19838 & n19839;
  assign n19841 = n50842 & n19840;
  assign n19842 = n50842 | n19840;
  assign n19843 = ~n19841 & n19842;
  assign n19844 = x116 & x195;
  assign n19845 = n19843 & n19844;
  assign n19846 = n19843 | n19844;
  assign n19847 = ~n19845 & n19846;
  assign n19848 = n50840 & n19847;
  assign n19849 = n50840 | n19847;
  assign n19850 = ~n19848 & n19849;
  assign n19851 = x115 & x196;
  assign n19852 = n19850 & n19851;
  assign n19853 = n19850 | n19851;
  assign n19854 = ~n19852 & n19853;
  assign n19855 = n50838 & n19854;
  assign n19856 = n50838 | n19854;
  assign n19857 = ~n19855 & n19856;
  assign n19858 = x114 & x197;
  assign n19859 = n19857 & n19858;
  assign n19860 = n19857 | n19858;
  assign n19861 = ~n19859 & n19860;
  assign n19862 = n50836 & n19861;
  assign n19863 = n50836 | n19861;
  assign n19864 = ~n19862 & n19863;
  assign n19865 = x113 & x198;
  assign n19866 = n19864 & n19865;
  assign n19867 = n19864 | n19865;
  assign n19868 = ~n19866 & n19867;
  assign n19869 = n19693 & n19868;
  assign n19870 = n19693 | n19868;
  assign n19871 = ~n19869 & n19870;
  assign n19872 = x112 & x199;
  assign n19873 = n19871 & n19872;
  assign n19874 = n19871 | n19872;
  assign n19875 = ~n19873 & n19874;
  assign n66916 = n19693 | n19865;
  assign n66917 = (n19693 & n19864) | (n19693 & n66916) | (n19864 & n66916);
  assign n50905 = (n19866 & n19868) | (n19866 & n66917) | (n19868 & n66917);
  assign n66918 = n19859 | n50836;
  assign n66919 = (n19859 & n19861) | (n19859 & n66918) | (n19861 & n66918);
  assign n19878 = n19852 | n19855;
  assign n19879 = n19845 | n19848;
  assign n19880 = n19838 | n19841;
  assign n19881 = n19831 | n19834;
  assign n50906 = n19824 | n19826;
  assign n50907 = (n19824 & n50846) | (n19824 & n50906) | (n50846 & n50906);
  assign n50908 = n19817 | n19819;
  assign n50909 = (n19817 & n50848) | (n19817 & n50908) | (n50848 & n50908);
  assign n50910 = n19810 | n19812;
  assign n50911 = (n19810 & n50850) | (n19810 & n50910) | (n50850 & n50910);
  assign n50912 = n19803 | n19805;
  assign n50913 = (n19803 & n50852) | (n19803 & n50912) | (n50852 & n50912);
  assign n50914 = n19796 | n19798;
  assign n50915 = (n19796 & n50854) | (n19796 & n50914) | (n50854 & n50914);
  assign n50916 = n19789 | n19791;
  assign n50917 = (n19789 & n50856) | (n19789 & n50916) | (n50856 & n50916);
  assign n50918 = n19782 | n19784;
  assign n50919 = (n19782 & n50858) | (n19782 & n50918) | (n50858 & n50918);
  assign n50923 = n19761 | n19763;
  assign n66920 = n19588 | n19761;
  assign n66921 = (n19761 & n19763) | (n19761 & n66920) | (n19763 & n66920);
  assign n66922 = (n50822 & n50923) | (n50822 & n66921) | (n50923 & n66921);
  assign n66923 = (n50821 & n50923) | (n50821 & n66921) | (n50923 & n66921);
  assign n66924 = (n66805 & n66922) | (n66805 & n66923) | (n66922 & n66923);
  assign n50792 = (n66767 & n66833) | (n66767 & n66835) | (n66833 & n66835);
  assign n19898 = x136 & x176;
  assign n19899 = x135 & x177;
  assign n19900 = n19898 & n19899;
  assign n19901 = n19898 | n19899;
  assign n19902 = ~n19900 & n19901;
  assign n66925 = n19719 | n19721;
  assign n66927 = n19902 & n66925;
  assign n66928 = n19719 & n19902;
  assign n66929 = (n66884 & n66927) | (n66884 & n66928) | (n66927 & n66928);
  assign n66931 = (n66885 & n66927) | (n66885 & n66928) | (n66927 & n66928);
  assign n66932 = (n66780 & n66929) | (n66780 & n66931) | (n66929 & n66931);
  assign n66933 = (n66778 & n66929) | (n66778 & n66931) | (n66929 & n66931);
  assign n66934 = (n66659 & n66932) | (n66659 & n66933) | (n66932 & n66933);
  assign n66935 = n19902 | n66925;
  assign n66936 = n19719 | n19902;
  assign n66937 = (n66884 & n66935) | (n66884 & n66936) | (n66935 & n66936);
  assign n66938 = (n66885 & n66935) | (n66885 & n66936) | (n66935 & n66936);
  assign n66939 = (n66780 & n66937) | (n66780 & n66938) | (n66937 & n66938);
  assign n66940 = (n66778 & n66937) | (n66778 & n66938) | (n66937 & n66938);
  assign n66941 = (n66659 & n66939) | (n66659 & n66940) | (n66939 & n66940);
  assign n19905 = ~n66934 & n66941;
  assign n19906 = x134 & x178;
  assign n19907 = n19905 & n19906;
  assign n19908 = n19905 | n19906;
  assign n19909 = ~n19907 & n19908;
  assign n50932 = n19726 | n19728;
  assign n50943 = n19909 & n50932;
  assign n50944 = n19726 & n19909;
  assign n66942 = (n50943 & n50944) | (n50943 & n66882) | (n50944 & n66882);
  assign n66943 = (n50943 & n50944) | (n50943 & n66881) | (n50944 & n66881);
  assign n66944 = (n66773 & n66942) | (n66773 & n66943) | (n66942 & n66943);
  assign n50946 = n19909 | n50932;
  assign n50947 = n19726 | n19909;
  assign n66945 = (n50946 & n50947) | (n50946 & n66882) | (n50947 & n66882);
  assign n66946 = (n50946 & n50947) | (n50946 & n66881) | (n50947 & n66881);
  assign n66947 = (n66773 & n66945) | (n66773 & n66946) | (n66945 & n66946);
  assign n19912 = ~n66944 & n66947;
  assign n19913 = x133 & x179;
  assign n19914 = n19912 & n19913;
  assign n19915 = n19912 | n19913;
  assign n19916 = ~n19914 & n19915;
  assign n66948 = n19733 | n19735;
  assign n66949 = (n19733 & n50870) | (n19733 & n66948) | (n50870 & n66948);
  assign n50949 = n19916 & n66949;
  assign n66950 = n19560 | n19733;
  assign n66951 = (n19733 & n19735) | (n19733 & n66950) | (n19735 & n66950);
  assign n50950 = n19916 & n66951;
  assign n50951 = (n50792 & n50949) | (n50792 & n50950) | (n50949 & n50950);
  assign n50952 = n19916 | n66949;
  assign n50953 = n19916 | n66951;
  assign n50954 = (n50792 & n50952) | (n50792 & n50953) | (n50952 & n50953);
  assign n19919 = ~n50951 & n50954;
  assign n19920 = x132 & x180;
  assign n19921 = n19919 & n19920;
  assign n19922 = n19919 | n19920;
  assign n19923 = ~n19921 & n19922;
  assign n50927 = n19740 | n19742;
  assign n50955 = n19923 & n50927;
  assign n50956 = n19740 & n19923;
  assign n66952 = (n50955 & n50956) | (n50955 & n66879) | (n50956 & n66879);
  assign n66953 = (n50955 & n50956) | (n50955 & n66877) | (n50956 & n66877);
  assign n66954 = (n66810 & n66952) | (n66810 & n66953) | (n66952 & n66953);
  assign n50958 = n19923 | n50927;
  assign n50959 = n19740 | n19923;
  assign n66955 = (n50958 & n50959) | (n50958 & n66879) | (n50959 & n66879);
  assign n66956 = (n50958 & n50959) | (n50958 & n66877) | (n50959 & n66877);
  assign n66957 = (n66810 & n66955) | (n66810 & n66956) | (n66955 & n66956);
  assign n19926 = ~n66954 & n66957;
  assign n19927 = x131 & x181;
  assign n19928 = n19926 & n19927;
  assign n19929 = n19926 | n19927;
  assign n19930 = ~n19928 & n19929;
  assign n50925 = n19747 | n19749;
  assign n50961 = n19930 & n50925;
  assign n50962 = n19747 & n19930;
  assign n50963 = (n66875 & n50961) | (n66875 & n50962) | (n50961 & n50962);
  assign n50964 = n19930 | n50925;
  assign n50965 = n19747 | n19930;
  assign n50966 = (n66875 & n50964) | (n66875 & n50965) | (n50964 & n50965);
  assign n19933 = ~n50963 & n50966;
  assign n19934 = x130 & x182;
  assign n19935 = n19933 & n19934;
  assign n19936 = n19933 | n19934;
  assign n19937 = ~n19935 & n19936;
  assign n50967 = n19754 & n19937;
  assign n66958 = (n19937 & n50891) | (n19937 & n50967) | (n50891 & n50967);
  assign n66959 = (n19937 & n50890) | (n19937 & n50967) | (n50890 & n50967);
  assign n66960 = (n66831 & n66958) | (n66831 & n66959) | (n66958 & n66959);
  assign n50969 = n19754 | n19937;
  assign n66961 = n50891 | n50969;
  assign n66962 = n50890 | n50969;
  assign n66963 = (n66831 & n66961) | (n66831 & n66962) | (n66961 & n66962);
  assign n19940 = ~n66960 & n66963;
  assign n19941 = x129 & x183;
  assign n19942 = n19940 & n19941;
  assign n19943 = n19940 | n19941;
  assign n19944 = ~n19942 & n19943;
  assign n19945 = n66924 & n19944;
  assign n19946 = n66924 | n19944;
  assign n19947 = ~n19945 & n19946;
  assign n19948 = x128 & x184;
  assign n19949 = n19947 & n19948;
  assign n19950 = n19947 | n19948;
  assign n19951 = ~n19949 & n19950;
  assign n50920 = n19768 | n19770;
  assign n50971 = n19951 & n50920;
  assign n50972 = n19768 & n19951;
  assign n50973 = (n66870 & n50971) | (n66870 & n50972) | (n50971 & n50972);
  assign n50974 = n19951 | n50920;
  assign n50975 = n19768 | n19951;
  assign n50976 = (n66870 & n50974) | (n66870 & n50975) | (n50974 & n50975);
  assign n19954 = ~n50973 & n50976;
  assign n19955 = x127 & x185;
  assign n19956 = n19954 & n19955;
  assign n19957 = n19954 | n19955;
  assign n19958 = ~n19956 & n19957;
  assign n50977 = n19775 & n19958;
  assign n66964 = (n19958 & n50900) | (n19958 & n50977) | (n50900 & n50977);
  assign n66965 = (n19777 & n19958) | (n19777 & n50977) | (n19958 & n50977);
  assign n66966 = (n50832 & n66964) | (n50832 & n66965) | (n66964 & n66965);
  assign n50979 = n19775 | n19958;
  assign n66967 = n50900 | n50979;
  assign n66968 = n19777 | n50979;
  assign n66969 = (n50832 & n66967) | (n50832 & n66968) | (n66967 & n66968);
  assign n19961 = ~n66966 & n66969;
  assign n19962 = x126 & x186;
  assign n19963 = n19961 & n19962;
  assign n19964 = n19961 | n19962;
  assign n19965 = ~n19963 & n19964;
  assign n19966 = n50919 & n19965;
  assign n19967 = n50919 | n19965;
  assign n19968 = ~n19966 & n19967;
  assign n19969 = x125 & x187;
  assign n19970 = n19968 & n19969;
  assign n19971 = n19968 | n19969;
  assign n19972 = ~n19970 & n19971;
  assign n19973 = n50917 & n19972;
  assign n19974 = n50917 | n19972;
  assign n19975 = ~n19973 & n19974;
  assign n19976 = x124 & x188;
  assign n19977 = n19975 & n19976;
  assign n19978 = n19975 | n19976;
  assign n19979 = ~n19977 & n19978;
  assign n19980 = n50915 & n19979;
  assign n19981 = n50915 | n19979;
  assign n19982 = ~n19980 & n19981;
  assign n19983 = x123 & x189;
  assign n19984 = n19982 & n19983;
  assign n19985 = n19982 | n19983;
  assign n19986 = ~n19984 & n19985;
  assign n19987 = n50913 & n19986;
  assign n19988 = n50913 | n19986;
  assign n19989 = ~n19987 & n19988;
  assign n19990 = x122 & x190;
  assign n19991 = n19989 & n19990;
  assign n19992 = n19989 | n19990;
  assign n19993 = ~n19991 & n19992;
  assign n19994 = n50911 & n19993;
  assign n19995 = n50911 | n19993;
  assign n19996 = ~n19994 & n19995;
  assign n19997 = x121 & x191;
  assign n19998 = n19996 & n19997;
  assign n19999 = n19996 | n19997;
  assign n20000 = ~n19998 & n19999;
  assign n20001 = n50909 & n20000;
  assign n20002 = n50909 | n20000;
  assign n20003 = ~n20001 & n20002;
  assign n20004 = x120 & x192;
  assign n20005 = n20003 & n20004;
  assign n20006 = n20003 | n20004;
  assign n20007 = ~n20005 & n20006;
  assign n20008 = n50907 & n20007;
  assign n20009 = n50907 | n20007;
  assign n20010 = ~n20008 & n20009;
  assign n20011 = x119 & x193;
  assign n20012 = n20010 & n20011;
  assign n20013 = n20010 | n20011;
  assign n20014 = ~n20012 & n20013;
  assign n20015 = n19881 & n20014;
  assign n20016 = n19881 | n20014;
  assign n20017 = ~n20015 & n20016;
  assign n20018 = x118 & x194;
  assign n20019 = n20017 & n20018;
  assign n20020 = n20017 | n20018;
  assign n20021 = ~n20019 & n20020;
  assign n20022 = n19880 & n20021;
  assign n20023 = n19880 | n20021;
  assign n20024 = ~n20022 & n20023;
  assign n20025 = x117 & x195;
  assign n20026 = n20024 & n20025;
  assign n20027 = n20024 | n20025;
  assign n20028 = ~n20026 & n20027;
  assign n20029 = n19879 & n20028;
  assign n20030 = n19879 | n20028;
  assign n20031 = ~n20029 & n20030;
  assign n20032 = x116 & x196;
  assign n20033 = n20031 & n20032;
  assign n20034 = n20031 | n20032;
  assign n20035 = ~n20033 & n20034;
  assign n20036 = n19878 & n20035;
  assign n20037 = n19878 | n20035;
  assign n20038 = ~n20036 & n20037;
  assign n20039 = x115 & x197;
  assign n20040 = n20038 & n20039;
  assign n20041 = n20038 | n20039;
  assign n20042 = ~n20040 & n20041;
  assign n20043 = n66919 & n20042;
  assign n20044 = n66919 | n20042;
  assign n20045 = ~n20043 & n20044;
  assign n20046 = x114 & x198;
  assign n20047 = n20045 & n20046;
  assign n20048 = n20045 | n20046;
  assign n20049 = ~n20047 & n20048;
  assign n20050 = n50905 & n20049;
  assign n20051 = n50905 | n20049;
  assign n20052 = ~n20050 & n20051;
  assign n20053 = x113 & x199;
  assign n20054 = n20052 & n20053;
  assign n20055 = n20052 | n20053;
  assign n20056 = ~n20054 & n20055;
  assign n20057 = n19873 & n20056;
  assign n20058 = n19873 | n20056;
  assign n20059 = ~n20057 & n20058;
  assign n20060 = x112 & x200;
  assign n20061 = n20059 & n20060;
  assign n20062 = n20059 | n20060;
  assign n20063 = ~n20061 & n20062;
  assign n66970 = n19873 | n20053;
  assign n66971 = (n19873 & n20052) | (n19873 & n66970) | (n20052 & n66970);
  assign n50982 = (n20054 & n20056) | (n20054 & n66971) | (n20056 & n66971);
  assign n50983 = n20047 | n50905;
  assign n50984 = (n20047 & n20049) | (n20047 & n50983) | (n20049 & n50983);
  assign n66972 = n20040 | n66919;
  assign n66973 = (n20040 & n20042) | (n20040 & n66972) | (n20042 & n66972);
  assign n20067 = n20033 | n20036;
  assign n20068 = n20026 | n20029;
  assign n20069 = n20019 | n20022;
  assign n50985 = n20012 | n20014;
  assign n50986 = (n19881 & n20012) | (n19881 & n50985) | (n20012 & n50985);
  assign n50987 = n20005 | n20007;
  assign n50988 = (n20005 & n50907) | (n20005 & n50987) | (n50907 & n50987);
  assign n50989 = n19998 | n20000;
  assign n50990 = (n19998 & n50909) | (n19998 & n50989) | (n50909 & n50989);
  assign n50991 = n19991 | n19993;
  assign n50992 = (n19991 & n50911) | (n19991 & n50991) | (n50911 & n50991);
  assign n50993 = n19984 | n19986;
  assign n50994 = (n19984 & n50913) | (n19984 & n50993) | (n50913 & n50993);
  assign n50995 = n19977 | n19979;
  assign n50996 = (n19977 & n50915) | (n19977 & n50995) | (n50915 & n50995);
  assign n50997 = n19970 | n19972;
  assign n50998 = (n19970 & n50917) | (n19970 & n50997) | (n50917 & n50997);
  assign n51002 = n19956 | n19958;
  assign n66974 = n19775 | n19956;
  assign n66975 = (n19956 & n19958) | (n19956 & n66974) | (n19958 & n66974);
  assign n66976 = (n50900 & n51002) | (n50900 & n66975) | (n51002 & n66975);
  assign n66977 = (n19777 & n51002) | (n19777 & n66975) | (n51002 & n66975);
  assign n66978 = (n50832 & n66976) | (n50832 & n66977) | (n66976 & n66977);
  assign n51007 = n19935 | n19937;
  assign n66979 = n19754 | n19935;
  assign n66980 = (n19935 & n19937) | (n19935 & n66979) | (n19937 & n66979);
  assign n66981 = (n50891 & n51007) | (n50891 & n66980) | (n51007 & n66980);
  assign n66982 = (n50890 & n51007) | (n50890 & n66980) | (n51007 & n66980);
  assign n66983 = (n66831 & n66981) | (n66831 & n66982) | (n66981 & n66982);
  assign n50869 = (n66810 & n66877) | (n66810 & n66879) | (n66877 & n66879);
  assign n51015 = n19900 | n66929;
  assign n51016 = n19900 | n66931;
  assign n66986 = (n51015 & n51016) | (n51015 & n66780) | (n51016 & n66780);
  assign n66987 = (n51015 & n51016) | (n51015 & n66778) | (n51016 & n66778);
  assign n66988 = (n66659 & n66986) | (n66659 & n66987) | (n66986 & n66987);
  assign n20087 = x137 & x176;
  assign n20088 = x136 & x177;
  assign n20089 = n20087 & n20088;
  assign n20090 = n20087 | n20088;
  assign n20091 = ~n20089 & n20090;
  assign n20092 = n66988 & n20091;
  assign n20093 = n66988 | n20091;
  assign n20094 = ~n20092 & n20093;
  assign n20095 = x135 & x178;
  assign n20096 = n20094 & n20095;
  assign n20097 = n20094 | n20095;
  assign n20098 = ~n20096 & n20097;
  assign n66989 = n19907 | n19909;
  assign n66990 = (n19907 & n50932) | (n19907 & n66989) | (n50932 & n66989);
  assign n51018 = n20098 & n66990;
  assign n66991 = n19726 | n19907;
  assign n66992 = (n19907 & n19909) | (n19907 & n66991) | (n19909 & n66991);
  assign n51019 = n20098 & n66992;
  assign n66993 = (n51018 & n51019) | (n51018 & n66882) | (n51019 & n66882);
  assign n66994 = (n51018 & n51019) | (n51018 & n66881) | (n51019 & n66881);
  assign n66995 = (n66773 & n66993) | (n66773 & n66994) | (n66993 & n66994);
  assign n51021 = n20098 | n66990;
  assign n51022 = n20098 | n66992;
  assign n66996 = (n51021 & n51022) | (n51021 & n66882) | (n51022 & n66882);
  assign n66997 = (n51021 & n51022) | (n51021 & n66881) | (n51022 & n66881);
  assign n66998 = (n66773 & n66996) | (n66773 & n66997) | (n66996 & n66997);
  assign n20101 = ~n66995 & n66998;
  assign n20102 = x134 & x179;
  assign n20103 = n20101 & n20102;
  assign n20104 = n20101 | n20102;
  assign n20105 = ~n20103 & n20104;
  assign n51024 = n19914 & n20105;
  assign n66999 = (n20105 & n50949) | (n20105 & n51024) | (n50949 & n51024);
  assign n67000 = (n20105 & n50950) | (n20105 & n51024) | (n50950 & n51024);
  assign n67001 = (n50792 & n66999) | (n50792 & n67000) | (n66999 & n67000);
  assign n51026 = n19914 | n20105;
  assign n67002 = n50949 | n51026;
  assign n67003 = n50950 | n51026;
  assign n67004 = (n50792 & n67002) | (n50792 & n67003) | (n67002 & n67003);
  assign n20108 = ~n67001 & n67004;
  assign n20109 = x133 & x180;
  assign n20110 = n20108 & n20109;
  assign n20111 = n20108 | n20109;
  assign n20112 = ~n20110 & n20111;
  assign n51009 = n19921 | n50955;
  assign n67005 = n20112 & n51009;
  assign n66984 = n19740 | n19921;
  assign n66985 = (n19921 & n19923) | (n19921 & n66984) | (n19923 & n66984);
  assign n67006 = n20112 & n66985;
  assign n67007 = (n50869 & n67005) | (n50869 & n67006) | (n67005 & n67006);
  assign n67008 = n20112 | n51009;
  assign n67009 = n20112 | n66985;
  assign n67010 = (n50869 & n67008) | (n50869 & n67009) | (n67008 & n67009);
  assign n20115 = ~n67007 & n67010;
  assign n20116 = x132 & x181;
  assign n20117 = n20115 & n20116;
  assign n20118 = n20115 | n20116;
  assign n20119 = ~n20117 & n20118;
  assign n51028 = n19928 & n20119;
  assign n67011 = (n20119 & n50961) | (n20119 & n51028) | (n50961 & n51028);
  assign n67012 = (n20119 & n50962) | (n20119 & n51028) | (n50962 & n51028);
  assign n67013 = (n66875 & n67011) | (n66875 & n67012) | (n67011 & n67012);
  assign n51030 = n19928 | n20119;
  assign n67014 = n50961 | n51030;
  assign n67015 = n50962 | n51030;
  assign n67016 = (n66875 & n67014) | (n66875 & n67015) | (n67014 & n67015);
  assign n20122 = ~n67013 & n67016;
  assign n20123 = x131 & x182;
  assign n20124 = n20122 & n20123;
  assign n20125 = n20122 | n20123;
  assign n20126 = ~n20124 & n20125;
  assign n20127 = n66983 & n20126;
  assign n20128 = n66983 | n20126;
  assign n20129 = ~n20127 & n20128;
  assign n20130 = x130 & x183;
  assign n20131 = n20129 & n20130;
  assign n20132 = n20129 | n20130;
  assign n20133 = ~n20131 & n20132;
  assign n51004 = n19942 | n19944;
  assign n51032 = n20133 & n51004;
  assign n51033 = n19942 & n20133;
  assign n51034 = (n66924 & n51032) | (n66924 & n51033) | (n51032 & n51033);
  assign n51035 = n20133 | n51004;
  assign n51036 = n19942 | n20133;
  assign n51037 = (n66924 & n51035) | (n66924 & n51036) | (n51035 & n51036);
  assign n20136 = ~n51034 & n51037;
  assign n20137 = x129 & x184;
  assign n20138 = n20136 & n20137;
  assign n20139 = n20136 | n20137;
  assign n20140 = ~n20138 & n20139;
  assign n51038 = n19949 & n20140;
  assign n67017 = (n20140 & n50972) | (n20140 & n51038) | (n50972 & n51038);
  assign n67018 = (n20140 & n50971) | (n20140 & n51038) | (n50971 & n51038);
  assign n67019 = (n66870 & n67017) | (n66870 & n67018) | (n67017 & n67018);
  assign n51040 = n19949 | n20140;
  assign n67020 = n50972 | n51040;
  assign n67021 = n50971 | n51040;
  assign n67022 = (n66870 & n67020) | (n66870 & n67021) | (n67020 & n67021);
  assign n20143 = ~n67019 & n67022;
  assign n20144 = x128 & x185;
  assign n20145 = n20143 & n20144;
  assign n20146 = n20143 | n20144;
  assign n20147 = ~n20145 & n20146;
  assign n20148 = n66978 & n20147;
  assign n20149 = n66978 | n20147;
  assign n20150 = ~n20148 & n20149;
  assign n20151 = x127 & x186;
  assign n20152 = n20150 & n20151;
  assign n20153 = n20150 | n20151;
  assign n20154 = ~n20152 & n20153;
  assign n50999 = n19963 | n19965;
  assign n67023 = n20154 & n50999;
  assign n67024 = n19963 & n20154;
  assign n67025 = (n50919 & n67023) | (n50919 & n67024) | (n67023 & n67024);
  assign n67026 = n20154 | n50999;
  assign n67027 = n19963 | n20154;
  assign n67028 = (n50919 & n67026) | (n50919 & n67027) | (n67026 & n67027);
  assign n20157 = ~n67025 & n67028;
  assign n20158 = x126 & x187;
  assign n20159 = n20157 & n20158;
  assign n20160 = n20157 | n20158;
  assign n20161 = ~n20159 & n20160;
  assign n20162 = n50998 & n20161;
  assign n20163 = n50998 | n20161;
  assign n20164 = ~n20162 & n20163;
  assign n20165 = x125 & x188;
  assign n20166 = n20164 & n20165;
  assign n20167 = n20164 | n20165;
  assign n20168 = ~n20166 & n20167;
  assign n20169 = n50996 & n20168;
  assign n20170 = n50996 | n20168;
  assign n20171 = ~n20169 & n20170;
  assign n20172 = x124 & x189;
  assign n20173 = n20171 & n20172;
  assign n20174 = n20171 | n20172;
  assign n20175 = ~n20173 & n20174;
  assign n20176 = n50994 & n20175;
  assign n20177 = n50994 | n20175;
  assign n20178 = ~n20176 & n20177;
  assign n20179 = x123 & x190;
  assign n20180 = n20178 & n20179;
  assign n20181 = n20178 | n20179;
  assign n20182 = ~n20180 & n20181;
  assign n20183 = n50992 & n20182;
  assign n20184 = n50992 | n20182;
  assign n20185 = ~n20183 & n20184;
  assign n20186 = x122 & x191;
  assign n20187 = n20185 & n20186;
  assign n20188 = n20185 | n20186;
  assign n20189 = ~n20187 & n20188;
  assign n20190 = n50990 & n20189;
  assign n20191 = n50990 | n20189;
  assign n20192 = ~n20190 & n20191;
  assign n20193 = x121 & x192;
  assign n20194 = n20192 & n20193;
  assign n20195 = n20192 | n20193;
  assign n20196 = ~n20194 & n20195;
  assign n20197 = n50988 & n20196;
  assign n20198 = n50988 | n20196;
  assign n20199 = ~n20197 & n20198;
  assign n20200 = x120 & x193;
  assign n20201 = n20199 & n20200;
  assign n20202 = n20199 | n20200;
  assign n20203 = ~n20201 & n20202;
  assign n20204 = n50986 & n20203;
  assign n20205 = n50986 | n20203;
  assign n20206 = ~n20204 & n20205;
  assign n20207 = x119 & x194;
  assign n20208 = n20206 & n20207;
  assign n20209 = n20206 | n20207;
  assign n20210 = ~n20208 & n20209;
  assign n20211 = n20069 & n20210;
  assign n20212 = n20069 | n20210;
  assign n20213 = ~n20211 & n20212;
  assign n20214 = x118 & x195;
  assign n20215 = n20213 & n20214;
  assign n20216 = n20213 | n20214;
  assign n20217 = ~n20215 & n20216;
  assign n20218 = n20068 & n20217;
  assign n20219 = n20068 | n20217;
  assign n20220 = ~n20218 & n20219;
  assign n20221 = x117 & x196;
  assign n20222 = n20220 & n20221;
  assign n20223 = n20220 | n20221;
  assign n20224 = ~n20222 & n20223;
  assign n20225 = n20067 & n20224;
  assign n20226 = n20067 | n20224;
  assign n20227 = ~n20225 & n20226;
  assign n20228 = x116 & x197;
  assign n20229 = n20227 & n20228;
  assign n20230 = n20227 | n20228;
  assign n20231 = ~n20229 & n20230;
  assign n20232 = n66973 & n20231;
  assign n20233 = n66973 | n20231;
  assign n20234 = ~n20232 & n20233;
  assign n20235 = x115 & x198;
  assign n20236 = n20234 & n20235;
  assign n20237 = n20234 | n20235;
  assign n20238 = ~n20236 & n20237;
  assign n20239 = n50984 & n20238;
  assign n20240 = n50984 | n20238;
  assign n20241 = ~n20239 & n20240;
  assign n20242 = x114 & x199;
  assign n20243 = n20241 & n20242;
  assign n20244 = n20241 | n20242;
  assign n20245 = ~n20243 & n20244;
  assign n20246 = n50982 & n20245;
  assign n20247 = n50982 | n20245;
  assign n20248 = ~n20246 & n20247;
  assign n20249 = x113 & x200;
  assign n20250 = n20248 & n20249;
  assign n20251 = n20248 | n20249;
  assign n20252 = ~n20250 & n20251;
  assign n20253 = n20061 & n20252;
  assign n20254 = n20061 | n20252;
  assign n20255 = ~n20253 & n20254;
  assign n20256 = x112 & x201;
  assign n20257 = n20255 & n20256;
  assign n20258 = n20255 | n20256;
  assign n20259 = ~n20257 & n20258;
  assign n67029 = n20061 | n20249;
  assign n67030 = (n20061 & n20248) | (n20061 & n67029) | (n20248 & n67029);
  assign n51043 = (n20250 & n20252) | (n20250 & n67030) | (n20252 & n67030);
  assign n51044 = n20243 | n50982;
  assign n51045 = (n20243 & n20245) | (n20243 & n51044) | (n20245 & n51044);
  assign n51046 = n20236 | n50984;
  assign n51047 = (n20236 & n20238) | (n20236 & n51046) | (n20238 & n51046);
  assign n67031 = n20229 | n66973;
  assign n67032 = (n20229 & n20231) | (n20229 & n67031) | (n20231 & n67031);
  assign n20264 = n20222 | n20225;
  assign n20265 = n20215 | n20218;
  assign n51048 = n20208 | n20210;
  assign n51049 = (n20069 & n20208) | (n20069 & n51048) | (n20208 & n51048);
  assign n51050 = n20201 | n20203;
  assign n51051 = (n20201 & n50986) | (n20201 & n51050) | (n50986 & n51050);
  assign n51052 = n20194 | n20196;
  assign n51053 = (n20194 & n50988) | (n20194 & n51052) | (n50988 & n51052);
  assign n51054 = n20187 | n20189;
  assign n51055 = (n20187 & n50990) | (n20187 & n51054) | (n50990 & n51054);
  assign n51056 = n20180 | n20182;
  assign n51057 = (n20180 & n50992) | (n20180 & n51056) | (n50992 & n51056);
  assign n51058 = n20173 | n20175;
  assign n51059 = (n20173 & n50994) | (n20173 & n51058) | (n50994 & n51058);
  assign n51060 = n20166 | n20168;
  assign n51061 = (n20166 & n50996) | (n20166 & n51060) | (n50996 & n51060);
  assign n51000 = (n19963 & n50919) | (n19963 & n50999) | (n50919 & n50999);
  assign n51069 = n20138 | n20140;
  assign n67033 = n19949 | n20138;
  assign n67034 = (n20138 & n20140) | (n20138 & n67033) | (n20140 & n67033);
  assign n67035 = (n50972 & n51069) | (n50972 & n67034) | (n51069 & n67034);
  assign n67036 = (n50971 & n51069) | (n50971 & n67034) | (n51069 & n67034);
  assign n67037 = (n66870 & n67035) | (n66870 & n67036) | (n67035 & n67036);
  assign n51074 = n20117 | n20119;
  assign n67038 = n19928 | n20117;
  assign n67039 = (n20117 & n20119) | (n20117 & n67038) | (n20119 & n67038);
  assign n67040 = (n50961 & n51074) | (n50961 & n67039) | (n51074 & n67039);
  assign n67041 = (n50962 & n51074) | (n50962 & n67039) | (n51074 & n67039);
  assign n67042 = (n66875 & n67040) | (n66875 & n67041) | (n67040 & n67041);
  assign n51082 = n20096 | n51019;
  assign n67043 = n20096 | n20098;
  assign n67044 = (n20096 & n66990) | (n20096 & n67043) | (n66990 & n67043);
  assign n67045 = (n51082 & n66882) | (n51082 & n67044) | (n66882 & n67044);
  assign n67046 = (n51082 & n66881) | (n51082 & n67044) | (n66881 & n67044);
  assign n67047 = (n66773 & n67045) | (n66773 & n67046) | (n67045 & n67046);
  assign n20284 = x138 & x176;
  assign n20285 = x137 & x177;
  assign n20286 = n20284 & n20285;
  assign n20287 = n20284 | n20285;
  assign n20288 = ~n20286 & n20287;
  assign n51084 = n20089 | n20091;
  assign n51086 = n20288 & n51084;
  assign n51087 = n20089 & n20288;
  assign n51088 = (n66988 & n51086) | (n66988 & n51087) | (n51086 & n51087);
  assign n51089 = n20288 | n51084;
  assign n51090 = n20089 | n20288;
  assign n51091 = (n66988 & n51089) | (n66988 & n51090) | (n51089 & n51090);
  assign n20291 = ~n51088 & n51091;
  assign n20292 = x136 & x178;
  assign n20293 = n20291 & n20292;
  assign n20294 = n20291 | n20292;
  assign n20295 = ~n20293 & n20294;
  assign n20296 = n67047 & n20295;
  assign n20297 = n67047 | n20295;
  assign n20298 = ~n20296 & n20297;
  assign n20299 = x135 & x179;
  assign n20300 = n20298 & n20299;
  assign n20301 = n20298 | n20299;
  assign n20302 = ~n20300 & n20301;
  assign n67048 = n19914 | n20103;
  assign n67049 = (n20103 & n20105) | (n20103 & n67048) | (n20105 & n67048);
  assign n51092 = n20302 & n67049;
  assign n51079 = n20103 | n20105;
  assign n51093 = n20302 & n51079;
  assign n67050 = (n50949 & n51092) | (n50949 & n51093) | (n51092 & n51093);
  assign n67051 = (n50950 & n51092) | (n50950 & n51093) | (n51092 & n51093);
  assign n67052 = (n50792 & n67050) | (n50792 & n67051) | (n67050 & n67051);
  assign n51095 = n20302 | n67049;
  assign n51096 = n20302 | n51079;
  assign n67053 = (n50949 & n51095) | (n50949 & n51096) | (n51095 & n51096);
  assign n67054 = (n50950 & n51095) | (n50950 & n51096) | (n51095 & n51096);
  assign n67055 = (n50792 & n67053) | (n50792 & n67054) | (n67053 & n67054);
  assign n20305 = ~n67052 & n67055;
  assign n20306 = x134 & x180;
  assign n20307 = n20305 & n20306;
  assign n20308 = n20305 | n20306;
  assign n20309 = ~n20307 & n20308;
  assign n51076 = n20110 | n20112;
  assign n51098 = n20309 & n51076;
  assign n51099 = n20110 & n20309;
  assign n67056 = (n51009 & n51098) | (n51009 & n51099) | (n51098 & n51099);
  assign n67057 = (n51098 & n51099) | (n51098 & n66985) | (n51099 & n66985);
  assign n67058 = (n50869 & n67056) | (n50869 & n67057) | (n67056 & n67057);
  assign n51101 = n20309 | n51076;
  assign n51102 = n20110 | n20309;
  assign n67059 = (n51009 & n51101) | (n51009 & n51102) | (n51101 & n51102);
  assign n67060 = (n51101 & n51102) | (n51101 & n66985) | (n51102 & n66985);
  assign n67061 = (n50869 & n67059) | (n50869 & n67060) | (n67059 & n67060);
  assign n20312 = ~n67058 & n67061;
  assign n20313 = x133 & x181;
  assign n20314 = n20312 & n20313;
  assign n20315 = n20312 | n20313;
  assign n20316 = ~n20314 & n20315;
  assign n20317 = n67042 & n20316;
  assign n20318 = n67042 | n20316;
  assign n20319 = ~n20317 & n20318;
  assign n20320 = x132 & x182;
  assign n20321 = n20319 & n20320;
  assign n20322 = n20319 | n20320;
  assign n20323 = ~n20321 & n20322;
  assign n51071 = n20124 | n20126;
  assign n51104 = n20323 & n51071;
  assign n51105 = n20124 & n20323;
  assign n51106 = (n66983 & n51104) | (n66983 & n51105) | (n51104 & n51105);
  assign n51107 = n20323 | n51071;
  assign n51108 = n20124 | n20323;
  assign n51109 = (n66983 & n51107) | (n66983 & n51108) | (n51107 & n51108);
  assign n20326 = ~n51106 & n51109;
  assign n20327 = x131 & x183;
  assign n20328 = n20326 & n20327;
  assign n20329 = n20326 | n20327;
  assign n20330 = ~n20328 & n20329;
  assign n51110 = n20131 & n20330;
  assign n67062 = (n20330 & n51033) | (n20330 & n51110) | (n51033 & n51110);
  assign n67063 = (n20330 & n51032) | (n20330 & n51110) | (n51032 & n51110);
  assign n67064 = (n66924 & n67062) | (n66924 & n67063) | (n67062 & n67063);
  assign n51112 = n20131 | n20330;
  assign n67065 = n51033 | n51112;
  assign n67066 = n51032 | n51112;
  assign n67067 = (n66924 & n67065) | (n66924 & n67066) | (n67065 & n67066);
  assign n20333 = ~n67064 & n67067;
  assign n20334 = x130 & x184;
  assign n20335 = n20333 & n20334;
  assign n20336 = n20333 | n20334;
  assign n20337 = ~n20335 & n20336;
  assign n20338 = n67037 & n20337;
  assign n20339 = n67037 | n20337;
  assign n20340 = ~n20338 & n20339;
  assign n20341 = x129 & x185;
  assign n20342 = n20340 & n20341;
  assign n20343 = n20340 | n20341;
  assign n20344 = ~n20342 & n20343;
  assign n51066 = n20145 | n20147;
  assign n51114 = n20344 & n51066;
  assign n51115 = n20145 & n20344;
  assign n51116 = (n66978 & n51114) | (n66978 & n51115) | (n51114 & n51115);
  assign n51117 = n20344 | n51066;
  assign n51118 = n20145 | n20344;
  assign n51119 = (n66978 & n51117) | (n66978 & n51118) | (n51117 & n51118);
  assign n20347 = ~n51116 & n51119;
  assign n20348 = x128 & x186;
  assign n20349 = n20347 & n20348;
  assign n20350 = n20347 | n20348;
  assign n20351 = ~n20349 & n20350;
  assign n51064 = n20152 | n20154;
  assign n67068 = n20351 & n51064;
  assign n67069 = n20152 & n20351;
  assign n67070 = (n51000 & n67068) | (n51000 & n67069) | (n67068 & n67069);
  assign n67071 = n20351 | n51064;
  assign n67072 = n20152 | n20351;
  assign n67073 = (n51000 & n67071) | (n51000 & n67072) | (n67071 & n67072);
  assign n20354 = ~n67070 & n67073;
  assign n20355 = x127 & x187;
  assign n20356 = n20354 & n20355;
  assign n20357 = n20354 | n20355;
  assign n20358 = ~n20356 & n20357;
  assign n51062 = n20159 | n20161;
  assign n67074 = n20358 & n51062;
  assign n67075 = n20159 & n20358;
  assign n67076 = (n50998 & n67074) | (n50998 & n67075) | (n67074 & n67075);
  assign n67077 = n20358 | n51062;
  assign n67078 = n20159 | n20358;
  assign n67079 = (n50998 & n67077) | (n50998 & n67078) | (n67077 & n67078);
  assign n20361 = ~n67076 & n67079;
  assign n20362 = x126 & x188;
  assign n20363 = n20361 & n20362;
  assign n20364 = n20361 | n20362;
  assign n20365 = ~n20363 & n20364;
  assign n20366 = n51061 & n20365;
  assign n20367 = n51061 | n20365;
  assign n20368 = ~n20366 & n20367;
  assign n20369 = x125 & x189;
  assign n20370 = n20368 & n20369;
  assign n20371 = n20368 | n20369;
  assign n20372 = ~n20370 & n20371;
  assign n20373 = n51059 & n20372;
  assign n20374 = n51059 | n20372;
  assign n20375 = ~n20373 & n20374;
  assign n20376 = x124 & x190;
  assign n20377 = n20375 & n20376;
  assign n20378 = n20375 | n20376;
  assign n20379 = ~n20377 & n20378;
  assign n20380 = n51057 & n20379;
  assign n20381 = n51057 | n20379;
  assign n20382 = ~n20380 & n20381;
  assign n20383 = x123 & x191;
  assign n20384 = n20382 & n20383;
  assign n20385 = n20382 | n20383;
  assign n20386 = ~n20384 & n20385;
  assign n20387 = n51055 & n20386;
  assign n20388 = n51055 | n20386;
  assign n20389 = ~n20387 & n20388;
  assign n20390 = x122 & x192;
  assign n20391 = n20389 & n20390;
  assign n20392 = n20389 | n20390;
  assign n20393 = ~n20391 & n20392;
  assign n20394 = n51053 & n20393;
  assign n20395 = n51053 | n20393;
  assign n20396 = ~n20394 & n20395;
  assign n20397 = x121 & x193;
  assign n20398 = n20396 & n20397;
  assign n20399 = n20396 | n20397;
  assign n20400 = ~n20398 & n20399;
  assign n20401 = n51051 & n20400;
  assign n20402 = n51051 | n20400;
  assign n20403 = ~n20401 & n20402;
  assign n20404 = x120 & x194;
  assign n20405 = n20403 & n20404;
  assign n20406 = n20403 | n20404;
  assign n20407 = ~n20405 & n20406;
  assign n20408 = n51049 & n20407;
  assign n20409 = n51049 | n20407;
  assign n20410 = ~n20408 & n20409;
  assign n20411 = x119 & x195;
  assign n20412 = n20410 & n20411;
  assign n20413 = n20410 | n20411;
  assign n20414 = ~n20412 & n20413;
  assign n20415 = n20265 & n20414;
  assign n20416 = n20265 | n20414;
  assign n20417 = ~n20415 & n20416;
  assign n20418 = x118 & x196;
  assign n20419 = n20417 & n20418;
  assign n20420 = n20417 | n20418;
  assign n20421 = ~n20419 & n20420;
  assign n20422 = n20264 & n20421;
  assign n20423 = n20264 | n20421;
  assign n20424 = ~n20422 & n20423;
  assign n20425 = x117 & x197;
  assign n20426 = n20424 & n20425;
  assign n20427 = n20424 | n20425;
  assign n20428 = ~n20426 & n20427;
  assign n20429 = n67032 & n20428;
  assign n20430 = n67032 | n20428;
  assign n20431 = ~n20429 & n20430;
  assign n20432 = x116 & x198;
  assign n20433 = n20431 & n20432;
  assign n20434 = n20431 | n20432;
  assign n20435 = ~n20433 & n20434;
  assign n20436 = n51047 & n20435;
  assign n20437 = n51047 | n20435;
  assign n20438 = ~n20436 & n20437;
  assign n20439 = x115 & x199;
  assign n20440 = n20438 & n20439;
  assign n20441 = n20438 | n20439;
  assign n20442 = ~n20440 & n20441;
  assign n20443 = n51045 & n20442;
  assign n20444 = n51045 | n20442;
  assign n20445 = ~n20443 & n20444;
  assign n20446 = x114 & x200;
  assign n20447 = n20445 & n20446;
  assign n20448 = n20445 | n20446;
  assign n20449 = ~n20447 & n20448;
  assign n20450 = n51043 & n20449;
  assign n20451 = n51043 | n20449;
  assign n20452 = ~n20450 & n20451;
  assign n20453 = x113 & x201;
  assign n20454 = n20452 & n20453;
  assign n20455 = n20452 | n20453;
  assign n20456 = ~n20454 & n20455;
  assign n20457 = n20257 & n20456;
  assign n20458 = n20257 | n20456;
  assign n20459 = ~n20457 & n20458;
  assign n20460 = x112 & x202;
  assign n20461 = n20459 & n20460;
  assign n20462 = n20459 | n20460;
  assign n20463 = ~n20461 & n20462;
  assign n67080 = n20257 | n20453;
  assign n67081 = (n20257 & n20452) | (n20257 & n67080) | (n20452 & n67080);
  assign n51121 = (n20454 & n20456) | (n20454 & n67081) | (n20456 & n67081);
  assign n51122 = n20447 | n51043;
  assign n51123 = (n20447 & n20449) | (n20447 & n51122) | (n20449 & n51122);
  assign n51124 = n20440 | n51045;
  assign n51125 = (n20440 & n20442) | (n20440 & n51124) | (n20442 & n51124);
  assign n51126 = n20433 | n51047;
  assign n51127 = (n20433 & n20435) | (n20433 & n51126) | (n20435 & n51126);
  assign n67082 = n20426 | n67032;
  assign n67083 = (n20426 & n20428) | (n20426 & n67082) | (n20428 & n67082);
  assign n20469 = n20419 | n20422;
  assign n51128 = n20412 | n20414;
  assign n51129 = (n20265 & n20412) | (n20265 & n51128) | (n20412 & n51128);
  assign n51130 = n20405 | n20407;
  assign n51131 = (n20405 & n51049) | (n20405 & n51130) | (n51049 & n51130);
  assign n51132 = n20398 | n20400;
  assign n51133 = (n20398 & n51051) | (n20398 & n51132) | (n51051 & n51132);
  assign n51134 = n20391 | n20393;
  assign n51135 = (n20391 & n51053) | (n20391 & n51134) | (n51053 & n51134);
  assign n51136 = n20384 | n20386;
  assign n51137 = (n20384 & n51055) | (n20384 & n51136) | (n51055 & n51136);
  assign n51138 = n20377 | n20379;
  assign n51139 = (n20377 & n51057) | (n20377 & n51138) | (n51057 & n51138);
  assign n51140 = n20370 | n20372;
  assign n51141 = (n20370 & n51059) | (n20370 & n51140) | (n51059 & n51140);
  assign n51063 = (n20159 & n50998) | (n20159 & n51062) | (n50998 & n51062);
  assign n51065 = (n20152 & n51000) | (n20152 & n51064) | (n51000 & n51064);
  assign n51151 = n20328 | n20330;
  assign n67084 = n20131 | n20328;
  assign n67085 = (n20328 & n20330) | (n20328 & n67084) | (n20330 & n67084);
  assign n67086 = (n51033 & n51151) | (n51033 & n67085) | (n51151 & n67085);
  assign n67087 = (n51032 & n51151) | (n51032 & n67085) | (n51151 & n67085);
  assign n67088 = (n66924 & n67086) | (n66924 & n67087) | (n67086 & n67087);
  assign n67089 = n20307 | n20309;
  assign n67090 = (n20307 & n51076) | (n20307 & n67089) | (n51076 & n67089);
  assign n67091 = n20110 | n20307;
  assign n67092 = (n20307 & n20309) | (n20307 & n67091) | (n20309 & n67091);
  assign n67093 = (n51009 & n67090) | (n51009 & n67092) | (n67090 & n67092);
  assign n67094 = (n66985 & n67090) | (n66985 & n67092) | (n67090 & n67092);
  assign n67095 = (n50869 & n67093) | (n50869 & n67094) | (n67093 & n67094);
  assign n51158 = n20300 | n51092;
  assign n51159 = n20300 | n51093;
  assign n67096 = (n50949 & n51158) | (n50949 & n51159) | (n51158 & n51159);
  assign n67097 = (n50950 & n51158) | (n50950 & n51159) | (n51158 & n51159);
  assign n67098 = (n50792 & n67096) | (n50792 & n67097) | (n67096 & n67097);
  assign n20489 = x139 & x176;
  assign n20490 = x138 & x177;
  assign n20491 = n20489 & n20490;
  assign n20492 = n20489 | n20490;
  assign n20493 = ~n20491 & n20492;
  assign n67099 = n20286 | n20288;
  assign n67100 = (n20286 & n51084) | (n20286 & n67099) | (n51084 & n67099);
  assign n51166 = n20493 & n67100;
  assign n67101 = n20089 | n20286;
  assign n67102 = (n20286 & n20288) | (n20286 & n67101) | (n20288 & n67101);
  assign n51167 = n20493 & n67102;
  assign n51168 = (n66988 & n51166) | (n66988 & n51167) | (n51166 & n51167);
  assign n51169 = n20493 | n67100;
  assign n51170 = n20493 | n67102;
  assign n51171 = (n66988 & n51169) | (n66988 & n51170) | (n51169 & n51170);
  assign n20496 = ~n51168 & n51171;
  assign n20497 = x137 & x178;
  assign n20498 = n20496 & n20497;
  assign n20499 = n20496 | n20497;
  assign n20500 = ~n20498 & n20499;
  assign n51161 = n20293 | n20295;
  assign n51172 = n20500 & n51161;
  assign n51173 = n20293 & n20500;
  assign n51174 = (n67047 & n51172) | (n67047 & n51173) | (n51172 & n51173);
  assign n51175 = n20500 | n51161;
  assign n51176 = n20293 | n20500;
  assign n51177 = (n67047 & n51175) | (n67047 & n51176) | (n51175 & n51176);
  assign n20503 = ~n51174 & n51177;
  assign n20504 = x136 & x179;
  assign n20505 = n20503 & n20504;
  assign n20506 = n20503 | n20504;
  assign n20507 = ~n20505 & n20506;
  assign n20508 = n67098 & n20507;
  assign n20509 = n67098 | n20507;
  assign n20510 = ~n20508 & n20509;
  assign n20511 = x135 & x180;
  assign n20512 = n20510 & n20511;
  assign n20513 = n20510 | n20511;
  assign n20514 = ~n20512 & n20513;
  assign n20515 = n67095 & n20514;
  assign n20516 = n67095 | n20514;
  assign n20517 = ~n20515 & n20516;
  assign n20518 = x134 & x181;
  assign n20519 = n20517 & n20518;
  assign n20520 = n20517 | n20518;
  assign n20521 = ~n20519 & n20520;
  assign n51153 = n20314 | n20316;
  assign n51178 = n20521 & n51153;
  assign n51179 = n20314 & n20521;
  assign n51180 = (n67042 & n51178) | (n67042 & n51179) | (n51178 & n51179);
  assign n51181 = n20521 | n51153;
  assign n51182 = n20314 | n20521;
  assign n51183 = (n67042 & n51181) | (n67042 & n51182) | (n51181 & n51182);
  assign n20524 = ~n51180 & n51183;
  assign n20525 = x133 & x182;
  assign n20526 = n20524 & n20525;
  assign n20527 = n20524 | n20525;
  assign n20528 = ~n20526 & n20527;
  assign n51184 = n20321 & n20528;
  assign n67103 = (n20528 & n51105) | (n20528 & n51184) | (n51105 & n51184);
  assign n67104 = (n20528 & n51104) | (n20528 & n51184) | (n51104 & n51184);
  assign n67105 = (n66983 & n67103) | (n66983 & n67104) | (n67103 & n67104);
  assign n51186 = n20321 | n20528;
  assign n67106 = n51105 | n51186;
  assign n67107 = n51104 | n51186;
  assign n67108 = (n66983 & n67106) | (n66983 & n67107) | (n67106 & n67107);
  assign n20531 = ~n67105 & n67108;
  assign n20532 = x132 & x183;
  assign n20533 = n20531 & n20532;
  assign n20534 = n20531 | n20532;
  assign n20535 = ~n20533 & n20534;
  assign n20536 = n67088 & n20535;
  assign n20537 = n67088 | n20535;
  assign n20538 = ~n20536 & n20537;
  assign n20539 = x131 & x184;
  assign n20540 = n20538 & n20539;
  assign n20541 = n20538 | n20539;
  assign n20542 = ~n20540 & n20541;
  assign n51148 = n20335 | n20337;
  assign n51188 = n20542 & n51148;
  assign n51189 = n20335 & n20542;
  assign n51190 = (n67037 & n51188) | (n67037 & n51189) | (n51188 & n51189);
  assign n51191 = n20542 | n51148;
  assign n51192 = n20335 | n20542;
  assign n51193 = (n67037 & n51191) | (n67037 & n51192) | (n51191 & n51192);
  assign n20545 = ~n51190 & n51193;
  assign n20546 = x130 & x185;
  assign n20547 = n20545 & n20546;
  assign n20548 = n20545 | n20546;
  assign n20549 = ~n20547 & n20548;
  assign n51194 = n20342 & n20549;
  assign n67109 = (n20549 & n51115) | (n20549 & n51194) | (n51115 & n51194);
  assign n67110 = (n20549 & n51114) | (n20549 & n51194) | (n51114 & n51194);
  assign n67111 = (n66978 & n67109) | (n66978 & n67110) | (n67109 & n67110);
  assign n51196 = n20342 | n20549;
  assign n67112 = n51115 | n51196;
  assign n67113 = n51114 | n51196;
  assign n67114 = (n66978 & n67112) | (n66978 & n67113) | (n67112 & n67113);
  assign n20552 = ~n67111 & n67114;
  assign n20553 = x129 & x186;
  assign n20554 = n20552 & n20553;
  assign n20555 = n20552 | n20553;
  assign n20556 = ~n20554 & n20555;
  assign n51146 = n20349 | n20351;
  assign n51198 = n20556 & n51146;
  assign n51199 = n20349 & n20556;
  assign n51200 = (n51065 & n51198) | (n51065 & n51199) | (n51198 & n51199);
  assign n51201 = n20556 | n51146;
  assign n51202 = n20349 | n20556;
  assign n51203 = (n51065 & n51201) | (n51065 & n51202) | (n51201 & n51202);
  assign n20559 = ~n51200 & n51203;
  assign n20560 = x128 & x187;
  assign n20561 = n20559 & n20560;
  assign n20562 = n20559 | n20560;
  assign n20563 = ~n20561 & n20562;
  assign n51144 = n20356 | n20358;
  assign n67115 = n20563 & n51144;
  assign n67116 = n20356 & n20563;
  assign n67117 = (n51063 & n67115) | (n51063 & n67116) | (n67115 & n67116);
  assign n67118 = n20563 | n51144;
  assign n67119 = n20356 | n20563;
  assign n67120 = (n51063 & n67118) | (n51063 & n67119) | (n67118 & n67119);
  assign n20566 = ~n67117 & n67120;
  assign n20567 = x127 & x188;
  assign n20568 = n20566 & n20567;
  assign n20569 = n20566 | n20567;
  assign n20570 = ~n20568 & n20569;
  assign n51142 = n20363 | n20365;
  assign n67121 = n20570 & n51142;
  assign n67122 = n20363 & n20570;
  assign n67123 = (n51061 & n67121) | (n51061 & n67122) | (n67121 & n67122);
  assign n67124 = n20570 | n51142;
  assign n67125 = n20363 | n20570;
  assign n67126 = (n51061 & n67124) | (n51061 & n67125) | (n67124 & n67125);
  assign n20573 = ~n67123 & n67126;
  assign n20574 = x126 & x189;
  assign n20575 = n20573 & n20574;
  assign n20576 = n20573 | n20574;
  assign n20577 = ~n20575 & n20576;
  assign n20578 = n51141 & n20577;
  assign n20579 = n51141 | n20577;
  assign n20580 = ~n20578 & n20579;
  assign n20581 = x125 & x190;
  assign n20582 = n20580 & n20581;
  assign n20583 = n20580 | n20581;
  assign n20584 = ~n20582 & n20583;
  assign n20585 = n51139 & n20584;
  assign n20586 = n51139 | n20584;
  assign n20587 = ~n20585 & n20586;
  assign n20588 = x124 & x191;
  assign n20589 = n20587 & n20588;
  assign n20590 = n20587 | n20588;
  assign n20591 = ~n20589 & n20590;
  assign n20592 = n51137 & n20591;
  assign n20593 = n51137 | n20591;
  assign n20594 = ~n20592 & n20593;
  assign n20595 = x123 & x192;
  assign n20596 = n20594 & n20595;
  assign n20597 = n20594 | n20595;
  assign n20598 = ~n20596 & n20597;
  assign n20599 = n51135 & n20598;
  assign n20600 = n51135 | n20598;
  assign n20601 = ~n20599 & n20600;
  assign n20602 = x122 & x193;
  assign n20603 = n20601 & n20602;
  assign n20604 = n20601 | n20602;
  assign n20605 = ~n20603 & n20604;
  assign n20606 = n51133 & n20605;
  assign n20607 = n51133 | n20605;
  assign n20608 = ~n20606 & n20607;
  assign n20609 = x121 & x194;
  assign n20610 = n20608 & n20609;
  assign n20611 = n20608 | n20609;
  assign n20612 = ~n20610 & n20611;
  assign n20613 = n51131 & n20612;
  assign n20614 = n51131 | n20612;
  assign n20615 = ~n20613 & n20614;
  assign n20616 = x120 & x195;
  assign n20617 = n20615 & n20616;
  assign n20618 = n20615 | n20616;
  assign n20619 = ~n20617 & n20618;
  assign n20620 = n51129 & n20619;
  assign n20621 = n51129 | n20619;
  assign n20622 = ~n20620 & n20621;
  assign n20623 = x119 & x196;
  assign n20624 = n20622 & n20623;
  assign n20625 = n20622 | n20623;
  assign n20626 = ~n20624 & n20625;
  assign n20627 = n20469 & n20626;
  assign n20628 = n20469 | n20626;
  assign n20629 = ~n20627 & n20628;
  assign n20630 = x118 & x197;
  assign n20631 = n20629 & n20630;
  assign n20632 = n20629 | n20630;
  assign n20633 = ~n20631 & n20632;
  assign n20634 = n67083 & n20633;
  assign n20635 = n67083 | n20633;
  assign n20636 = ~n20634 & n20635;
  assign n20637 = x117 & x198;
  assign n20638 = n20636 & n20637;
  assign n20639 = n20636 | n20637;
  assign n20640 = ~n20638 & n20639;
  assign n20641 = n51127 & n20640;
  assign n20642 = n51127 | n20640;
  assign n20643 = ~n20641 & n20642;
  assign n20644 = x116 & x199;
  assign n20645 = n20643 & n20644;
  assign n20646 = n20643 | n20644;
  assign n20647 = ~n20645 & n20646;
  assign n20648 = n51125 & n20647;
  assign n20649 = n51125 | n20647;
  assign n20650 = ~n20648 & n20649;
  assign n20651 = x115 & x200;
  assign n20652 = n20650 & n20651;
  assign n20653 = n20650 | n20651;
  assign n20654 = ~n20652 & n20653;
  assign n20655 = n51123 & n20654;
  assign n20656 = n51123 | n20654;
  assign n20657 = ~n20655 & n20656;
  assign n20658 = x114 & x201;
  assign n20659 = n20657 & n20658;
  assign n20660 = n20657 | n20658;
  assign n20661 = ~n20659 & n20660;
  assign n20662 = n51121 & n20661;
  assign n20663 = n51121 | n20661;
  assign n20664 = ~n20662 & n20663;
  assign n20665 = x113 & x202;
  assign n20666 = n20664 & n20665;
  assign n20667 = n20664 | n20665;
  assign n20668 = ~n20666 & n20667;
  assign n20669 = n20461 & n20668;
  assign n20670 = n20461 | n20668;
  assign n20671 = ~n20669 & n20670;
  assign n20672 = x112 & x203;
  assign n20673 = n20671 & n20672;
  assign n20674 = n20671 | n20672;
  assign n20675 = ~n20673 & n20674;
  assign n67127 = n20461 | n20665;
  assign n67128 = (n20461 & n20664) | (n20461 & n67127) | (n20664 & n67127);
  assign n51205 = (n20666 & n20668) | (n20666 & n67128) | (n20668 & n67128);
  assign n51206 = n20659 | n51121;
  assign n51207 = (n20659 & n20661) | (n20659 & n51206) | (n20661 & n51206);
  assign n51208 = n20652 | n51123;
  assign n51209 = (n20652 & n20654) | (n20652 & n51208) | (n20654 & n51208);
  assign n51210 = n20645 | n51125;
  assign n51211 = (n20645 & n20647) | (n20645 & n51210) | (n20647 & n51210);
  assign n51212 = n20638 | n51127;
  assign n51213 = (n20638 & n20640) | (n20638 & n51212) | (n20640 & n51212);
  assign n67129 = n20631 | n67083;
  assign n67130 = (n20631 & n20633) | (n20631 & n67129) | (n20633 & n67129);
  assign n51214 = n20624 | n20626;
  assign n51215 = (n20469 & n20624) | (n20469 & n51214) | (n20624 & n51214);
  assign n51216 = n20617 | n20619;
  assign n51217 = (n20617 & n51129) | (n20617 & n51216) | (n51129 & n51216);
  assign n51218 = n20610 | n20612;
  assign n51219 = (n20610 & n51131) | (n20610 & n51218) | (n51131 & n51218);
  assign n51220 = n20603 | n20605;
  assign n51221 = (n20603 & n51133) | (n20603 & n51220) | (n51133 & n51220);
  assign n51222 = n20596 | n20598;
  assign n51223 = (n20596 & n51135) | (n20596 & n51222) | (n51135 & n51222);
  assign n51224 = n20589 | n20591;
  assign n51225 = (n20589 & n51137) | (n20589 & n51224) | (n51137 & n51224);
  assign n51226 = n20582 | n20584;
  assign n51227 = (n20582 & n51139) | (n20582 & n51226) | (n51139 & n51226);
  assign n51143 = (n20363 & n51061) | (n20363 & n51142) | (n51061 & n51142);
  assign n51145 = (n20356 & n51063) | (n20356 & n51144) | (n51063 & n51144);
  assign n51235 = n20547 | n20549;
  assign n67131 = n20342 | n20547;
  assign n67132 = (n20547 & n20549) | (n20547 & n67131) | (n20549 & n67131);
  assign n67133 = (n51115 & n51235) | (n51115 & n67132) | (n51235 & n67132);
  assign n67134 = (n51114 & n51235) | (n51114 & n67132) | (n51235 & n67132);
  assign n67135 = (n66978 & n67133) | (n66978 & n67134) | (n67133 & n67134);
  assign n51240 = n20526 | n20528;
  assign n67136 = n20321 | n20526;
  assign n67137 = (n20526 & n20528) | (n20526 & n67136) | (n20528 & n67136);
  assign n67138 = (n51105 & n51240) | (n51105 & n67137) | (n51240 & n67137);
  assign n67139 = (n51104 & n51240) | (n51104 & n67137) | (n51240 & n67137);
  assign n67140 = (n66983 & n67138) | (n66983 & n67139) | (n67138 & n67139);
  assign n67141 = n20314 | n20519;
  assign n67142 = (n20519 & n20521) | (n20519 & n67141) | (n20521 & n67141);
  assign n51243 = n20519 | n51178;
  assign n51244 = (n67042 & n67142) | (n67042 & n51243) | (n67142 & n51243);
  assign n20702 = x140 & x176;
  assign n20703 = x139 & x177;
  assign n20704 = n20702 & n20703;
  assign n20705 = n20702 | n20703;
  assign n20706 = ~n20704 & n20705;
  assign n67143 = n20491 | n20493;
  assign n67145 = n20706 & n67143;
  assign n67146 = n20491 & n20706;
  assign n67147 = (n67100 & n67145) | (n67100 & n67146) | (n67145 & n67146);
  assign n67148 = (n20491 & n67102) | (n20491 & n67143) | (n67102 & n67143);
  assign n51256 = n20706 & n67148;
  assign n51257 = (n66988 & n67147) | (n66988 & n51256) | (n67147 & n51256);
  assign n67149 = n20706 | n67143;
  assign n67150 = n20491 | n20706;
  assign n67151 = (n67100 & n67149) | (n67100 & n67150) | (n67149 & n67150);
  assign n51259 = n20706 | n67148;
  assign n51260 = (n66988 & n67151) | (n66988 & n51259) | (n67151 & n51259);
  assign n20709 = ~n51257 & n51260;
  assign n20710 = x138 & x178;
  assign n20711 = n20709 & n20710;
  assign n20712 = n20709 | n20710;
  assign n20713 = ~n20711 & n20712;
  assign n67152 = n20498 | n20500;
  assign n67153 = (n20498 & n51161) | (n20498 & n67152) | (n51161 & n67152);
  assign n51261 = n20713 & n67153;
  assign n67154 = n20293 | n20498;
  assign n67155 = (n20498 & n20500) | (n20498 & n67154) | (n20500 & n67154);
  assign n51262 = n20713 & n67155;
  assign n51263 = (n67047 & n51261) | (n67047 & n51262) | (n51261 & n51262);
  assign n51264 = n20713 | n67153;
  assign n51265 = n20713 | n67155;
  assign n51266 = (n67047 & n51264) | (n67047 & n51265) | (n51264 & n51265);
  assign n20716 = ~n51263 & n51266;
  assign n20717 = x137 & x179;
  assign n20718 = n20716 & n20717;
  assign n20719 = n20716 | n20717;
  assign n20720 = ~n20718 & n20719;
  assign n51247 = n20505 | n20507;
  assign n51267 = n20720 & n51247;
  assign n51268 = n20505 & n20720;
  assign n51269 = (n67098 & n51267) | (n67098 & n51268) | (n51267 & n51268);
  assign n51270 = n20720 | n51247;
  assign n51271 = n20505 | n20720;
  assign n51272 = (n67098 & n51270) | (n67098 & n51271) | (n51270 & n51271);
  assign n20723 = ~n51269 & n51272;
  assign n20724 = x136 & x180;
  assign n20725 = n20723 & n20724;
  assign n20726 = n20723 | n20724;
  assign n20727 = ~n20725 & n20726;
  assign n51245 = n20512 | n20514;
  assign n51273 = n20727 & n51245;
  assign n51274 = n20512 & n20727;
  assign n51275 = (n67095 & n51273) | (n67095 & n51274) | (n51273 & n51274);
  assign n51276 = n20727 | n51245;
  assign n51277 = n20512 | n20727;
  assign n51278 = (n67095 & n51276) | (n67095 & n51277) | (n51276 & n51277);
  assign n20730 = ~n51275 & n51278;
  assign n20731 = x135 & x181;
  assign n20732 = n20730 & n20731;
  assign n20733 = n20730 | n20731;
  assign n20734 = ~n20732 & n20733;
  assign n20735 = n51244 & n20734;
  assign n20736 = n51244 | n20734;
  assign n20737 = ~n20735 & n20736;
  assign n20738 = x134 & x182;
  assign n20739 = n20737 & n20738;
  assign n20740 = n20737 | n20738;
  assign n20741 = ~n20739 & n20740;
  assign n20742 = n67140 & n20741;
  assign n20743 = n67140 | n20741;
  assign n20744 = ~n20742 & n20743;
  assign n20745 = x133 & x183;
  assign n20746 = n20744 & n20745;
  assign n20747 = n20744 | n20745;
  assign n20748 = ~n20746 & n20747;
  assign n51237 = n20533 | n20535;
  assign n51279 = n20748 & n51237;
  assign n51280 = n20533 & n20748;
  assign n51281 = (n67088 & n51279) | (n67088 & n51280) | (n51279 & n51280);
  assign n51282 = n20748 | n51237;
  assign n51283 = n20533 | n20748;
  assign n51284 = (n67088 & n51282) | (n67088 & n51283) | (n51282 & n51283);
  assign n20751 = ~n51281 & n51284;
  assign n20752 = x132 & x184;
  assign n20753 = n20751 & n20752;
  assign n20754 = n20751 | n20752;
  assign n20755 = ~n20753 & n20754;
  assign n51285 = n20540 & n20755;
  assign n67156 = (n20755 & n51189) | (n20755 & n51285) | (n51189 & n51285);
  assign n67157 = (n20755 & n51188) | (n20755 & n51285) | (n51188 & n51285);
  assign n67158 = (n67037 & n67156) | (n67037 & n67157) | (n67156 & n67157);
  assign n51287 = n20540 | n20755;
  assign n67159 = n51189 | n51287;
  assign n67160 = n51188 | n51287;
  assign n67161 = (n67037 & n67159) | (n67037 & n67160) | (n67159 & n67160);
  assign n20758 = ~n67158 & n67161;
  assign n20759 = x131 & x185;
  assign n20760 = n20758 & n20759;
  assign n20761 = n20758 | n20759;
  assign n20762 = ~n20760 & n20761;
  assign n20763 = n67135 & n20762;
  assign n20764 = n67135 | n20762;
  assign n20765 = ~n20763 & n20764;
  assign n20766 = x130 & x186;
  assign n20767 = n20765 & n20766;
  assign n20768 = n20765 | n20766;
  assign n20769 = ~n20767 & n20768;
  assign n51289 = n20554 & n20769;
  assign n67162 = (n20769 & n51198) | (n20769 & n51289) | (n51198 & n51289);
  assign n67163 = (n20769 & n51199) | (n20769 & n51289) | (n51199 & n51289);
  assign n67164 = (n51065 & n67162) | (n51065 & n67163) | (n67162 & n67163);
  assign n51291 = n20554 | n20769;
  assign n67165 = n51198 | n51291;
  assign n67166 = n51199 | n51291;
  assign n67167 = (n51065 & n67165) | (n51065 & n67166) | (n67165 & n67166);
  assign n20772 = ~n67164 & n67167;
  assign n20773 = x129 & x187;
  assign n20774 = n20772 & n20773;
  assign n20775 = n20772 | n20773;
  assign n20776 = ~n20774 & n20775;
  assign n51232 = n20561 | n20563;
  assign n51293 = n20776 & n51232;
  assign n51294 = n20561 & n20776;
  assign n51295 = (n51145 & n51293) | (n51145 & n51294) | (n51293 & n51294);
  assign n51296 = n20776 | n51232;
  assign n51297 = n20561 | n20776;
  assign n51298 = (n51145 & n51296) | (n51145 & n51297) | (n51296 & n51297);
  assign n20779 = ~n51295 & n51298;
  assign n20780 = x128 & x188;
  assign n20781 = n20779 & n20780;
  assign n20782 = n20779 | n20780;
  assign n20783 = ~n20781 & n20782;
  assign n51230 = n20568 | n20570;
  assign n67168 = n20783 & n51230;
  assign n67169 = n20568 & n20783;
  assign n67170 = (n51143 & n67168) | (n51143 & n67169) | (n67168 & n67169);
  assign n67171 = n20783 | n51230;
  assign n67172 = n20568 | n20783;
  assign n67173 = (n51143 & n67171) | (n51143 & n67172) | (n67171 & n67172);
  assign n20786 = ~n67170 & n67173;
  assign n20787 = x127 & x189;
  assign n20788 = n20786 & n20787;
  assign n20789 = n20786 | n20787;
  assign n20790 = ~n20788 & n20789;
  assign n51228 = n20575 | n20577;
  assign n67174 = n20790 & n51228;
  assign n67175 = n20575 & n20790;
  assign n67176 = (n51141 & n67174) | (n51141 & n67175) | (n67174 & n67175);
  assign n67177 = n20790 | n51228;
  assign n67178 = n20575 | n20790;
  assign n67179 = (n51141 & n67177) | (n51141 & n67178) | (n67177 & n67178);
  assign n20793 = ~n67176 & n67179;
  assign n20794 = x126 & x190;
  assign n20795 = n20793 & n20794;
  assign n20796 = n20793 | n20794;
  assign n20797 = ~n20795 & n20796;
  assign n20798 = n51227 & n20797;
  assign n20799 = n51227 | n20797;
  assign n20800 = ~n20798 & n20799;
  assign n20801 = x125 & x191;
  assign n20802 = n20800 & n20801;
  assign n20803 = n20800 | n20801;
  assign n20804 = ~n20802 & n20803;
  assign n20805 = n51225 & n20804;
  assign n20806 = n51225 | n20804;
  assign n20807 = ~n20805 & n20806;
  assign n20808 = x124 & x192;
  assign n20809 = n20807 & n20808;
  assign n20810 = n20807 | n20808;
  assign n20811 = ~n20809 & n20810;
  assign n20812 = n51223 & n20811;
  assign n20813 = n51223 | n20811;
  assign n20814 = ~n20812 & n20813;
  assign n20815 = x123 & x193;
  assign n20816 = n20814 & n20815;
  assign n20817 = n20814 | n20815;
  assign n20818 = ~n20816 & n20817;
  assign n20819 = n51221 & n20818;
  assign n20820 = n51221 | n20818;
  assign n20821 = ~n20819 & n20820;
  assign n20822 = x122 & x194;
  assign n20823 = n20821 & n20822;
  assign n20824 = n20821 | n20822;
  assign n20825 = ~n20823 & n20824;
  assign n20826 = n51219 & n20825;
  assign n20827 = n51219 | n20825;
  assign n20828 = ~n20826 & n20827;
  assign n20829 = x121 & x195;
  assign n20830 = n20828 & n20829;
  assign n20831 = n20828 | n20829;
  assign n20832 = ~n20830 & n20831;
  assign n20833 = n51217 & n20832;
  assign n20834 = n51217 | n20832;
  assign n20835 = ~n20833 & n20834;
  assign n20836 = x120 & x196;
  assign n20837 = n20835 & n20836;
  assign n20838 = n20835 | n20836;
  assign n20839 = ~n20837 & n20838;
  assign n20840 = n51215 & n20839;
  assign n20841 = n51215 | n20839;
  assign n20842 = ~n20840 & n20841;
  assign n20843 = x119 & x197;
  assign n20844 = n20842 & n20843;
  assign n20845 = n20842 | n20843;
  assign n20846 = ~n20844 & n20845;
  assign n20847 = n67130 & n20846;
  assign n20848 = n67130 | n20846;
  assign n20849 = ~n20847 & n20848;
  assign n20850 = x118 & x198;
  assign n20851 = n20849 & n20850;
  assign n20852 = n20849 | n20850;
  assign n20853 = ~n20851 & n20852;
  assign n20854 = n51213 & n20853;
  assign n20855 = n51213 | n20853;
  assign n20856 = ~n20854 & n20855;
  assign n20857 = x117 & x199;
  assign n20858 = n20856 & n20857;
  assign n20859 = n20856 | n20857;
  assign n20860 = ~n20858 & n20859;
  assign n20861 = n51211 & n20860;
  assign n20862 = n51211 | n20860;
  assign n20863 = ~n20861 & n20862;
  assign n20864 = x116 & x200;
  assign n20865 = n20863 & n20864;
  assign n20866 = n20863 | n20864;
  assign n20867 = ~n20865 & n20866;
  assign n20868 = n51209 & n20867;
  assign n20869 = n51209 | n20867;
  assign n20870 = ~n20868 & n20869;
  assign n20871 = x115 & x201;
  assign n20872 = n20870 & n20871;
  assign n20873 = n20870 | n20871;
  assign n20874 = ~n20872 & n20873;
  assign n20875 = n51207 & n20874;
  assign n20876 = n51207 | n20874;
  assign n20877 = ~n20875 & n20876;
  assign n20878 = x114 & x202;
  assign n20879 = n20877 & n20878;
  assign n20880 = n20877 | n20878;
  assign n20881 = ~n20879 & n20880;
  assign n20882 = n51205 & n20881;
  assign n20883 = n51205 | n20881;
  assign n20884 = ~n20882 & n20883;
  assign n20885 = x113 & x203;
  assign n20886 = n20884 & n20885;
  assign n20887 = n20884 | n20885;
  assign n20888 = ~n20886 & n20887;
  assign n20889 = n20673 & n20888;
  assign n20890 = n20673 | n20888;
  assign n20891 = ~n20889 & n20890;
  assign n20892 = x112 & x204;
  assign n20893 = n20891 & n20892;
  assign n20894 = n20891 | n20892;
  assign n20895 = ~n20893 & n20894;
  assign n51299 = n20673 | n20886;
  assign n51300 = (n20886 & n20888) | (n20886 & n51299) | (n20888 & n51299);
  assign n51301 = n20879 | n51205;
  assign n51302 = (n20879 & n20881) | (n20879 & n51301) | (n20881 & n51301);
  assign n51303 = n20872 | n51207;
  assign n51304 = (n20872 & n20874) | (n20872 & n51303) | (n20874 & n51303);
  assign n51305 = n20865 | n51209;
  assign n51306 = (n20865 & n20867) | (n20865 & n51305) | (n20867 & n51305);
  assign n51307 = n20858 | n51211;
  assign n51308 = (n20858 & n20860) | (n20858 & n51307) | (n20860 & n51307);
  assign n51309 = n20851 | n51213;
  assign n51310 = (n20851 & n20853) | (n20851 & n51309) | (n20853 & n51309);
  assign n51311 = n20844 | n20846;
  assign n51312 = (n67130 & n20844) | (n67130 & n51311) | (n20844 & n51311);
  assign n51313 = n20837 | n20839;
  assign n51314 = (n20837 & n51215) | (n20837 & n51313) | (n51215 & n51313);
  assign n51315 = n20830 | n20832;
  assign n51316 = (n20830 & n51217) | (n20830 & n51315) | (n51217 & n51315);
  assign n51317 = n20823 | n20825;
  assign n51318 = (n20823 & n51219) | (n20823 & n51317) | (n51219 & n51317);
  assign n51319 = n20816 | n20818;
  assign n51320 = (n20816 & n51221) | (n20816 & n51319) | (n51221 & n51319);
  assign n51321 = n20809 | n20811;
  assign n51322 = (n20809 & n51223) | (n20809 & n51321) | (n51223 & n51321);
  assign n51323 = n20802 | n20804;
  assign n51324 = (n20802 & n51225) | (n20802 & n51323) | (n51225 & n51323);
  assign n51229 = (n20575 & n51141) | (n20575 & n51228) | (n51141 & n51228);
  assign n51231 = (n20568 & n51143) | (n20568 & n51230) | (n51143 & n51230);
  assign n51334 = n20753 | n20755;
  assign n67180 = n20540 | n20753;
  assign n67181 = (n20753 & n20755) | (n20753 & n67180) | (n20755 & n67180);
  assign n67182 = (n51189 & n51334) | (n51189 & n67181) | (n51334 & n67181);
  assign n67183 = (n51188 & n51334) | (n51188 & n67181) | (n51334 & n67181);
  assign n67184 = (n67037 & n67182) | (n67037 & n67183) | (n67182 & n67183);
  assign n20923 = x141 & x176;
  assign n20924 = x140 & x177;
  assign n20925 = n20923 & n20924;
  assign n20926 = n20923 | n20924;
  assign n20927 = ~n20925 & n20926;
  assign n67192 = n20704 & n20927;
  assign n67193 = (n20927 & n67147) | (n20927 & n67192) | (n67147 & n67192);
  assign n67194 = n20704 | n20706;
  assign n67196 = n20927 & n67194;
  assign n67197 = (n67148 & n67192) | (n67148 & n67196) | (n67192 & n67196);
  assign n51354 = (n66988 & n67193) | (n66988 & n67197) | (n67193 & n67197);
  assign n67198 = n20704 | n20927;
  assign n67199 = n67147 | n67198;
  assign n67200 = n20927 | n67194;
  assign n67201 = (n67148 & n67198) | (n67148 & n67200) | (n67198 & n67200);
  assign n51357 = (n66988 & n67199) | (n66988 & n67201) | (n67199 & n67201);
  assign n20930 = ~n51354 & n51357;
  assign n20931 = x139 & x178;
  assign n20932 = n20930 & n20931;
  assign n20933 = n20930 | n20931;
  assign n20934 = ~n20932 & n20933;
  assign n67189 = n20711 | n20713;
  assign n67190 = (n20711 & n67153) | (n20711 & n67189) | (n67153 & n67189);
  assign n67202 = n20934 & n67190;
  assign n67191 = (n20711 & n67155) | (n20711 & n67189) | (n67155 & n67189);
  assign n67203 = n20934 & n67191;
  assign n67204 = (n67047 & n67202) | (n67047 & n67203) | (n67202 & n67203);
  assign n67205 = n20934 | n67190;
  assign n67206 = n20934 | n67191;
  assign n67207 = (n67047 & n67205) | (n67047 & n67206) | (n67205 & n67206);
  assign n20937 = ~n67204 & n67207;
  assign n20938 = x138 & x179;
  assign n20939 = n20937 & n20938;
  assign n20940 = n20937 | n20938;
  assign n20941 = ~n20939 & n20940;
  assign n67208 = n20718 | n20720;
  assign n67209 = (n20718 & n51247) | (n20718 & n67208) | (n51247 & n67208);
  assign n51358 = n20941 & n67209;
  assign n67210 = n20505 | n20718;
  assign n67211 = (n20718 & n20720) | (n20718 & n67210) | (n20720 & n67210);
  assign n51359 = n20941 & n67211;
  assign n51360 = (n67098 & n51358) | (n67098 & n51359) | (n51358 & n51359);
  assign n51361 = n20941 | n67209;
  assign n51362 = n20941 | n67211;
  assign n51363 = (n67098 & n51361) | (n67098 & n51362) | (n51361 & n51362);
  assign n20944 = ~n51360 & n51363;
  assign n20945 = x137 & x180;
  assign n20946 = n20944 & n20945;
  assign n20947 = n20944 | n20945;
  assign n20948 = ~n20946 & n20947;
  assign n67185 = n20725 | n20727;
  assign n67186 = (n20725 & n51245) | (n20725 & n67185) | (n51245 & n67185);
  assign n67212 = n20948 & n67186;
  assign n67187 = n20512 | n20725;
  assign n67188 = (n20725 & n20727) | (n20725 & n67187) | (n20727 & n67187);
  assign n67213 = n20948 & n67188;
  assign n67214 = (n67095 & n67212) | (n67095 & n67213) | (n67212 & n67213);
  assign n67215 = n20948 | n67186;
  assign n67216 = n20948 | n67188;
  assign n67217 = (n67095 & n67215) | (n67095 & n67216) | (n67215 & n67216);
  assign n20951 = ~n67214 & n67217;
  assign n20952 = x136 & x181;
  assign n20953 = n20951 & n20952;
  assign n20954 = n20951 | n20952;
  assign n20955 = ~n20953 & n20954;
  assign n51338 = n20732 | n20734;
  assign n51364 = n20955 & n51338;
  assign n51365 = n20732 & n20955;
  assign n51366 = (n51244 & n51364) | (n51244 & n51365) | (n51364 & n51365);
  assign n51367 = n20955 | n51338;
  assign n51368 = n20732 | n20955;
  assign n51369 = (n51244 & n51367) | (n51244 & n51368) | (n51367 & n51368);
  assign n20958 = ~n51366 & n51369;
  assign n20959 = x135 & x182;
  assign n20960 = n20958 & n20959;
  assign n20961 = n20958 | n20959;
  assign n20962 = ~n20960 & n20961;
  assign n51336 = n20739 | n20741;
  assign n51370 = n20962 & n51336;
  assign n51371 = n20739 & n20962;
  assign n51372 = (n67140 & n51370) | (n67140 & n51371) | (n51370 & n51371);
  assign n51373 = n20962 | n51336;
  assign n51374 = n20739 | n20962;
  assign n51375 = (n67140 & n51373) | (n67140 & n51374) | (n51373 & n51374);
  assign n20965 = ~n51372 & n51375;
  assign n20966 = x134 & x183;
  assign n20967 = n20965 & n20966;
  assign n20968 = n20965 | n20966;
  assign n20969 = ~n20967 & n20968;
  assign n51376 = n20746 & n20969;
  assign n67218 = (n20969 & n51280) | (n20969 & n51376) | (n51280 & n51376);
  assign n67219 = (n20969 & n51279) | (n20969 & n51376) | (n51279 & n51376);
  assign n67220 = (n67088 & n67218) | (n67088 & n67219) | (n67218 & n67219);
  assign n51378 = n20746 | n20969;
  assign n67221 = n51280 | n51378;
  assign n67222 = n51279 | n51378;
  assign n67223 = (n67088 & n67221) | (n67088 & n67222) | (n67221 & n67222);
  assign n20972 = ~n67220 & n67223;
  assign n20973 = x133 & x184;
  assign n20974 = n20972 & n20973;
  assign n20975 = n20972 | n20973;
  assign n20976 = ~n20974 & n20975;
  assign n20977 = n67184 & n20976;
  assign n20978 = n67184 | n20976;
  assign n20979 = ~n20977 & n20978;
  assign n20980 = x132 & x185;
  assign n20981 = n20979 & n20980;
  assign n20982 = n20979 | n20980;
  assign n20983 = ~n20981 & n20982;
  assign n51331 = n20760 | n20762;
  assign n51380 = n20983 & n51331;
  assign n51381 = n20760 & n20983;
  assign n51382 = (n67135 & n51380) | (n67135 & n51381) | (n51380 & n51381);
  assign n51383 = n20983 | n51331;
  assign n51384 = n20760 | n20983;
  assign n51385 = (n67135 & n51383) | (n67135 & n51384) | (n51383 & n51384);
  assign n20986 = ~n51382 & n51385;
  assign n20987 = x131 & x186;
  assign n20988 = n20986 & n20987;
  assign n20989 = n20986 | n20987;
  assign n20990 = ~n20988 & n20989;
  assign n51386 = n20767 & n20990;
  assign n51387 = (n20990 & n67164) | (n20990 & n51386) | (n67164 & n51386);
  assign n51388 = n20767 | n20990;
  assign n51389 = n67164 | n51388;
  assign n20993 = ~n51387 & n51389;
  assign n20994 = x130 & x187;
  assign n20995 = n20993 & n20994;
  assign n20996 = n20993 | n20994;
  assign n20997 = ~n20995 & n20996;
  assign n51390 = n20774 & n20997;
  assign n51391 = (n20997 & n51295) | (n20997 & n51390) | (n51295 & n51390);
  assign n51392 = n20774 | n20997;
  assign n51393 = n51295 | n51392;
  assign n21000 = ~n51391 & n51393;
  assign n21001 = x129 & x188;
  assign n21002 = n21000 & n21001;
  assign n21003 = n21000 | n21001;
  assign n21004 = ~n21002 & n21003;
  assign n51329 = n20781 | n20783;
  assign n51394 = n21004 & n51329;
  assign n51395 = n20781 & n21004;
  assign n51396 = (n51231 & n51394) | (n51231 & n51395) | (n51394 & n51395);
  assign n51397 = n21004 | n51329;
  assign n51398 = n20781 | n21004;
  assign n51399 = (n51231 & n51397) | (n51231 & n51398) | (n51397 & n51398);
  assign n21007 = ~n51396 & n51399;
  assign n21008 = x128 & x189;
  assign n21009 = n21007 & n21008;
  assign n21010 = n21007 | n21008;
  assign n21011 = ~n21009 & n21010;
  assign n51327 = n20788 | n20790;
  assign n67224 = n21011 & n51327;
  assign n67225 = n20788 & n21011;
  assign n67226 = (n51229 & n67224) | (n51229 & n67225) | (n67224 & n67225);
  assign n67227 = n21011 | n51327;
  assign n67228 = n20788 | n21011;
  assign n67229 = (n51229 & n67227) | (n51229 & n67228) | (n67227 & n67228);
  assign n21014 = ~n67226 & n67229;
  assign n21015 = x127 & x190;
  assign n21016 = n21014 & n21015;
  assign n21017 = n21014 | n21015;
  assign n21018 = ~n21016 & n21017;
  assign n51325 = n20795 | n20797;
  assign n67230 = n21018 & n51325;
  assign n67231 = n20795 & n21018;
  assign n67232 = (n51227 & n67230) | (n51227 & n67231) | (n67230 & n67231);
  assign n67233 = n21018 | n51325;
  assign n67234 = n20795 | n21018;
  assign n67235 = (n51227 & n67233) | (n51227 & n67234) | (n67233 & n67234);
  assign n21021 = ~n67232 & n67235;
  assign n21022 = x126 & x191;
  assign n21023 = n21021 & n21022;
  assign n21024 = n21021 | n21022;
  assign n21025 = ~n21023 & n21024;
  assign n21026 = n51324 & n21025;
  assign n21027 = n51324 | n21025;
  assign n21028 = ~n21026 & n21027;
  assign n21029 = x125 & x192;
  assign n21030 = n21028 & n21029;
  assign n21031 = n21028 | n21029;
  assign n21032 = ~n21030 & n21031;
  assign n21033 = n51322 & n21032;
  assign n21034 = n51322 | n21032;
  assign n21035 = ~n21033 & n21034;
  assign n21036 = x124 & x193;
  assign n21037 = n21035 & n21036;
  assign n21038 = n21035 | n21036;
  assign n21039 = ~n21037 & n21038;
  assign n21040 = n51320 & n21039;
  assign n21041 = n51320 | n21039;
  assign n21042 = ~n21040 & n21041;
  assign n21043 = x123 & x194;
  assign n21044 = n21042 & n21043;
  assign n21045 = n21042 | n21043;
  assign n21046 = ~n21044 & n21045;
  assign n21047 = n51318 & n21046;
  assign n21048 = n51318 | n21046;
  assign n21049 = ~n21047 & n21048;
  assign n21050 = x122 & x195;
  assign n21051 = n21049 & n21050;
  assign n21052 = n21049 | n21050;
  assign n21053 = ~n21051 & n21052;
  assign n21054 = n51316 & n21053;
  assign n21055 = n51316 | n21053;
  assign n21056 = ~n21054 & n21055;
  assign n21057 = x121 & x196;
  assign n21058 = n21056 & n21057;
  assign n21059 = n21056 | n21057;
  assign n21060 = ~n21058 & n21059;
  assign n21061 = n51314 & n21060;
  assign n21062 = n51314 | n21060;
  assign n21063 = ~n21061 & n21062;
  assign n21064 = x120 & x197;
  assign n21065 = n21063 & n21064;
  assign n21066 = n21063 | n21064;
  assign n21067 = ~n21065 & n21066;
  assign n21068 = n51312 & n21067;
  assign n21069 = n51312 | n21067;
  assign n21070 = ~n21068 & n21069;
  assign n21071 = x119 & x198;
  assign n21072 = n21070 & n21071;
  assign n21073 = n21070 | n21071;
  assign n21074 = ~n21072 & n21073;
  assign n21075 = n51310 & n21074;
  assign n21076 = n51310 | n21074;
  assign n21077 = ~n21075 & n21076;
  assign n21078 = x118 & x199;
  assign n21079 = n21077 & n21078;
  assign n21080 = n21077 | n21078;
  assign n21081 = ~n21079 & n21080;
  assign n21082 = n51308 & n21081;
  assign n21083 = n51308 | n21081;
  assign n21084 = ~n21082 & n21083;
  assign n21085 = x117 & x200;
  assign n21086 = n21084 & n21085;
  assign n21087 = n21084 | n21085;
  assign n21088 = ~n21086 & n21087;
  assign n21089 = n51306 & n21088;
  assign n21090 = n51306 | n21088;
  assign n21091 = ~n21089 & n21090;
  assign n21092 = x116 & x201;
  assign n21093 = n21091 & n21092;
  assign n21094 = n21091 | n21092;
  assign n21095 = ~n21093 & n21094;
  assign n21096 = n51304 & n21095;
  assign n21097 = n51304 | n21095;
  assign n21098 = ~n21096 & n21097;
  assign n21099 = x115 & x202;
  assign n21100 = n21098 & n21099;
  assign n21101 = n21098 | n21099;
  assign n21102 = ~n21100 & n21101;
  assign n21103 = n51302 & n21102;
  assign n21104 = n51302 | n21102;
  assign n21105 = ~n21103 & n21104;
  assign n21106 = x114 & x203;
  assign n21107 = n21105 & n21106;
  assign n21108 = n21105 | n21106;
  assign n21109 = ~n21107 & n21108;
  assign n21110 = n51300 & n21109;
  assign n21111 = n51300 | n21109;
  assign n21112 = ~n21110 & n21111;
  assign n21113 = x113 & x204;
  assign n21114 = n21112 & n21113;
  assign n21115 = n21112 | n21113;
  assign n21116 = ~n21114 & n21115;
  assign n21117 = n20893 & n21116;
  assign n21118 = n20893 | n21116;
  assign n21119 = ~n21117 & n21118;
  assign n21120 = x112 & x205;
  assign n21121 = n21119 & n21120;
  assign n21122 = n21119 | n21120;
  assign n21123 = ~n21121 & n21122;
  assign n67236 = n20893 | n21113;
  assign n67237 = (n20893 & n21112) | (n20893 & n67236) | (n21112 & n67236);
  assign n51401 = (n21114 & n21116) | (n21114 & n67237) | (n21116 & n67237);
  assign n67238 = n21107 | n51300;
  assign n67239 = (n21107 & n21109) | (n21107 & n67238) | (n21109 & n67238);
  assign n21126 = n21100 | n21103;
  assign n21127 = n21093 | n21096;
  assign n21128 = n21086 | n21089;
  assign n21129 = n21079 | n21082;
  assign n21130 = n21072 | n21075;
  assign n51402 = n21065 | n21067;
  assign n51403 = (n21065 & n51312) | (n21065 & n51402) | (n51312 & n51402);
  assign n51404 = n21058 | n21060;
  assign n51405 = (n21058 & n51314) | (n21058 & n51404) | (n51314 & n51404);
  assign n51406 = n21051 | n21053;
  assign n51407 = (n21051 & n51316) | (n21051 & n51406) | (n51316 & n51406);
  assign n51408 = n21044 | n21046;
  assign n51409 = (n21044 & n51318) | (n21044 & n51408) | (n51318 & n51408);
  assign n51410 = n21037 | n21039;
  assign n51411 = (n21037 & n51320) | (n21037 & n51410) | (n51320 & n51410);
  assign n51412 = n21030 | n21032;
  assign n51413 = (n21030 & n51322) | (n21030 & n51412) | (n51322 & n51412);
  assign n51326 = (n20795 & n51227) | (n20795 & n51325) | (n51227 & n51325);
  assign n51328 = (n20788 & n51229) | (n20788 & n51327) | (n51229 & n51327);
  assign n51426 = n20967 | n20969;
  assign n67242 = n20746 | n20967;
  assign n67243 = (n20967 & n20969) | (n20967 & n67242) | (n20969 & n67242);
  assign n67244 = (n51280 & n51426) | (n51280 & n67243) | (n51426 & n67243);
  assign n67245 = (n51279 & n51426) | (n51279 & n67243) | (n51426 & n67243);
  assign n67246 = (n67088 & n67244) | (n67088 & n67245) | (n67244 & n67245);
  assign n21152 = x142 & x176;
  assign n21153 = x141 & x177;
  assign n21154 = n21152 & n21153;
  assign n21155 = n21152 | n21153;
  assign n21156 = ~n21154 & n21155;
  assign n51436 = n20925 | n67197;
  assign n67254 = n21156 & n51436;
  assign n67251 = n20925 | n67192;
  assign n67252 = n20925 | n20927;
  assign n67253 = (n67147 & n67251) | (n67147 & n67252) | (n67251 & n67252);
  assign n67255 = n21156 & n67253;
  assign n67256 = (n66988 & n67254) | (n66988 & n67255) | (n67254 & n67255);
  assign n67257 = n21156 | n51436;
  assign n67258 = n21156 | n67253;
  assign n67259 = (n66988 & n67257) | (n66988 & n67258) | (n67257 & n67258);
  assign n21159 = ~n67256 & n67259;
  assign n21160 = x140 & x178;
  assign n21161 = n21159 & n21160;
  assign n21162 = n21159 | n21160;
  assign n21163 = ~n21161 & n21162;
  assign n51433 = n20932 | n20934;
  assign n51438 = n21163 & n51433;
  assign n51439 = n20932 & n21163;
  assign n67260 = (n51438 & n51439) | (n51438 & n67190) | (n51439 & n67190);
  assign n67261 = (n51438 & n51439) | (n51438 & n67191) | (n51439 & n67191);
  assign n67262 = (n67047 & n67260) | (n67047 & n67261) | (n67260 & n67261);
  assign n51441 = n21163 | n51433;
  assign n51442 = n20932 | n21163;
  assign n67263 = (n51441 & n51442) | (n51441 & n67190) | (n51442 & n67190);
  assign n67264 = (n51441 & n51442) | (n51441 & n67191) | (n51442 & n67191);
  assign n67265 = (n67047 & n67263) | (n67047 & n67264) | (n67263 & n67264);
  assign n21166 = ~n67262 & n67265;
  assign n21167 = x139 & x179;
  assign n21168 = n21166 & n21167;
  assign n21169 = n21166 | n21167;
  assign n21170 = ~n21168 & n21169;
  assign n51444 = n20939 & n21170;
  assign n67266 = (n21170 & n51358) | (n21170 & n51444) | (n51358 & n51444);
  assign n67267 = (n21170 & n51359) | (n21170 & n51444) | (n51359 & n51444);
  assign n67268 = (n67098 & n67266) | (n67098 & n67267) | (n67266 & n67267);
  assign n51446 = n20939 | n21170;
  assign n67269 = n51358 | n51446;
  assign n67270 = n51359 | n51446;
  assign n67271 = (n67098 & n67269) | (n67098 & n67270) | (n67269 & n67270);
  assign n21173 = ~n67268 & n67271;
  assign n21174 = x138 & x180;
  assign n21175 = n21173 & n21174;
  assign n21176 = n21173 | n21174;
  assign n21177 = ~n21175 & n21176;
  assign n51431 = n20946 | n20948;
  assign n51448 = n21177 & n51431;
  assign n51449 = n20946 & n21177;
  assign n67272 = (n51448 & n51449) | (n51448 & n67186) | (n51449 & n67186);
  assign n67273 = (n51448 & n51449) | (n51448 & n67188) | (n51449 & n67188);
  assign n67274 = (n67095 & n67272) | (n67095 & n67273) | (n67272 & n67273);
  assign n51451 = n21177 | n51431;
  assign n51452 = n20946 | n21177;
  assign n67275 = (n51451 & n51452) | (n51451 & n67186) | (n51452 & n67186);
  assign n67276 = (n51451 & n51452) | (n51451 & n67188) | (n51452 & n67188);
  assign n67277 = (n67095 & n67275) | (n67095 & n67276) | (n67275 & n67276);
  assign n21180 = ~n67274 & n67277;
  assign n21181 = x137 & x181;
  assign n21182 = n21180 & n21181;
  assign n21183 = n21180 | n21181;
  assign n21184 = ~n21182 & n21183;
  assign n67249 = n20953 | n20955;
  assign n67250 = (n20953 & n51338) | (n20953 & n67249) | (n51338 & n67249);
  assign n67278 = n21184 & n67250;
  assign n67247 = n20732 | n20953;
  assign n67248 = (n20953 & n20955) | (n20953 & n67247) | (n20955 & n67247);
  assign n67279 = n21184 & n67248;
  assign n67280 = (n51244 & n67278) | (n51244 & n67279) | (n67278 & n67279);
  assign n67281 = n21184 | n67250;
  assign n67282 = n21184 | n67248;
  assign n67283 = (n51244 & n67281) | (n51244 & n67282) | (n67281 & n67282);
  assign n21187 = ~n67280 & n67283;
  assign n21188 = x136 & x182;
  assign n21189 = n21187 & n21188;
  assign n21190 = n21187 | n21188;
  assign n21191 = ~n21189 & n21190;
  assign n51454 = n20960 & n21191;
  assign n51455 = (n21191 & n51372) | (n21191 & n51454) | (n51372 & n51454);
  assign n51456 = n20960 | n21191;
  assign n51457 = n51372 | n51456;
  assign n21194 = ~n51455 & n51457;
  assign n21195 = x135 & x183;
  assign n21196 = n21194 & n21195;
  assign n21197 = n21194 | n21195;
  assign n21198 = ~n21196 & n21197;
  assign n21199 = n67246 & n21198;
  assign n21200 = n67246 | n21198;
  assign n21201 = ~n21199 & n21200;
  assign n21202 = x134 & x184;
  assign n21203 = n21201 & n21202;
  assign n21204 = n21201 | n21202;
  assign n21205 = ~n21203 & n21204;
  assign n51423 = n20974 | n20976;
  assign n51458 = n21205 & n51423;
  assign n51459 = n20974 & n21205;
  assign n51460 = (n67184 & n51458) | (n67184 & n51459) | (n51458 & n51459);
  assign n51461 = n21205 | n51423;
  assign n51462 = n20974 | n21205;
  assign n51463 = (n67184 & n51461) | (n67184 & n51462) | (n51461 & n51462);
  assign n21208 = ~n51460 & n51463;
  assign n21209 = x133 & x185;
  assign n21210 = n21208 & n21209;
  assign n21211 = n21208 | n21209;
  assign n21212 = ~n21210 & n21211;
  assign n51464 = n20981 & n21212;
  assign n67284 = (n21212 & n51381) | (n21212 & n51464) | (n51381 & n51464);
  assign n67285 = (n21212 & n51380) | (n21212 & n51464) | (n51380 & n51464);
  assign n67286 = (n67135 & n67284) | (n67135 & n67285) | (n67284 & n67285);
  assign n51466 = n20981 | n21212;
  assign n67287 = n51381 | n51466;
  assign n67288 = n51380 | n51466;
  assign n67289 = (n67135 & n67287) | (n67135 & n67288) | (n67287 & n67288);
  assign n21215 = ~n67286 & n67289;
  assign n21216 = x132 & x186;
  assign n21217 = n21215 & n21216;
  assign n21218 = n21215 | n21216;
  assign n21219 = ~n21217 & n21218;
  assign n51421 = n20988 | n20990;
  assign n67290 = n21219 & n51421;
  assign n67240 = n20767 | n20988;
  assign n67241 = (n20988 & n20990) | (n20988 & n67240) | (n20990 & n67240);
  assign n67291 = n21219 & n67241;
  assign n67292 = (n67164 & n67290) | (n67164 & n67291) | (n67290 & n67291);
  assign n67293 = n21219 | n51421;
  assign n67294 = n21219 | n67241;
  assign n67295 = (n67164 & n67293) | (n67164 & n67294) | (n67293 & n67294);
  assign n21222 = ~n67292 & n67295;
  assign n21223 = x131 & x187;
  assign n21224 = n21222 & n21223;
  assign n21225 = n21222 | n21223;
  assign n21226 = ~n21224 & n21225;
  assign n51468 = n20995 & n21226;
  assign n67296 = (n21226 & n51390) | (n21226 & n51468) | (n51390 & n51468);
  assign n67297 = (n20997 & n21226) | (n20997 & n51468) | (n21226 & n51468);
  assign n67298 = (n51295 & n67296) | (n51295 & n67297) | (n67296 & n67297);
  assign n51470 = n20995 | n21226;
  assign n67299 = n51390 | n51470;
  assign n67300 = n20997 | n51470;
  assign n67301 = (n51295 & n67299) | (n51295 & n67300) | (n67299 & n67300);
  assign n21229 = ~n67298 & n67301;
  assign n21230 = x130 & x188;
  assign n21231 = n21229 & n21230;
  assign n21232 = n21229 | n21230;
  assign n21233 = ~n21231 & n21232;
  assign n51472 = n21002 & n21233;
  assign n51473 = (n21233 & n51396) | (n21233 & n51472) | (n51396 & n51472);
  assign n51474 = n21002 | n21233;
  assign n51475 = n51396 | n51474;
  assign n21236 = ~n51473 & n51475;
  assign n21237 = x129 & x189;
  assign n21238 = n21236 & n21237;
  assign n21239 = n21236 | n21237;
  assign n21240 = ~n21238 & n21239;
  assign n51418 = n21009 | n21011;
  assign n51476 = n21240 & n51418;
  assign n51477 = n21009 & n21240;
  assign n51478 = (n51328 & n51476) | (n51328 & n51477) | (n51476 & n51477);
  assign n51479 = n21240 | n51418;
  assign n51480 = n21009 | n21240;
  assign n51481 = (n51328 & n51479) | (n51328 & n51480) | (n51479 & n51480);
  assign n21243 = ~n51478 & n51481;
  assign n21244 = x128 & x190;
  assign n21245 = n21243 & n21244;
  assign n21246 = n21243 | n21244;
  assign n21247 = ~n21245 & n21246;
  assign n51416 = n21016 | n21018;
  assign n67302 = n21247 & n51416;
  assign n67303 = n21016 & n21247;
  assign n67304 = (n51326 & n67302) | (n51326 & n67303) | (n67302 & n67303);
  assign n67305 = n21247 | n51416;
  assign n67306 = n21016 | n21247;
  assign n67307 = (n51326 & n67305) | (n51326 & n67306) | (n67305 & n67306);
  assign n21250 = ~n67304 & n67307;
  assign n21251 = x127 & x191;
  assign n21252 = n21250 & n21251;
  assign n21253 = n21250 | n21251;
  assign n21254 = ~n21252 & n21253;
  assign n51414 = n21023 | n21025;
  assign n67308 = n21254 & n51414;
  assign n67309 = n21023 & n21254;
  assign n67310 = (n51324 & n67308) | (n51324 & n67309) | (n67308 & n67309);
  assign n67311 = n21254 | n51414;
  assign n67312 = n21023 | n21254;
  assign n67313 = (n51324 & n67311) | (n51324 & n67312) | (n67311 & n67312);
  assign n21257 = ~n67310 & n67313;
  assign n21258 = x126 & x192;
  assign n21259 = n21257 & n21258;
  assign n21260 = n21257 | n21258;
  assign n21261 = ~n21259 & n21260;
  assign n21262 = n51413 & n21261;
  assign n21263 = n51413 | n21261;
  assign n21264 = ~n21262 & n21263;
  assign n21265 = x125 & x193;
  assign n21266 = n21264 & n21265;
  assign n21267 = n21264 | n21265;
  assign n21268 = ~n21266 & n21267;
  assign n21269 = n51411 & n21268;
  assign n21270 = n51411 | n21268;
  assign n21271 = ~n21269 & n21270;
  assign n21272 = x124 & x194;
  assign n21273 = n21271 & n21272;
  assign n21274 = n21271 | n21272;
  assign n21275 = ~n21273 & n21274;
  assign n21276 = n51409 & n21275;
  assign n21277 = n51409 | n21275;
  assign n21278 = ~n21276 & n21277;
  assign n21279 = x123 & x195;
  assign n21280 = n21278 & n21279;
  assign n21281 = n21278 | n21279;
  assign n21282 = ~n21280 & n21281;
  assign n21283 = n51407 & n21282;
  assign n21284 = n51407 | n21282;
  assign n21285 = ~n21283 & n21284;
  assign n21286 = x122 & x196;
  assign n21287 = n21285 & n21286;
  assign n21288 = n21285 | n21286;
  assign n21289 = ~n21287 & n21288;
  assign n21290 = n51405 & n21289;
  assign n21291 = n51405 | n21289;
  assign n21292 = ~n21290 & n21291;
  assign n21293 = x121 & x197;
  assign n21294 = n21292 & n21293;
  assign n21295 = n21292 | n21293;
  assign n21296 = ~n21294 & n21295;
  assign n21297 = n51403 & n21296;
  assign n21298 = n51403 | n21296;
  assign n21299 = ~n21297 & n21298;
  assign n21300 = x120 & x198;
  assign n21301 = n21299 & n21300;
  assign n21302 = n21299 | n21300;
  assign n21303 = ~n21301 & n21302;
  assign n21304 = n21130 & n21303;
  assign n21305 = n21130 | n21303;
  assign n21306 = ~n21304 & n21305;
  assign n21307 = x119 & x199;
  assign n21308 = n21306 & n21307;
  assign n21309 = n21306 | n21307;
  assign n21310 = ~n21308 & n21309;
  assign n21311 = n21129 & n21310;
  assign n21312 = n21129 | n21310;
  assign n21313 = ~n21311 & n21312;
  assign n21314 = x118 & x200;
  assign n21315 = n21313 & n21314;
  assign n21316 = n21313 | n21314;
  assign n21317 = ~n21315 & n21316;
  assign n21318 = n21128 & n21317;
  assign n21319 = n21128 | n21317;
  assign n21320 = ~n21318 & n21319;
  assign n21321 = x117 & x201;
  assign n21322 = n21320 & n21321;
  assign n21323 = n21320 | n21321;
  assign n21324 = ~n21322 & n21323;
  assign n21325 = n21127 & n21324;
  assign n21326 = n21127 | n21324;
  assign n21327 = ~n21325 & n21326;
  assign n21328 = x116 & x202;
  assign n21329 = n21327 & n21328;
  assign n21330 = n21327 | n21328;
  assign n21331 = ~n21329 & n21330;
  assign n21332 = n21126 & n21331;
  assign n21333 = n21126 | n21331;
  assign n21334 = ~n21332 & n21333;
  assign n21335 = x115 & x203;
  assign n21336 = n21334 & n21335;
  assign n21337 = n21334 | n21335;
  assign n21338 = ~n21336 & n21337;
  assign n21339 = n67239 & n21338;
  assign n21340 = n67239 | n21338;
  assign n21341 = ~n21339 & n21340;
  assign n21342 = x114 & x204;
  assign n21343 = n21341 & n21342;
  assign n21344 = n21341 | n21342;
  assign n21345 = ~n21343 & n21344;
  assign n21346 = n51401 & n21345;
  assign n21347 = n51401 | n21345;
  assign n21348 = ~n21346 & n21347;
  assign n21349 = x113 & x205;
  assign n21350 = n21348 & n21349;
  assign n21351 = n21348 | n21349;
  assign n21352 = ~n21350 & n21351;
  assign n21353 = n21121 & n21352;
  assign n21354 = n21121 | n21352;
  assign n21355 = ~n21353 & n21354;
  assign n21356 = x112 & x206;
  assign n21357 = n21355 & n21356;
  assign n21358 = n21355 | n21356;
  assign n21359 = ~n21357 & n21358;
  assign n67314 = n21121 | n21349;
  assign n67315 = (n21121 & n21348) | (n21121 & n67314) | (n21348 & n67314);
  assign n51483 = (n21350 & n21352) | (n21350 & n67315) | (n21352 & n67315);
  assign n51484 = n21343 | n51401;
  assign n51485 = (n21343 & n21345) | (n21343 & n51484) | (n21345 & n51484);
  assign n67316 = n21336 | n67239;
  assign n67317 = (n21336 & n21338) | (n21336 & n67316) | (n21338 & n67316);
  assign n21363 = n21329 | n21332;
  assign n21364 = n21322 | n21325;
  assign n21365 = n21315 | n21318;
  assign n21366 = n21308 | n21311;
  assign n51486 = n21301 | n21303;
  assign n51487 = (n21130 & n21301) | (n21130 & n51486) | (n21301 & n51486);
  assign n51488 = n21294 | n21296;
  assign n51489 = (n21294 & n51403) | (n21294 & n51488) | (n51403 & n51488);
  assign n51490 = n21287 | n21289;
  assign n51491 = (n21287 & n51405) | (n21287 & n51490) | (n51405 & n51490);
  assign n51492 = n21280 | n21282;
  assign n51493 = (n21280 & n51407) | (n21280 & n51492) | (n51407 & n51492);
  assign n51494 = n21273 | n21275;
  assign n51495 = (n21273 & n51409) | (n21273 & n51494) | (n51409 & n51494);
  assign n51496 = n21266 | n21268;
  assign n51497 = (n21266 & n51411) | (n21266 & n51496) | (n51411 & n51496);
  assign n51415 = (n21023 & n51324) | (n21023 & n51414) | (n51324 & n51414);
  assign n51417 = (n21016 & n51326) | (n21016 & n51416) | (n51326 & n51416);
  assign n51507 = n21210 | n21212;
  assign n67318 = n20981 | n21210;
  assign n67319 = (n21210 & n21212) | (n21210 & n67318) | (n21212 & n67318);
  assign n67320 = (n51381 & n51507) | (n51381 & n67319) | (n51507 & n67319);
  assign n67321 = (n51380 & n51507) | (n51380 & n67319) | (n51507 & n67319);
  assign n67322 = (n67135 & n67320) | (n67135 & n67321) | (n67320 & n67321);
  assign n51342 = (n67095 & n67186) | (n67095 & n67188) | (n67186 & n67188);
  assign n21389 = x143 & x176;
  assign n21390 = x142 & x177;
  assign n21391 = n21389 & n21390;
  assign n21392 = n21389 | n21390;
  assign n21393 = ~n21391 & n21392;
  assign n51525 = n21154 | n21156;
  assign n51527 = n21393 & n51525;
  assign n51528 = n21154 & n21393;
  assign n67325 = (n51436 & n51527) | (n51436 & n51528) | (n51527 & n51528);
  assign n67326 = (n51527 & n51528) | (n51527 & n67253) | (n51528 & n67253);
  assign n67327 = (n66988 & n67325) | (n66988 & n67326) | (n67325 & n67326);
  assign n51530 = n21393 | n51525;
  assign n51531 = n21154 | n21393;
  assign n67328 = (n51436 & n51530) | (n51436 & n51531) | (n51530 & n51531);
  assign n67329 = (n51530 & n51531) | (n51530 & n67253) | (n51531 & n67253);
  assign n67330 = (n66988 & n67328) | (n66988 & n67329) | (n67328 & n67329);
  assign n21396 = ~n67327 & n67330;
  assign n21397 = x141 & x178;
  assign n21398 = n21396 & n21397;
  assign n21399 = n21396 | n21397;
  assign n21400 = ~n21398 & n21399;
  assign n67331 = n21161 | n21163;
  assign n67332 = (n21161 & n51433) | (n21161 & n67331) | (n51433 & n67331);
  assign n51533 = n21400 & n67332;
  assign n67333 = n20932 | n21161;
  assign n67334 = (n21161 & n21163) | (n21161 & n67333) | (n21163 & n67333);
  assign n51534 = n21400 & n67334;
  assign n67335 = (n51533 & n51534) | (n51533 & n67190) | (n51534 & n67190);
  assign n67336 = (n51533 & n51534) | (n51533 & n67191) | (n51534 & n67191);
  assign n67337 = (n67047 & n67335) | (n67047 & n67336) | (n67335 & n67336);
  assign n51536 = n21400 | n67332;
  assign n51537 = n21400 | n67334;
  assign n67338 = (n51536 & n51537) | (n51536 & n67190) | (n51537 & n67190);
  assign n67339 = (n51536 & n51537) | (n51536 & n67191) | (n51537 & n67191);
  assign n67340 = (n67047 & n67338) | (n67047 & n67339) | (n67338 & n67339);
  assign n21403 = ~n67337 & n67340;
  assign n21404 = x140 & x179;
  assign n21405 = n21403 & n21404;
  assign n21406 = n21403 | n21404;
  assign n21407 = ~n21405 & n21406;
  assign n67341 = n20939 | n21168;
  assign n67342 = (n21168 & n21170) | (n21168 & n67341) | (n21170 & n67341);
  assign n51539 = n21407 & n67342;
  assign n51520 = n21168 | n21170;
  assign n51540 = n21407 & n51520;
  assign n67343 = (n51358 & n51539) | (n51358 & n51540) | (n51539 & n51540);
  assign n67344 = (n51359 & n51539) | (n51359 & n51540) | (n51539 & n51540);
  assign n67345 = (n67098 & n67343) | (n67098 & n67344) | (n67343 & n67344);
  assign n51542 = n21407 | n67342;
  assign n51543 = n21407 | n51520;
  assign n67346 = (n51358 & n51542) | (n51358 & n51543) | (n51542 & n51543);
  assign n67347 = (n51359 & n51542) | (n51359 & n51543) | (n51542 & n51543);
  assign n67348 = (n67098 & n67346) | (n67098 & n67347) | (n67346 & n67347);
  assign n21410 = ~n67345 & n67348;
  assign n21411 = x139 & x180;
  assign n21412 = n21410 & n21411;
  assign n21413 = n21410 | n21411;
  assign n21414 = ~n21412 & n21413;
  assign n67349 = n21175 | n21177;
  assign n67350 = (n21175 & n51431) | (n21175 & n67349) | (n51431 & n67349);
  assign n51545 = n21414 & n67350;
  assign n67351 = n20946 | n21175;
  assign n67352 = (n21175 & n21177) | (n21175 & n67351) | (n21177 & n67351);
  assign n51546 = n21414 & n67352;
  assign n51547 = (n51342 & n51545) | (n51342 & n51546) | (n51545 & n51546);
  assign n51548 = n21414 | n67350;
  assign n51549 = n21414 | n67352;
  assign n51550 = (n51342 & n51548) | (n51342 & n51549) | (n51548 & n51549);
  assign n21417 = ~n51547 & n51550;
  assign n21418 = x138 & x181;
  assign n21419 = n21417 & n21418;
  assign n21420 = n21417 | n21418;
  assign n21421 = ~n21419 & n21420;
  assign n51514 = n21182 | n21184;
  assign n51551 = n21421 & n51514;
  assign n51552 = n21182 & n21421;
  assign n67353 = (n51551 & n51552) | (n51551 & n67250) | (n51552 & n67250);
  assign n67354 = (n51551 & n51552) | (n51551 & n67248) | (n51552 & n67248);
  assign n67355 = (n51244 & n67353) | (n51244 & n67354) | (n67353 & n67354);
  assign n51554 = n21421 | n51514;
  assign n51555 = n21182 | n21421;
  assign n67356 = (n51554 & n51555) | (n51554 & n67250) | (n51555 & n67250);
  assign n67357 = (n51554 & n51555) | (n51554 & n67248) | (n51555 & n67248);
  assign n67358 = (n51244 & n67356) | (n51244 & n67357) | (n67356 & n67357);
  assign n21424 = ~n67355 & n67358;
  assign n21425 = x137 & x182;
  assign n21426 = n21424 & n21425;
  assign n21427 = n21424 | n21425;
  assign n21428 = ~n21426 & n21427;
  assign n51512 = n21189 | n21191;
  assign n67359 = n21428 & n51512;
  assign n67323 = n20960 | n21189;
  assign n67324 = (n21189 & n21191) | (n21189 & n67323) | (n21191 & n67323);
  assign n67360 = n21428 & n67324;
  assign n67361 = (n51372 & n67359) | (n51372 & n67360) | (n67359 & n67360);
  assign n67362 = n21428 | n51512;
  assign n67363 = n21428 | n67324;
  assign n67364 = (n51372 & n67362) | (n51372 & n67363) | (n67362 & n67363);
  assign n21431 = ~n67361 & n67364;
  assign n21432 = x136 & x183;
  assign n21433 = n21431 & n21432;
  assign n21434 = n21431 | n21432;
  assign n21435 = ~n21433 & n21434;
  assign n51509 = n21196 | n21198;
  assign n51557 = n21435 & n51509;
  assign n51558 = n21196 & n21435;
  assign n51559 = (n67246 & n51557) | (n67246 & n51558) | (n51557 & n51558);
  assign n51560 = n21435 | n51509;
  assign n51561 = n21196 | n21435;
  assign n51562 = (n67246 & n51560) | (n67246 & n51561) | (n51560 & n51561);
  assign n21438 = ~n51559 & n51562;
  assign n21439 = x135 & x184;
  assign n21440 = n21438 & n21439;
  assign n21441 = n21438 | n21439;
  assign n21442 = ~n21440 & n21441;
  assign n51563 = n21203 & n21442;
  assign n67365 = (n21442 & n51459) | (n21442 & n51563) | (n51459 & n51563);
  assign n67366 = (n21442 & n51458) | (n21442 & n51563) | (n51458 & n51563);
  assign n67367 = (n67184 & n67365) | (n67184 & n67366) | (n67365 & n67366);
  assign n51565 = n21203 | n21442;
  assign n67368 = n51459 | n51565;
  assign n67369 = n51458 | n51565;
  assign n67370 = (n67184 & n67368) | (n67184 & n67369) | (n67368 & n67369);
  assign n21445 = ~n67367 & n67370;
  assign n21446 = x134 & x185;
  assign n21447 = n21445 & n21446;
  assign n21448 = n21445 | n21446;
  assign n21449 = ~n21447 & n21448;
  assign n21450 = n67322 & n21449;
  assign n21451 = n67322 | n21449;
  assign n21452 = ~n21450 & n21451;
  assign n21453 = x133 & x186;
  assign n21454 = n21452 & n21453;
  assign n21455 = n21452 | n21453;
  assign n21456 = ~n21454 & n21455;
  assign n51504 = n21217 | n21219;
  assign n51567 = n21456 & n51504;
  assign n51568 = n21217 & n21456;
  assign n67371 = (n51421 & n51567) | (n51421 & n51568) | (n51567 & n51568);
  assign n67372 = (n51567 & n51568) | (n51567 & n67241) | (n51568 & n67241);
  assign n67373 = (n67164 & n67371) | (n67164 & n67372) | (n67371 & n67372);
  assign n51570 = n21456 | n51504;
  assign n51571 = n21217 | n21456;
  assign n67374 = (n51421 & n51570) | (n51421 & n51571) | (n51570 & n51571);
  assign n67375 = (n51570 & n51571) | (n51570 & n67241) | (n51571 & n67241);
  assign n67376 = (n67164 & n67374) | (n67164 & n67375) | (n67374 & n67375);
  assign n21459 = ~n67373 & n67376;
  assign n21460 = x132 & x187;
  assign n21461 = n21459 & n21460;
  assign n21462 = n21459 | n21460;
  assign n21463 = ~n21461 & n21462;
  assign n51573 = n21224 & n21463;
  assign n51574 = (n21463 & n67298) | (n21463 & n51573) | (n67298 & n51573);
  assign n51575 = n21224 | n21463;
  assign n51576 = n67298 | n51575;
  assign n21466 = ~n51574 & n51576;
  assign n21467 = x131 & x188;
  assign n21468 = n21466 & n21467;
  assign n21469 = n21466 | n21467;
  assign n21470 = ~n21468 & n21469;
  assign n51577 = n21231 & n21470;
  assign n51578 = (n21470 & n51473) | (n21470 & n51577) | (n51473 & n51577);
  assign n51579 = n21231 | n21470;
  assign n51580 = n51473 | n51579;
  assign n21473 = ~n51578 & n51580;
  assign n21474 = x130 & x189;
  assign n21475 = n21473 & n21474;
  assign n21476 = n21473 | n21474;
  assign n21477 = ~n21475 & n21476;
  assign n51581 = n21238 & n21477;
  assign n51582 = (n21477 & n51478) | (n21477 & n51581) | (n51478 & n51581);
  assign n51583 = n21238 | n21477;
  assign n51584 = n51478 | n51583;
  assign n21480 = ~n51582 & n51584;
  assign n21481 = x129 & x190;
  assign n21482 = n21480 & n21481;
  assign n21483 = n21480 | n21481;
  assign n21484 = ~n21482 & n21483;
  assign n51502 = n21245 | n21247;
  assign n51585 = n21484 & n51502;
  assign n51586 = n21245 & n21484;
  assign n51587 = (n51417 & n51585) | (n51417 & n51586) | (n51585 & n51586);
  assign n51588 = n21484 | n51502;
  assign n51589 = n21245 | n21484;
  assign n51590 = (n51417 & n51588) | (n51417 & n51589) | (n51588 & n51589);
  assign n21487 = ~n51587 & n51590;
  assign n21488 = x128 & x191;
  assign n21489 = n21487 & n21488;
  assign n21490 = n21487 | n21488;
  assign n21491 = ~n21489 & n21490;
  assign n51500 = n21252 | n21254;
  assign n67377 = n21491 & n51500;
  assign n67378 = n21252 & n21491;
  assign n67379 = (n51415 & n67377) | (n51415 & n67378) | (n67377 & n67378);
  assign n67380 = n21491 | n51500;
  assign n67381 = n21252 | n21491;
  assign n67382 = (n51415 & n67380) | (n51415 & n67381) | (n67380 & n67381);
  assign n21494 = ~n67379 & n67382;
  assign n21495 = x127 & x192;
  assign n21496 = n21494 & n21495;
  assign n21497 = n21494 | n21495;
  assign n21498 = ~n21496 & n21497;
  assign n51498 = n21259 | n21261;
  assign n67383 = n21498 & n51498;
  assign n67384 = n21259 & n21498;
  assign n67385 = (n51413 & n67383) | (n51413 & n67384) | (n67383 & n67384);
  assign n67386 = n21498 | n51498;
  assign n67387 = n21259 | n21498;
  assign n67388 = (n51413 & n67386) | (n51413 & n67387) | (n67386 & n67387);
  assign n21501 = ~n67385 & n67388;
  assign n21502 = x126 & x193;
  assign n21503 = n21501 & n21502;
  assign n21504 = n21501 | n21502;
  assign n21505 = ~n21503 & n21504;
  assign n21506 = n51497 & n21505;
  assign n21507 = n51497 | n21505;
  assign n21508 = ~n21506 & n21507;
  assign n21509 = x125 & x194;
  assign n21510 = n21508 & n21509;
  assign n21511 = n21508 | n21509;
  assign n21512 = ~n21510 & n21511;
  assign n21513 = n51495 & n21512;
  assign n21514 = n51495 | n21512;
  assign n21515 = ~n21513 & n21514;
  assign n21516 = x124 & x195;
  assign n21517 = n21515 & n21516;
  assign n21518 = n21515 | n21516;
  assign n21519 = ~n21517 & n21518;
  assign n21520 = n51493 & n21519;
  assign n21521 = n51493 | n21519;
  assign n21522 = ~n21520 & n21521;
  assign n21523 = x123 & x196;
  assign n21524 = n21522 & n21523;
  assign n21525 = n21522 | n21523;
  assign n21526 = ~n21524 & n21525;
  assign n21527 = n51491 & n21526;
  assign n21528 = n51491 | n21526;
  assign n21529 = ~n21527 & n21528;
  assign n21530 = x122 & x197;
  assign n21531 = n21529 & n21530;
  assign n21532 = n21529 | n21530;
  assign n21533 = ~n21531 & n21532;
  assign n21534 = n51489 & n21533;
  assign n21535 = n51489 | n21533;
  assign n21536 = ~n21534 & n21535;
  assign n21537 = x121 & x198;
  assign n21538 = n21536 & n21537;
  assign n21539 = n21536 | n21537;
  assign n21540 = ~n21538 & n21539;
  assign n21541 = n51487 & n21540;
  assign n21542 = n51487 | n21540;
  assign n21543 = ~n21541 & n21542;
  assign n21544 = x120 & x199;
  assign n21545 = n21543 & n21544;
  assign n21546 = n21543 | n21544;
  assign n21547 = ~n21545 & n21546;
  assign n21548 = n21366 & n21547;
  assign n21549 = n21366 | n21547;
  assign n21550 = ~n21548 & n21549;
  assign n21551 = x119 & x200;
  assign n21552 = n21550 & n21551;
  assign n21553 = n21550 | n21551;
  assign n21554 = ~n21552 & n21553;
  assign n21555 = n21365 & n21554;
  assign n21556 = n21365 | n21554;
  assign n21557 = ~n21555 & n21556;
  assign n21558 = x118 & x201;
  assign n21559 = n21557 & n21558;
  assign n21560 = n21557 | n21558;
  assign n21561 = ~n21559 & n21560;
  assign n21562 = n21364 & n21561;
  assign n21563 = n21364 | n21561;
  assign n21564 = ~n21562 & n21563;
  assign n21565 = x117 & x202;
  assign n21566 = n21564 & n21565;
  assign n21567 = n21564 | n21565;
  assign n21568 = ~n21566 & n21567;
  assign n21569 = n21363 & n21568;
  assign n21570 = n21363 | n21568;
  assign n21571 = ~n21569 & n21570;
  assign n21572 = x116 & x203;
  assign n21573 = n21571 & n21572;
  assign n21574 = n21571 | n21572;
  assign n21575 = ~n21573 & n21574;
  assign n21576 = n67317 & n21575;
  assign n21577 = n67317 | n21575;
  assign n21578 = ~n21576 & n21577;
  assign n21579 = x115 & x204;
  assign n21580 = n21578 & n21579;
  assign n21581 = n21578 | n21579;
  assign n21582 = ~n21580 & n21581;
  assign n21583 = n51485 & n21582;
  assign n21584 = n51485 | n21582;
  assign n21585 = ~n21583 & n21584;
  assign n21586 = x114 & x205;
  assign n21587 = n21585 & n21586;
  assign n21588 = n21585 | n21586;
  assign n21589 = ~n21587 & n21588;
  assign n21590 = n51483 & n21589;
  assign n21591 = n51483 | n21589;
  assign n21592 = ~n21590 & n21591;
  assign n21593 = x113 & x206;
  assign n21594 = n21592 & n21593;
  assign n21595 = n21592 | n21593;
  assign n21596 = ~n21594 & n21595;
  assign n21597 = n21357 & n21596;
  assign n21598 = n21357 | n21596;
  assign n21599 = ~n21597 & n21598;
  assign n21600 = x112 & x207;
  assign n21601 = n21599 & n21600;
  assign n21602 = n21599 | n21600;
  assign n21603 = ~n21601 & n21602;
  assign n67389 = n21357 | n21593;
  assign n67390 = (n21357 & n21592) | (n21357 & n67389) | (n21592 & n67389);
  assign n51592 = (n21594 & n21596) | (n21594 & n67390) | (n21596 & n67390);
  assign n51593 = n21587 | n51483;
  assign n51594 = (n21587 & n21589) | (n21587 & n51593) | (n21589 & n51593);
  assign n51595 = n21580 | n51485;
  assign n51596 = (n21580 & n21582) | (n21580 & n51595) | (n21582 & n51595);
  assign n67391 = n21573 | n67317;
  assign n67392 = (n21573 & n21575) | (n21573 & n67391) | (n21575 & n67391);
  assign n21608 = n21566 | n21569;
  assign n21609 = n21559 | n21562;
  assign n21610 = n21552 | n21555;
  assign n51597 = n21545 | n21547;
  assign n51598 = (n21366 & n21545) | (n21366 & n51597) | (n21545 & n51597);
  assign n51599 = n21538 | n21540;
  assign n51600 = (n21538 & n51487) | (n21538 & n51599) | (n51487 & n51599);
  assign n51601 = n21531 | n21533;
  assign n51602 = (n21531 & n51489) | (n21531 & n51601) | (n51489 & n51601);
  assign n51603 = n21524 | n21526;
  assign n51604 = (n21524 & n51491) | (n21524 & n51603) | (n51491 & n51603);
  assign n51605 = n21517 | n21519;
  assign n51606 = (n21517 & n51493) | (n21517 & n51605) | (n51493 & n51605);
  assign n51607 = n21510 | n21512;
  assign n51608 = (n21510 & n51495) | (n21510 & n51607) | (n51495 & n51607);
  assign n51499 = (n21259 & n51413) | (n21259 & n51498) | (n51413 & n51498);
  assign n51501 = (n21252 & n51415) | (n21252 & n51500) | (n51415 & n51500);
  assign n51621 = n21440 | n21442;
  assign n67395 = n21203 | n21440;
  assign n67396 = (n21440 & n21442) | (n21440 & n67395) | (n21442 & n67395);
  assign n67397 = (n51459 & n51621) | (n51459 & n67396) | (n51621 & n67396);
  assign n67398 = (n51458 & n51621) | (n51458 & n67396) | (n51621 & n67396);
  assign n67399 = (n67184 & n67397) | (n67184 & n67398) | (n67397 & n67398);
  assign n51430 = (n51244 & n67248) | (n51244 & n67250) | (n67248 & n67250);
  assign n67402 = n21405 | n21407;
  assign n67403 = (n21405 & n67342) | (n21405 & n67402) | (n67342 & n67402);
  assign n67404 = (n21405 & n51520) | (n21405 & n67402) | (n51520 & n67402);
  assign n67405 = (n51358 & n67403) | (n51358 & n67404) | (n67403 & n67404);
  assign n67406 = (n51359 & n67403) | (n51359 & n67404) | (n67403 & n67404);
  assign n67407 = (n67098 & n67405) | (n67098 & n67406) | (n67405 & n67406);
  assign n21634 = x144 & x176;
  assign n21635 = x143 & x177;
  assign n21636 = n21634 & n21635;
  assign n21637 = n21634 | n21635;
  assign n21638 = ~n21636 & n21637;
  assign n67408 = n21391 | n21393;
  assign n67409 = (n21391 & n51525) | (n21391 & n67408) | (n51525 & n67408);
  assign n51637 = n21638 & n67409;
  assign n67410 = n21154 | n21391;
  assign n67411 = (n21391 & n21393) | (n21391 & n67410) | (n21393 & n67410);
  assign n51638 = n21638 & n67411;
  assign n67412 = (n51436 & n51637) | (n51436 & n51638) | (n51637 & n51638);
  assign n67413 = (n51637 & n51638) | (n51637 & n67253) | (n51638 & n67253);
  assign n67414 = (n66988 & n67412) | (n66988 & n67413) | (n67412 & n67413);
  assign n51640 = n21638 | n67409;
  assign n51641 = n21638 | n67411;
  assign n67415 = (n51436 & n51640) | (n51436 & n51641) | (n51640 & n51641);
  assign n67416 = (n51640 & n51641) | (n51640 & n67253) | (n51641 & n67253);
  assign n67417 = (n66988 & n67415) | (n66988 & n67416) | (n67415 & n67416);
  assign n21641 = ~n67414 & n67417;
  assign n21642 = x142 & x178;
  assign n21643 = n21641 & n21642;
  assign n21644 = n21641 | n21642;
  assign n21645 = ~n21643 & n21644;
  assign n67418 = n21398 | n21400;
  assign n67423 = (n21398 & n67334) | (n21398 & n67418) | (n67334 & n67418);
  assign n51644 = n21645 & n67423;
  assign n67420 = n21645 & n67418;
  assign n67421 = n21398 & n21645;
  assign n67422 = (n67332 & n67420) | (n67332 & n67421) | (n67420 & n67421);
  assign n67424 = (n51644 & n67190) | (n51644 & n67422) | (n67190 & n67422);
  assign n67425 = (n51644 & n67191) | (n51644 & n67422) | (n67191 & n67422);
  assign n67426 = (n67047 & n67424) | (n67047 & n67425) | (n67424 & n67425);
  assign n51647 = n21645 | n67423;
  assign n67427 = n21645 | n67418;
  assign n67428 = n21398 | n21645;
  assign n67429 = (n67332 & n67427) | (n67332 & n67428) | (n67427 & n67428);
  assign n67430 = (n51647 & n67190) | (n51647 & n67429) | (n67190 & n67429);
  assign n67431 = (n51647 & n67191) | (n51647 & n67429) | (n67191 & n67429);
  assign n67432 = (n67047 & n67430) | (n67047 & n67431) | (n67430 & n67431);
  assign n21648 = ~n67426 & n67432;
  assign n21649 = x141 & x179;
  assign n21650 = n21648 & n21649;
  assign n21651 = n21648 | n21649;
  assign n21652 = ~n21650 & n21651;
  assign n21653 = n67407 & n21652;
  assign n21654 = n67407 | n21652;
  assign n21655 = ~n21653 & n21654;
  assign n21656 = x140 & x180;
  assign n21657 = n21655 & n21656;
  assign n21658 = n21655 | n21656;
  assign n21659 = ~n21657 & n21658;
  assign n51649 = n21412 & n21659;
  assign n67433 = (n21659 & n51545) | (n21659 & n51649) | (n51545 & n51649);
  assign n67434 = (n21659 & n51546) | (n21659 & n51649) | (n51546 & n51649);
  assign n67435 = (n51342 & n67433) | (n51342 & n67434) | (n67433 & n67434);
  assign n51651 = n21412 | n21659;
  assign n67436 = n51545 | n51651;
  assign n67437 = n51546 | n51651;
  assign n67438 = (n51342 & n67436) | (n51342 & n67437) | (n67436 & n67437);
  assign n21662 = ~n67435 & n67438;
  assign n21663 = x139 & x181;
  assign n21664 = n21662 & n21663;
  assign n21665 = n21662 | n21663;
  assign n21666 = ~n21664 & n21665;
  assign n51625 = n21419 | n51551;
  assign n67439 = n21666 & n51625;
  assign n67400 = n21182 | n21419;
  assign n67401 = (n21419 & n21421) | (n21419 & n67400) | (n21421 & n67400);
  assign n67440 = n21666 & n67401;
  assign n67441 = (n51430 & n67439) | (n51430 & n67440) | (n67439 & n67440);
  assign n67442 = n21666 | n51625;
  assign n67443 = n21666 | n67401;
  assign n67444 = (n51430 & n67442) | (n51430 & n67443) | (n67442 & n67443);
  assign n21669 = ~n67441 & n67444;
  assign n21670 = x138 & x182;
  assign n21671 = n21669 & n21670;
  assign n21672 = n21669 | n21670;
  assign n21673 = ~n21671 & n21672;
  assign n51623 = n21426 | n21428;
  assign n51653 = n21673 & n51623;
  assign n51654 = n21426 & n21673;
  assign n67445 = (n51512 & n51653) | (n51512 & n51654) | (n51653 & n51654);
  assign n67446 = (n51653 & n51654) | (n51653 & n67324) | (n51654 & n67324);
  assign n67447 = (n51372 & n67445) | (n51372 & n67446) | (n67445 & n67446);
  assign n51656 = n21673 | n51623;
  assign n51657 = n21426 | n21673;
  assign n67448 = (n51512 & n51656) | (n51512 & n51657) | (n51656 & n51657);
  assign n67449 = (n51656 & n51657) | (n51656 & n67324) | (n51657 & n67324);
  assign n67450 = (n51372 & n67448) | (n51372 & n67449) | (n67448 & n67449);
  assign n21676 = ~n67447 & n67450;
  assign n21677 = x137 & x183;
  assign n21678 = n21676 & n21677;
  assign n21679 = n21676 | n21677;
  assign n21680 = ~n21678 & n21679;
  assign n51659 = n21433 & n21680;
  assign n51660 = (n21680 & n51559) | (n21680 & n51659) | (n51559 & n51659);
  assign n51661 = n21433 | n21680;
  assign n51662 = n51559 | n51661;
  assign n21683 = ~n51660 & n51662;
  assign n21684 = x136 & x184;
  assign n21685 = n21683 & n21684;
  assign n21686 = n21683 | n21684;
  assign n21687 = ~n21685 & n21686;
  assign n21688 = n67399 & n21687;
  assign n21689 = n67399 | n21687;
  assign n21690 = ~n21688 & n21689;
  assign n21691 = x135 & x185;
  assign n21692 = n21690 & n21691;
  assign n21693 = n21690 | n21691;
  assign n21694 = ~n21692 & n21693;
  assign n51618 = n21447 | n21449;
  assign n51663 = n21694 & n51618;
  assign n51664 = n21447 & n21694;
  assign n51665 = (n67322 & n51663) | (n67322 & n51664) | (n51663 & n51664);
  assign n51666 = n21694 | n51618;
  assign n51667 = n21447 | n21694;
  assign n51668 = (n67322 & n51666) | (n67322 & n51667) | (n51666 & n51667);
  assign n21697 = ~n51665 & n51668;
  assign n21698 = x134 & x186;
  assign n21699 = n21697 & n21698;
  assign n21700 = n21697 | n21698;
  assign n21701 = ~n21699 & n21700;
  assign n51669 = n21454 & n21701;
  assign n51670 = (n21701 & n67373) | (n21701 & n51669) | (n67373 & n51669);
  assign n51671 = n21454 | n21701;
  assign n51672 = n67373 | n51671;
  assign n21704 = ~n51670 & n51672;
  assign n21705 = x133 & x187;
  assign n21706 = n21704 & n21705;
  assign n21707 = n21704 | n21705;
  assign n21708 = ~n21706 & n21707;
  assign n51616 = n21461 | n21463;
  assign n67451 = n21708 & n51616;
  assign n67393 = n21224 | n21461;
  assign n67394 = (n21461 & n21463) | (n21461 & n67393) | (n21463 & n67393);
  assign n67452 = n21708 & n67394;
  assign n67453 = (n67298 & n67451) | (n67298 & n67452) | (n67451 & n67452);
  assign n67454 = n21708 | n51616;
  assign n67455 = n21708 | n67394;
  assign n67456 = (n67298 & n67454) | (n67298 & n67455) | (n67454 & n67455);
  assign n21711 = ~n67453 & n67456;
  assign n21712 = x132 & x188;
  assign n21713 = n21711 & n21712;
  assign n21714 = n21711 | n21712;
  assign n21715 = ~n21713 & n21714;
  assign n51673 = n21468 & n21715;
  assign n67457 = (n21715 & n51577) | (n21715 & n51673) | (n51577 & n51673);
  assign n67458 = (n21470 & n21715) | (n21470 & n51673) | (n21715 & n51673);
  assign n67459 = (n51473 & n67457) | (n51473 & n67458) | (n67457 & n67458);
  assign n51675 = n21468 | n21715;
  assign n67460 = n51577 | n51675;
  assign n67461 = n21470 | n51675;
  assign n67462 = (n51473 & n67460) | (n51473 & n67461) | (n67460 & n67461);
  assign n21718 = ~n67459 & n67462;
  assign n21719 = x131 & x189;
  assign n21720 = n21718 & n21719;
  assign n21721 = n21718 | n21719;
  assign n21722 = ~n21720 & n21721;
  assign n51677 = n21475 & n21722;
  assign n51678 = (n21722 & n51582) | (n21722 & n51677) | (n51582 & n51677);
  assign n51679 = n21475 | n21722;
  assign n51680 = n51582 | n51679;
  assign n21725 = ~n51678 & n51680;
  assign n21726 = x130 & x190;
  assign n21727 = n21725 & n21726;
  assign n21728 = n21725 | n21726;
  assign n21729 = ~n21727 & n21728;
  assign n51681 = n21482 & n21729;
  assign n51682 = (n21729 & n51587) | (n21729 & n51681) | (n51587 & n51681);
  assign n51683 = n21482 | n21729;
  assign n51684 = n51587 | n51683;
  assign n21732 = ~n51682 & n51684;
  assign n21733 = x129 & x191;
  assign n21734 = n21732 & n21733;
  assign n21735 = n21732 | n21733;
  assign n21736 = ~n21734 & n21735;
  assign n51613 = n21489 | n21491;
  assign n51685 = n21736 & n51613;
  assign n51686 = n21489 & n21736;
  assign n51687 = (n51501 & n51685) | (n51501 & n51686) | (n51685 & n51686);
  assign n51688 = n21736 | n51613;
  assign n51689 = n21489 | n21736;
  assign n51690 = (n51501 & n51688) | (n51501 & n51689) | (n51688 & n51689);
  assign n21739 = ~n51687 & n51690;
  assign n21740 = x128 & x192;
  assign n21741 = n21739 & n21740;
  assign n21742 = n21739 | n21740;
  assign n21743 = ~n21741 & n21742;
  assign n51611 = n21496 | n21498;
  assign n67463 = n21743 & n51611;
  assign n67464 = n21496 & n21743;
  assign n67465 = (n51499 & n67463) | (n51499 & n67464) | (n67463 & n67464);
  assign n67466 = n21743 | n51611;
  assign n67467 = n21496 | n21743;
  assign n67468 = (n51499 & n67466) | (n51499 & n67467) | (n67466 & n67467);
  assign n21746 = ~n67465 & n67468;
  assign n21747 = x127 & x193;
  assign n21748 = n21746 & n21747;
  assign n21749 = n21746 | n21747;
  assign n21750 = ~n21748 & n21749;
  assign n51609 = n21503 | n21505;
  assign n67469 = n21750 & n51609;
  assign n67470 = n21503 & n21750;
  assign n67471 = (n51497 & n67469) | (n51497 & n67470) | (n67469 & n67470);
  assign n67472 = n21750 | n51609;
  assign n67473 = n21503 | n21750;
  assign n67474 = (n51497 & n67472) | (n51497 & n67473) | (n67472 & n67473);
  assign n21753 = ~n67471 & n67474;
  assign n21754 = x126 & x194;
  assign n21755 = n21753 & n21754;
  assign n21756 = n21753 | n21754;
  assign n21757 = ~n21755 & n21756;
  assign n21758 = n51608 & n21757;
  assign n21759 = n51608 | n21757;
  assign n21760 = ~n21758 & n21759;
  assign n21761 = x125 & x195;
  assign n21762 = n21760 & n21761;
  assign n21763 = n21760 | n21761;
  assign n21764 = ~n21762 & n21763;
  assign n21765 = n51606 & n21764;
  assign n21766 = n51606 | n21764;
  assign n21767 = ~n21765 & n21766;
  assign n21768 = x124 & x196;
  assign n21769 = n21767 & n21768;
  assign n21770 = n21767 | n21768;
  assign n21771 = ~n21769 & n21770;
  assign n21772 = n51604 & n21771;
  assign n21773 = n51604 | n21771;
  assign n21774 = ~n21772 & n21773;
  assign n21775 = x123 & x197;
  assign n21776 = n21774 & n21775;
  assign n21777 = n21774 | n21775;
  assign n21778 = ~n21776 & n21777;
  assign n21779 = n51602 & n21778;
  assign n21780 = n51602 | n21778;
  assign n21781 = ~n21779 & n21780;
  assign n21782 = x122 & x198;
  assign n21783 = n21781 & n21782;
  assign n21784 = n21781 | n21782;
  assign n21785 = ~n21783 & n21784;
  assign n21786 = n51600 & n21785;
  assign n21787 = n51600 | n21785;
  assign n21788 = ~n21786 & n21787;
  assign n21789 = x121 & x199;
  assign n21790 = n21788 & n21789;
  assign n21791 = n21788 | n21789;
  assign n21792 = ~n21790 & n21791;
  assign n21793 = n51598 & n21792;
  assign n21794 = n51598 | n21792;
  assign n21795 = ~n21793 & n21794;
  assign n21796 = x120 & x200;
  assign n21797 = n21795 & n21796;
  assign n21798 = n21795 | n21796;
  assign n21799 = ~n21797 & n21798;
  assign n21800 = n21610 & n21799;
  assign n21801 = n21610 | n21799;
  assign n21802 = ~n21800 & n21801;
  assign n21803 = x119 & x201;
  assign n21804 = n21802 & n21803;
  assign n21805 = n21802 | n21803;
  assign n21806 = ~n21804 & n21805;
  assign n21807 = n21609 & n21806;
  assign n21808 = n21609 | n21806;
  assign n21809 = ~n21807 & n21808;
  assign n21810 = x118 & x202;
  assign n21811 = n21809 & n21810;
  assign n21812 = n21809 | n21810;
  assign n21813 = ~n21811 & n21812;
  assign n21814 = n21608 & n21813;
  assign n21815 = n21608 | n21813;
  assign n21816 = ~n21814 & n21815;
  assign n21817 = x117 & x203;
  assign n21818 = n21816 & n21817;
  assign n21819 = n21816 | n21817;
  assign n21820 = ~n21818 & n21819;
  assign n21821 = n67392 & n21820;
  assign n21822 = n67392 | n21820;
  assign n21823 = ~n21821 & n21822;
  assign n21824 = x116 & x204;
  assign n21825 = n21823 & n21824;
  assign n21826 = n21823 | n21824;
  assign n21827 = ~n21825 & n21826;
  assign n21828 = n51596 & n21827;
  assign n21829 = n51596 | n21827;
  assign n21830 = ~n21828 & n21829;
  assign n21831 = x115 & x205;
  assign n21832 = n21830 & n21831;
  assign n21833 = n21830 | n21831;
  assign n21834 = ~n21832 & n21833;
  assign n21835 = n51594 & n21834;
  assign n21836 = n51594 | n21834;
  assign n21837 = ~n21835 & n21836;
  assign n21838 = x114 & x206;
  assign n21839 = n21837 & n21838;
  assign n21840 = n21837 | n21838;
  assign n21841 = ~n21839 & n21840;
  assign n21842 = n51592 & n21841;
  assign n21843 = n51592 | n21841;
  assign n21844 = ~n21842 & n21843;
  assign n21845 = x113 & x207;
  assign n21846 = n21844 & n21845;
  assign n21847 = n21844 | n21845;
  assign n21848 = ~n21846 & n21847;
  assign n21849 = n21601 & n21848;
  assign n21850 = n21601 | n21848;
  assign n21851 = ~n21849 & n21850;
  assign n21852 = x112 & x208;
  assign n21853 = n21851 & n21852;
  assign n21854 = n21851 | n21852;
  assign n21855 = ~n21853 & n21854;
  assign n67475 = n21601 | n21845;
  assign n67476 = (n21601 & n21844) | (n21601 & n67475) | (n21844 & n67475);
  assign n51692 = (n21846 & n21848) | (n21846 & n67476) | (n21848 & n67476);
  assign n51693 = n21839 | n51592;
  assign n51694 = (n21839 & n21841) | (n21839 & n51693) | (n21841 & n51693);
  assign n51695 = n21832 | n51594;
  assign n51696 = (n21832 & n21834) | (n21832 & n51695) | (n21834 & n51695);
  assign n51697 = n21825 | n51596;
  assign n51698 = (n21825 & n21827) | (n21825 & n51697) | (n21827 & n51697);
  assign n67477 = n21818 | n67392;
  assign n67478 = (n21818 & n21820) | (n21818 & n67477) | (n21820 & n67477);
  assign n21861 = n21811 | n21814;
  assign n21862 = n21804 | n21807;
  assign n51699 = n21797 | n21799;
  assign n51700 = (n21610 & n21797) | (n21610 & n51699) | (n21797 & n51699);
  assign n51701 = n21790 | n21792;
  assign n51702 = (n21790 & n51598) | (n21790 & n51701) | (n51598 & n51701);
  assign n51703 = n21783 | n21785;
  assign n51704 = (n21783 & n51600) | (n21783 & n51703) | (n51600 & n51703);
  assign n51705 = n21776 | n21778;
  assign n51706 = (n21776 & n51602) | (n21776 & n51705) | (n51602 & n51705);
  assign n51707 = n21769 | n21771;
  assign n51708 = (n21769 & n51604) | (n21769 & n51707) | (n51604 & n51707);
  assign n51709 = n21762 | n21764;
  assign n51710 = (n21762 & n51606) | (n21762 & n51709) | (n51606 & n51709);
  assign n51610 = (n21503 & n51497) | (n21503 & n51609) | (n51497 & n51609);
  assign n51612 = (n21496 & n51499) | (n21496 & n51611) | (n51499 & n51611);
  assign n51617 = (n67298 & n67394) | (n67298 & n51616) | (n67394 & n51616);
  assign n51513 = (n51372 & n67324) | (n51372 & n51512) | (n67324 & n51512);
  assign n21887 = x145 & x176;
  assign n21888 = x144 & x177;
  assign n21889 = n21887 & n21888;
  assign n21890 = n21887 | n21888;
  assign n21891 = ~n21889 & n21890;
  assign n67485 = n21636 | n21638;
  assign n67490 = (n21636 & n67411) | (n21636 & n67485) | (n67411 & n67485);
  assign n51741 = n21891 & n67490;
  assign n67487 = n21891 & n67485;
  assign n67488 = n21636 & n21891;
  assign n67489 = (n67409 & n67487) | (n67409 & n67488) | (n67487 & n67488);
  assign n67491 = (n51436 & n51741) | (n51436 & n67489) | (n51741 & n67489);
  assign n67492 = (n51741 & n67253) | (n51741 & n67489) | (n67253 & n67489);
  assign n67493 = (n66988 & n67491) | (n66988 & n67492) | (n67491 & n67492);
  assign n51744 = n21891 | n67490;
  assign n67494 = n21891 | n67485;
  assign n67495 = n21636 | n21891;
  assign n67496 = (n67409 & n67494) | (n67409 & n67495) | (n67494 & n67495);
  assign n67497 = (n51436 & n51744) | (n51436 & n67496) | (n51744 & n67496);
  assign n67498 = (n51744 & n67253) | (n51744 & n67496) | (n67253 & n67496);
  assign n67499 = (n66988 & n67497) | (n66988 & n67498) | (n67497 & n67498);
  assign n21894 = ~n67493 & n67499;
  assign n21895 = x143 & x178;
  assign n21896 = n21894 & n21895;
  assign n21897 = n21894 | n21895;
  assign n21898 = ~n21896 & n21897;
  assign n51746 = n21643 & n21898;
  assign n51747 = (n21898 & n67426) | (n21898 & n51746) | (n67426 & n51746);
  assign n51748 = n21643 | n21898;
  assign n51749 = n67426 | n51748;
  assign n21901 = ~n51747 & n51749;
  assign n21902 = x142 & x179;
  assign n21903 = n21901 & n21902;
  assign n21904 = n21901 | n21902;
  assign n21905 = ~n21903 & n21904;
  assign n51735 = n21650 | n21652;
  assign n51750 = n21905 & n51735;
  assign n51751 = n21650 & n21905;
  assign n51752 = (n67407 & n51750) | (n67407 & n51751) | (n51750 & n51751);
  assign n51753 = n21905 | n51735;
  assign n51754 = n21650 | n21905;
  assign n51755 = (n67407 & n51753) | (n67407 & n51754) | (n51753 & n51754);
  assign n21908 = ~n51752 & n51755;
  assign n21909 = x141 & x180;
  assign n21910 = n21908 & n21909;
  assign n21911 = n21908 | n21909;
  assign n21912 = ~n21910 & n21911;
  assign n67500 = n21412 | n21657;
  assign n67501 = (n21657 & n21659) | (n21657 & n67500) | (n21659 & n67500);
  assign n51756 = n21912 & n67501;
  assign n51733 = n21657 | n21659;
  assign n51757 = n21912 & n51733;
  assign n67502 = (n51545 & n51756) | (n51545 & n51757) | (n51756 & n51757);
  assign n67503 = (n51546 & n51756) | (n51546 & n51757) | (n51756 & n51757);
  assign n67504 = (n51342 & n67502) | (n51342 & n67503) | (n67502 & n67503);
  assign n51759 = n21912 | n67501;
  assign n51760 = n21912 | n51733;
  assign n67505 = (n51545 & n51759) | (n51545 & n51760) | (n51759 & n51760);
  assign n67506 = (n51546 & n51759) | (n51546 & n51760) | (n51759 & n51760);
  assign n67507 = (n51342 & n67505) | (n51342 & n67506) | (n67505 & n67506);
  assign n21915 = ~n67504 & n67507;
  assign n21916 = x140 & x181;
  assign n21917 = n21915 & n21916;
  assign n21918 = n21915 | n21916;
  assign n21919 = ~n21917 & n21918;
  assign n51730 = n21664 | n21666;
  assign n51762 = n21919 & n51730;
  assign n51763 = n21664 & n21919;
  assign n67508 = (n51625 & n51762) | (n51625 & n51763) | (n51762 & n51763);
  assign n67509 = (n51762 & n51763) | (n51762 & n67401) | (n51763 & n67401);
  assign n67510 = (n51430 & n67508) | (n51430 & n67509) | (n67508 & n67509);
  assign n51765 = n21919 | n51730;
  assign n51766 = n21664 | n21919;
  assign n67511 = (n51625 & n51765) | (n51625 & n51766) | (n51765 & n51766);
  assign n67512 = (n51765 & n51766) | (n51765 & n67401) | (n51766 & n67401);
  assign n67513 = (n51430 & n67511) | (n51430 & n67512) | (n67511 & n67512);
  assign n21922 = ~n67510 & n67513;
  assign n21923 = x139 & x182;
  assign n21924 = n21922 & n21923;
  assign n21925 = n21922 | n21923;
  assign n21926 = ~n21924 & n21925;
  assign n51728 = n21671 | n51653;
  assign n67514 = n21926 & n51728;
  assign n67483 = n21426 | n21671;
  assign n67484 = (n21671 & n21673) | (n21671 & n67483) | (n21673 & n67483);
  assign n67515 = n21926 & n67484;
  assign n67516 = (n51513 & n67514) | (n51513 & n67515) | (n67514 & n67515);
  assign n67517 = n21926 | n51728;
  assign n67518 = n21926 | n67484;
  assign n67519 = (n51513 & n67517) | (n51513 & n67518) | (n67517 & n67518);
  assign n21929 = ~n67516 & n67519;
  assign n21930 = x138 & x183;
  assign n21931 = n21929 & n21930;
  assign n21932 = n21929 | n21930;
  assign n21933 = ~n21931 & n21932;
  assign n51725 = n21678 | n21680;
  assign n67520 = n21933 & n51725;
  assign n67481 = n21433 | n21678;
  assign n67482 = (n21678 & n21680) | (n21678 & n67481) | (n21680 & n67481);
  assign n67521 = n21933 & n67482;
  assign n67522 = (n51559 & n67520) | (n51559 & n67521) | (n67520 & n67521);
  assign n67523 = n21933 | n51725;
  assign n67524 = n21933 | n67482;
  assign n67525 = (n51559 & n67523) | (n51559 & n67524) | (n67523 & n67524);
  assign n21936 = ~n67522 & n67525;
  assign n21937 = x137 & x184;
  assign n21938 = n21936 & n21937;
  assign n21939 = n21936 | n21937;
  assign n21940 = ~n21938 & n21939;
  assign n51722 = n21685 | n21687;
  assign n51768 = n21940 & n51722;
  assign n51769 = n21685 & n21940;
  assign n51770 = (n67399 & n51768) | (n67399 & n51769) | (n51768 & n51769);
  assign n51771 = n21940 | n51722;
  assign n51772 = n21685 | n21940;
  assign n51773 = (n67399 & n51771) | (n67399 & n51772) | (n51771 & n51772);
  assign n21943 = ~n51770 & n51773;
  assign n21944 = x136 & x185;
  assign n21945 = n21943 & n21944;
  assign n21946 = n21943 | n21944;
  assign n21947 = ~n21945 & n21946;
  assign n51774 = n21692 & n21947;
  assign n67526 = (n21947 & n51664) | (n21947 & n51774) | (n51664 & n51774);
  assign n67527 = (n21947 & n51663) | (n21947 & n51774) | (n51663 & n51774);
  assign n67528 = (n67322 & n67526) | (n67322 & n67527) | (n67526 & n67527);
  assign n51776 = n21692 | n21947;
  assign n67529 = n51664 | n51776;
  assign n67530 = n51663 | n51776;
  assign n67531 = (n67322 & n67529) | (n67322 & n67530) | (n67529 & n67530);
  assign n21950 = ~n67528 & n67531;
  assign n21951 = x135 & x186;
  assign n21952 = n21950 & n21951;
  assign n21953 = n21950 | n21951;
  assign n21954 = ~n21952 & n21953;
  assign n51720 = n21699 | n21701;
  assign n67532 = n21954 & n51720;
  assign n67479 = n21454 | n21699;
  assign n67480 = (n21699 & n21701) | (n21699 & n67479) | (n21701 & n67479);
  assign n67533 = n21954 & n67480;
  assign n67534 = (n67373 & n67532) | (n67373 & n67533) | (n67532 & n67533);
  assign n67535 = n21954 | n51720;
  assign n67536 = n21954 | n67480;
  assign n67537 = (n67373 & n67535) | (n67373 & n67536) | (n67535 & n67536);
  assign n21957 = ~n67534 & n67537;
  assign n21958 = x134 & x187;
  assign n21959 = n21957 & n21958;
  assign n21960 = n21957 | n21958;
  assign n21961 = ~n21959 & n21960;
  assign n51717 = n21706 | n21708;
  assign n51778 = n21961 & n51717;
  assign n51779 = n21706 & n21961;
  assign n51780 = (n51617 & n51778) | (n51617 & n51779) | (n51778 & n51779);
  assign n51781 = n21961 | n51717;
  assign n51782 = n21706 | n21961;
  assign n51783 = (n51617 & n51781) | (n51617 & n51782) | (n51781 & n51782);
  assign n21964 = ~n51780 & n51783;
  assign n21965 = x133 & x188;
  assign n21966 = n21964 & n21965;
  assign n21967 = n21964 | n21965;
  assign n21968 = ~n21966 & n21967;
  assign n51784 = n21713 & n21968;
  assign n51785 = (n21968 & n67459) | (n21968 & n51784) | (n67459 & n51784);
  assign n51786 = n21713 | n21968;
  assign n51787 = n67459 | n51786;
  assign n21971 = ~n51785 & n51787;
  assign n21972 = x132 & x189;
  assign n21973 = n21971 & n21972;
  assign n21974 = n21971 | n21972;
  assign n21975 = ~n21973 & n21974;
  assign n51788 = n21720 & n21975;
  assign n51789 = (n21975 & n51678) | (n21975 & n51788) | (n51678 & n51788);
  assign n51790 = n21720 | n21975;
  assign n51791 = n51678 | n51790;
  assign n21978 = ~n51789 & n51791;
  assign n21979 = x131 & x190;
  assign n21980 = n21978 & n21979;
  assign n21981 = n21978 | n21979;
  assign n21982 = ~n21980 & n21981;
  assign n51792 = n21727 & n21982;
  assign n51793 = (n21982 & n51682) | (n21982 & n51792) | (n51682 & n51792);
  assign n51794 = n21727 | n21982;
  assign n51795 = n51682 | n51794;
  assign n21985 = ~n51793 & n51795;
  assign n21986 = x130 & x191;
  assign n21987 = n21985 & n21986;
  assign n21988 = n21985 | n21986;
  assign n21989 = ~n21987 & n21988;
  assign n51796 = n21734 & n21989;
  assign n51797 = (n21989 & n51687) | (n21989 & n51796) | (n51687 & n51796);
  assign n51798 = n21734 | n21989;
  assign n51799 = n51687 | n51798;
  assign n21992 = ~n51797 & n51799;
  assign n21993 = x129 & x192;
  assign n21994 = n21992 & n21993;
  assign n21995 = n21992 | n21993;
  assign n21996 = ~n21994 & n21995;
  assign n51715 = n21741 | n21743;
  assign n51800 = n21996 & n51715;
  assign n51801 = n21741 & n21996;
  assign n51802 = (n51612 & n51800) | (n51612 & n51801) | (n51800 & n51801);
  assign n51803 = n21996 | n51715;
  assign n51804 = n21741 | n21996;
  assign n51805 = (n51612 & n51803) | (n51612 & n51804) | (n51803 & n51804);
  assign n21999 = ~n51802 & n51805;
  assign n22000 = x128 & x193;
  assign n22001 = n21999 & n22000;
  assign n22002 = n21999 | n22000;
  assign n22003 = ~n22001 & n22002;
  assign n51713 = n21748 | n21750;
  assign n67538 = n22003 & n51713;
  assign n67539 = n21748 & n22003;
  assign n67540 = (n51610 & n67538) | (n51610 & n67539) | (n67538 & n67539);
  assign n67541 = n22003 | n51713;
  assign n67542 = n21748 | n22003;
  assign n67543 = (n51610 & n67541) | (n51610 & n67542) | (n67541 & n67542);
  assign n22006 = ~n67540 & n67543;
  assign n22007 = x127 & x194;
  assign n22008 = n22006 & n22007;
  assign n22009 = n22006 | n22007;
  assign n22010 = ~n22008 & n22009;
  assign n51711 = n21755 | n21757;
  assign n67544 = n22010 & n51711;
  assign n67545 = n21755 & n22010;
  assign n67546 = (n51608 & n67544) | (n51608 & n67545) | (n67544 & n67545);
  assign n67547 = n22010 | n51711;
  assign n67548 = n21755 | n22010;
  assign n67549 = (n51608 & n67547) | (n51608 & n67548) | (n67547 & n67548);
  assign n22013 = ~n67546 & n67549;
  assign n22014 = x126 & x195;
  assign n22015 = n22013 & n22014;
  assign n22016 = n22013 | n22014;
  assign n22017 = ~n22015 & n22016;
  assign n22018 = n51710 & n22017;
  assign n22019 = n51710 | n22017;
  assign n22020 = ~n22018 & n22019;
  assign n22021 = x125 & x196;
  assign n22022 = n22020 & n22021;
  assign n22023 = n22020 | n22021;
  assign n22024 = ~n22022 & n22023;
  assign n22025 = n51708 & n22024;
  assign n22026 = n51708 | n22024;
  assign n22027 = ~n22025 & n22026;
  assign n22028 = x124 & x197;
  assign n22029 = n22027 & n22028;
  assign n22030 = n22027 | n22028;
  assign n22031 = ~n22029 & n22030;
  assign n22032 = n51706 & n22031;
  assign n22033 = n51706 | n22031;
  assign n22034 = ~n22032 & n22033;
  assign n22035 = x123 & x198;
  assign n22036 = n22034 & n22035;
  assign n22037 = n22034 | n22035;
  assign n22038 = ~n22036 & n22037;
  assign n22039 = n51704 & n22038;
  assign n22040 = n51704 | n22038;
  assign n22041 = ~n22039 & n22040;
  assign n22042 = x122 & x199;
  assign n22043 = n22041 & n22042;
  assign n22044 = n22041 | n22042;
  assign n22045 = ~n22043 & n22044;
  assign n22046 = n51702 & n22045;
  assign n22047 = n51702 | n22045;
  assign n22048 = ~n22046 & n22047;
  assign n22049 = x121 & x200;
  assign n22050 = n22048 & n22049;
  assign n22051 = n22048 | n22049;
  assign n22052 = ~n22050 & n22051;
  assign n22053 = n51700 & n22052;
  assign n22054 = n51700 | n22052;
  assign n22055 = ~n22053 & n22054;
  assign n22056 = x120 & x201;
  assign n22057 = n22055 & n22056;
  assign n22058 = n22055 | n22056;
  assign n22059 = ~n22057 & n22058;
  assign n22060 = n21862 & n22059;
  assign n22061 = n21862 | n22059;
  assign n22062 = ~n22060 & n22061;
  assign n22063 = x119 & x202;
  assign n22064 = n22062 & n22063;
  assign n22065 = n22062 | n22063;
  assign n22066 = ~n22064 & n22065;
  assign n22067 = n21861 & n22066;
  assign n22068 = n21861 | n22066;
  assign n22069 = ~n22067 & n22068;
  assign n22070 = x118 & x203;
  assign n22071 = n22069 & n22070;
  assign n22072 = n22069 | n22070;
  assign n22073 = ~n22071 & n22072;
  assign n22074 = n67478 & n22073;
  assign n22075 = n67478 | n22073;
  assign n22076 = ~n22074 & n22075;
  assign n22077 = x117 & x204;
  assign n22078 = n22076 & n22077;
  assign n22079 = n22076 | n22077;
  assign n22080 = ~n22078 & n22079;
  assign n22081 = n51698 & n22080;
  assign n22082 = n51698 | n22080;
  assign n22083 = ~n22081 & n22082;
  assign n22084 = x116 & x205;
  assign n22085 = n22083 & n22084;
  assign n22086 = n22083 | n22084;
  assign n22087 = ~n22085 & n22086;
  assign n22088 = n51696 & n22087;
  assign n22089 = n51696 | n22087;
  assign n22090 = ~n22088 & n22089;
  assign n22091 = x115 & x206;
  assign n22092 = n22090 & n22091;
  assign n22093 = n22090 | n22091;
  assign n22094 = ~n22092 & n22093;
  assign n22095 = n51694 & n22094;
  assign n22096 = n51694 | n22094;
  assign n22097 = ~n22095 & n22096;
  assign n22098 = x114 & x207;
  assign n22099 = n22097 & n22098;
  assign n22100 = n22097 | n22098;
  assign n22101 = ~n22099 & n22100;
  assign n22102 = n51692 & n22101;
  assign n22103 = n51692 | n22101;
  assign n22104 = ~n22102 & n22103;
  assign n22105 = x113 & x208;
  assign n22106 = n22104 & n22105;
  assign n22107 = n22104 | n22105;
  assign n22108 = ~n22106 & n22107;
  assign n22109 = n21853 & n22108;
  assign n22110 = n21853 | n22108;
  assign n22111 = ~n22109 & n22110;
  assign n22112 = x112 & x209;
  assign n22113 = n22111 & n22112;
  assign n22114 = n22111 | n22112;
  assign n22115 = ~n22113 & n22114;
  assign n67550 = n21853 | n22105;
  assign n67551 = (n21853 & n22104) | (n21853 & n67550) | (n22104 & n67550);
  assign n51807 = (n22106 & n22108) | (n22106 & n67551) | (n22108 & n67551);
  assign n51808 = n22099 | n51692;
  assign n51809 = (n22099 & n22101) | (n22099 & n51808) | (n22101 & n51808);
  assign n51810 = n22092 | n51694;
  assign n51811 = (n22092 & n22094) | (n22092 & n51810) | (n22094 & n51810);
  assign n51812 = n22085 | n51696;
  assign n51813 = (n22085 & n22087) | (n22085 & n51812) | (n22087 & n51812);
  assign n51814 = n22078 | n51698;
  assign n51815 = (n22078 & n22080) | (n22078 & n51814) | (n22080 & n51814);
  assign n67552 = n22071 | n67478;
  assign n67553 = (n22071 & n22073) | (n22071 & n67552) | (n22073 & n67552);
  assign n22122 = n22064 | n22067;
  assign n51816 = n22057 | n22059;
  assign n51817 = (n21862 & n22057) | (n21862 & n51816) | (n22057 & n51816);
  assign n51818 = n22050 | n22052;
  assign n51819 = (n22050 & n51700) | (n22050 & n51818) | (n51700 & n51818);
  assign n51820 = n22043 | n22045;
  assign n51821 = (n22043 & n51702) | (n22043 & n51820) | (n51702 & n51820);
  assign n51822 = n22036 | n22038;
  assign n51823 = (n22036 & n51704) | (n22036 & n51822) | (n51704 & n51822);
  assign n51824 = n22029 | n22031;
  assign n51825 = (n22029 & n51706) | (n22029 & n51824) | (n51706 & n51824);
  assign n51826 = n22022 | n22024;
  assign n51827 = (n22022 & n51708) | (n22022 & n51826) | (n51708 & n51826);
  assign n51712 = (n21755 & n51608) | (n21755 & n51711) | (n51608 & n51711);
  assign n51714 = (n21748 & n51610) | (n21748 & n51713) | (n51610 & n51713);
  assign n51840 = n21945 | n21947;
  assign n67556 = n21692 | n21945;
  assign n67557 = (n21945 & n21947) | (n21945 & n67556) | (n21947 & n67556);
  assign n67558 = (n51664 & n51840) | (n51664 & n67557) | (n51840 & n67557);
  assign n67559 = (n51663 & n51840) | (n51663 & n67557) | (n51840 & n67557);
  assign n67560 = (n67322 & n67558) | (n67322 & n67559) | (n67558 & n67559);
  assign n51726 = (n51559 & n67482) | (n51559 & n51725) | (n67482 & n51725);
  assign n67561 = n21917 | n21919;
  assign n67562 = (n21917 & n51730) | (n21917 & n67561) | (n51730 & n67561);
  assign n67563 = n21664 | n21917;
  assign n67564 = (n21917 & n21919) | (n21917 & n67563) | (n21919 & n67563);
  assign n67565 = (n51625 & n67562) | (n51625 & n67564) | (n67562 & n67564);
  assign n67566 = (n67401 & n67562) | (n67401 & n67564) | (n67562 & n67564);
  assign n67567 = (n51430 & n67565) | (n51430 & n67566) | (n67565 & n67566);
  assign n22148 = x146 & x176;
  assign n22149 = x145 & x177;
  assign n22150 = n22148 & n22149;
  assign n22151 = n22148 | n22149;
  assign n22152 = ~n22150 & n22151;
  assign n67568 = n21889 & n22152;
  assign n67569 = (n22152 & n67489) | (n22152 & n67568) | (n67489 & n67568);
  assign n67570 = n21889 | n21891;
  assign n67572 = n22152 & n67570;
  assign n67573 = (n67490 & n67568) | (n67490 & n67572) | (n67568 & n67572);
  assign n67574 = (n51436 & n67569) | (n51436 & n67573) | (n67569 & n67573);
  assign n67575 = (n67253 & n67569) | (n67253 & n67573) | (n67569 & n67573);
  assign n67576 = (n66988 & n67574) | (n66988 & n67575) | (n67574 & n67575);
  assign n67577 = n21889 | n22152;
  assign n67578 = n67489 | n67577;
  assign n67579 = n22152 | n67570;
  assign n67580 = (n67490 & n67577) | (n67490 & n67579) | (n67577 & n67579);
  assign n67581 = (n51436 & n67578) | (n51436 & n67580) | (n67578 & n67580);
  assign n67582 = (n67253 & n67578) | (n67253 & n67580) | (n67578 & n67580);
  assign n67583 = (n66988 & n67581) | (n66988 & n67582) | (n67581 & n67582);
  assign n22155 = ~n67576 & n67583;
  assign n22156 = x144 & x178;
  assign n22157 = n22155 & n22156;
  assign n22158 = n22155 | n22156;
  assign n22159 = ~n22157 & n22158;
  assign n67584 = n21643 | n21896;
  assign n67585 = (n21896 & n21898) | (n21896 & n67584) | (n21898 & n67584);
  assign n51864 = n22159 & n67585;
  assign n51853 = n21896 | n21898;
  assign n51865 = n22159 & n51853;
  assign n51866 = (n67426 & n51864) | (n67426 & n51865) | (n51864 & n51865);
  assign n51867 = n22159 | n67585;
  assign n51868 = n22159 | n51853;
  assign n51869 = (n67426 & n51867) | (n67426 & n51868) | (n51867 & n51868);
  assign n22162 = ~n51866 & n51869;
  assign n22163 = x143 & x179;
  assign n22164 = n22162 & n22163;
  assign n22165 = n22162 | n22163;
  assign n22166 = ~n22164 & n22165;
  assign n67586 = n21903 & n22166;
  assign n67587 = (n22166 & n51750) | (n22166 & n67586) | (n51750 & n67586);
  assign n67588 = n21650 | n21903;
  assign n67589 = (n21903 & n21905) | (n21903 & n67588) | (n21905 & n67588);
  assign n51871 = n22166 & n67589;
  assign n51872 = (n67407 & n67587) | (n67407 & n51871) | (n67587 & n51871);
  assign n67590 = n21903 | n22166;
  assign n67591 = n51750 | n67590;
  assign n51874 = n22166 | n67589;
  assign n51875 = (n67407 & n67591) | (n67407 & n51874) | (n67591 & n51874);
  assign n22169 = ~n51872 & n51875;
  assign n22170 = x142 & x180;
  assign n22171 = n22169 & n22170;
  assign n22172 = n22169 | n22170;
  assign n22173 = ~n22171 & n22172;
  assign n51876 = n21910 & n22173;
  assign n51877 = (n22173 & n67504) | (n22173 & n51876) | (n67504 & n51876);
  assign n51878 = n21910 | n22173;
  assign n51879 = n67504 | n51878;
  assign n22176 = ~n51877 & n51879;
  assign n22177 = x141 & x181;
  assign n22178 = n22176 & n22177;
  assign n22179 = n22176 | n22177;
  assign n22180 = ~n22178 & n22179;
  assign n22181 = n67567 & n22180;
  assign n22182 = n67567 | n22180;
  assign n22183 = ~n22181 & n22182;
  assign n22184 = x140 & x182;
  assign n22185 = n22183 & n22184;
  assign n22186 = n22183 | n22184;
  assign n22187 = ~n22185 & n22186;
  assign n51844 = n21924 | n21926;
  assign n51880 = n22187 & n51844;
  assign n51881 = n21924 & n22187;
  assign n67592 = (n51728 & n51880) | (n51728 & n51881) | (n51880 & n51881);
  assign n67593 = (n51880 & n51881) | (n51880 & n67484) | (n51881 & n67484);
  assign n67594 = (n51513 & n67592) | (n51513 & n67593) | (n67592 & n67593);
  assign n51883 = n22187 | n51844;
  assign n51884 = n21924 | n22187;
  assign n67595 = (n51728 & n51883) | (n51728 & n51884) | (n51883 & n51884);
  assign n67596 = (n51883 & n51884) | (n51883 & n67484) | (n51884 & n67484);
  assign n67597 = (n51513 & n67595) | (n51513 & n67596) | (n67595 & n67596);
  assign n22190 = ~n67594 & n67597;
  assign n22191 = x139 & x183;
  assign n22192 = n22190 & n22191;
  assign n22193 = n22190 | n22191;
  assign n22194 = ~n22192 & n22193;
  assign n51842 = n21931 | n21933;
  assign n51886 = n22194 & n51842;
  assign n51887 = n21931 & n22194;
  assign n51888 = (n51726 & n51886) | (n51726 & n51887) | (n51886 & n51887);
  assign n51889 = n22194 | n51842;
  assign n51890 = n21931 | n22194;
  assign n51891 = (n51726 & n51889) | (n51726 & n51890) | (n51889 & n51890);
  assign n22197 = ~n51888 & n51891;
  assign n22198 = x138 & x184;
  assign n22199 = n22197 & n22198;
  assign n22200 = n22197 | n22198;
  assign n22201 = ~n22199 & n22200;
  assign n51892 = n21938 & n22201;
  assign n51893 = (n22201 & n51770) | (n22201 & n51892) | (n51770 & n51892);
  assign n51894 = n21938 | n22201;
  assign n51895 = n51770 | n51894;
  assign n22204 = ~n51893 & n51895;
  assign n22205 = x137 & x185;
  assign n22206 = n22204 & n22205;
  assign n22207 = n22204 | n22205;
  assign n22208 = ~n22206 & n22207;
  assign n22209 = n67560 & n22208;
  assign n22210 = n67560 | n22208;
  assign n22211 = ~n22209 & n22210;
  assign n22212 = x136 & x186;
  assign n22213 = n22211 & n22212;
  assign n22214 = n22211 | n22212;
  assign n22215 = ~n22213 & n22214;
  assign n51837 = n21952 | n21954;
  assign n51896 = n22215 & n51837;
  assign n51897 = n21952 & n22215;
  assign n67598 = (n51720 & n51896) | (n51720 & n51897) | (n51896 & n51897);
  assign n67599 = (n51896 & n51897) | (n51896 & n67480) | (n51897 & n67480);
  assign n67600 = (n67373 & n67598) | (n67373 & n67599) | (n67598 & n67599);
  assign n51899 = n22215 | n51837;
  assign n51900 = n21952 | n22215;
  assign n67601 = (n51720 & n51899) | (n51720 & n51900) | (n51899 & n51900);
  assign n67602 = (n51899 & n51900) | (n51899 & n67480) | (n51900 & n67480);
  assign n67603 = (n67373 & n67601) | (n67373 & n67602) | (n67601 & n67602);
  assign n22218 = ~n67600 & n67603;
  assign n22219 = x135 & x187;
  assign n22220 = n22218 & n22219;
  assign n22221 = n22218 | n22219;
  assign n22222 = ~n22220 & n22221;
  assign n51902 = n21959 & n22222;
  assign n67604 = (n22222 & n51778) | (n22222 & n51902) | (n51778 & n51902);
  assign n67605 = (n22222 & n51779) | (n22222 & n51902) | (n51779 & n51902);
  assign n67606 = (n51617 & n67604) | (n51617 & n67605) | (n67604 & n67605);
  assign n51904 = n21959 | n22222;
  assign n67607 = n51778 | n51904;
  assign n67608 = n51779 | n51904;
  assign n67609 = (n51617 & n67607) | (n51617 & n67608) | (n67607 & n67608);
  assign n22225 = ~n67606 & n67609;
  assign n22226 = x134 & x188;
  assign n22227 = n22225 & n22226;
  assign n22228 = n22225 | n22226;
  assign n22229 = ~n22227 & n22228;
  assign n51835 = n21966 | n21968;
  assign n67610 = n22229 & n51835;
  assign n67554 = n21713 | n21966;
  assign n67555 = (n21966 & n21968) | (n21966 & n67554) | (n21968 & n67554);
  assign n67611 = n22229 & n67555;
  assign n67612 = (n67459 & n67610) | (n67459 & n67611) | (n67610 & n67611);
  assign n67613 = n22229 | n51835;
  assign n67614 = n22229 | n67555;
  assign n67615 = (n67459 & n67613) | (n67459 & n67614) | (n67613 & n67614);
  assign n22232 = ~n67612 & n67615;
  assign n22233 = x133 & x189;
  assign n22234 = n22232 & n22233;
  assign n22235 = n22232 | n22233;
  assign n22236 = ~n22234 & n22235;
  assign n51906 = n21973 & n22236;
  assign n67616 = (n22236 & n51788) | (n22236 & n51906) | (n51788 & n51906);
  assign n67617 = (n21975 & n22236) | (n21975 & n51906) | (n22236 & n51906);
  assign n67618 = (n51678 & n67616) | (n51678 & n67617) | (n67616 & n67617);
  assign n51908 = n21973 | n22236;
  assign n67619 = n51788 | n51908;
  assign n67620 = n21975 | n51908;
  assign n67621 = (n51678 & n67619) | (n51678 & n67620) | (n67619 & n67620);
  assign n22239 = ~n67618 & n67621;
  assign n22240 = x132 & x190;
  assign n22241 = n22239 & n22240;
  assign n22242 = n22239 | n22240;
  assign n22243 = ~n22241 & n22242;
  assign n51910 = n21980 & n22243;
  assign n51911 = (n22243 & n51793) | (n22243 & n51910) | (n51793 & n51910);
  assign n51912 = n21980 | n22243;
  assign n51913 = n51793 | n51912;
  assign n22246 = ~n51911 & n51913;
  assign n22247 = x131 & x191;
  assign n22248 = n22246 & n22247;
  assign n22249 = n22246 | n22247;
  assign n22250 = ~n22248 & n22249;
  assign n51914 = n21987 & n22250;
  assign n51915 = (n22250 & n51797) | (n22250 & n51914) | (n51797 & n51914);
  assign n51916 = n21987 | n22250;
  assign n51917 = n51797 | n51916;
  assign n22253 = ~n51915 & n51917;
  assign n22254 = x130 & x192;
  assign n22255 = n22253 & n22254;
  assign n22256 = n22253 | n22254;
  assign n22257 = ~n22255 & n22256;
  assign n51918 = n21994 & n22257;
  assign n51919 = (n22257 & n51802) | (n22257 & n51918) | (n51802 & n51918);
  assign n51920 = n21994 | n22257;
  assign n51921 = n51802 | n51920;
  assign n22260 = ~n51919 & n51921;
  assign n22261 = x129 & x193;
  assign n22262 = n22260 & n22261;
  assign n22263 = n22260 | n22261;
  assign n22264 = ~n22262 & n22263;
  assign n51832 = n22001 | n22003;
  assign n51922 = n22264 & n51832;
  assign n51923 = n22001 & n22264;
  assign n51924 = (n51714 & n51922) | (n51714 & n51923) | (n51922 & n51923);
  assign n51925 = n22264 | n51832;
  assign n51926 = n22001 | n22264;
  assign n51927 = (n51714 & n51925) | (n51714 & n51926) | (n51925 & n51926);
  assign n22267 = ~n51924 & n51927;
  assign n22268 = x128 & x194;
  assign n22269 = n22267 & n22268;
  assign n22270 = n22267 | n22268;
  assign n22271 = ~n22269 & n22270;
  assign n51830 = n22008 | n22010;
  assign n67622 = n22271 & n51830;
  assign n67623 = n22008 & n22271;
  assign n67624 = (n51712 & n67622) | (n51712 & n67623) | (n67622 & n67623);
  assign n67625 = n22271 | n51830;
  assign n67626 = n22008 | n22271;
  assign n67627 = (n51712 & n67625) | (n51712 & n67626) | (n67625 & n67626);
  assign n22274 = ~n67624 & n67627;
  assign n22275 = x127 & x195;
  assign n22276 = n22274 & n22275;
  assign n22277 = n22274 | n22275;
  assign n22278 = ~n22276 & n22277;
  assign n51828 = n22015 | n22017;
  assign n67628 = n22278 & n51828;
  assign n67629 = n22015 & n22278;
  assign n67630 = (n51710 & n67628) | (n51710 & n67629) | (n67628 & n67629);
  assign n67631 = n22278 | n51828;
  assign n67632 = n22015 | n22278;
  assign n67633 = (n51710 & n67631) | (n51710 & n67632) | (n67631 & n67632);
  assign n22281 = ~n67630 & n67633;
  assign n22282 = x126 & x196;
  assign n22283 = n22281 & n22282;
  assign n22284 = n22281 | n22282;
  assign n22285 = ~n22283 & n22284;
  assign n22286 = n51827 & n22285;
  assign n22287 = n51827 | n22285;
  assign n22288 = ~n22286 & n22287;
  assign n22289 = x125 & x197;
  assign n22290 = n22288 & n22289;
  assign n22291 = n22288 | n22289;
  assign n22292 = ~n22290 & n22291;
  assign n22293 = n51825 & n22292;
  assign n22294 = n51825 | n22292;
  assign n22295 = ~n22293 & n22294;
  assign n22296 = x124 & x198;
  assign n22297 = n22295 & n22296;
  assign n22298 = n22295 | n22296;
  assign n22299 = ~n22297 & n22298;
  assign n22300 = n51823 & n22299;
  assign n22301 = n51823 | n22299;
  assign n22302 = ~n22300 & n22301;
  assign n22303 = x123 & x199;
  assign n22304 = n22302 & n22303;
  assign n22305 = n22302 | n22303;
  assign n22306 = ~n22304 & n22305;
  assign n22307 = n51821 & n22306;
  assign n22308 = n51821 | n22306;
  assign n22309 = ~n22307 & n22308;
  assign n22310 = x122 & x200;
  assign n22311 = n22309 & n22310;
  assign n22312 = n22309 | n22310;
  assign n22313 = ~n22311 & n22312;
  assign n22314 = n51819 & n22313;
  assign n22315 = n51819 | n22313;
  assign n22316 = ~n22314 & n22315;
  assign n22317 = x121 & x201;
  assign n22318 = n22316 & n22317;
  assign n22319 = n22316 | n22317;
  assign n22320 = ~n22318 & n22319;
  assign n22321 = n51817 & n22320;
  assign n22322 = n51817 | n22320;
  assign n22323 = ~n22321 & n22322;
  assign n22324 = x120 & x202;
  assign n22325 = n22323 & n22324;
  assign n22326 = n22323 | n22324;
  assign n22327 = ~n22325 & n22326;
  assign n22328 = n22122 & n22327;
  assign n22329 = n22122 | n22327;
  assign n22330 = ~n22328 & n22329;
  assign n22331 = x119 & x203;
  assign n22332 = n22330 & n22331;
  assign n22333 = n22330 | n22331;
  assign n22334 = ~n22332 & n22333;
  assign n22335 = n67553 & n22334;
  assign n22336 = n67553 | n22334;
  assign n22337 = ~n22335 & n22336;
  assign n22338 = x118 & x204;
  assign n22339 = n22337 & n22338;
  assign n22340 = n22337 | n22338;
  assign n22341 = ~n22339 & n22340;
  assign n22342 = n51815 & n22341;
  assign n22343 = n51815 | n22341;
  assign n22344 = ~n22342 & n22343;
  assign n22345 = x117 & x205;
  assign n22346 = n22344 & n22345;
  assign n22347 = n22344 | n22345;
  assign n22348 = ~n22346 & n22347;
  assign n22349 = n51813 & n22348;
  assign n22350 = n51813 | n22348;
  assign n22351 = ~n22349 & n22350;
  assign n22352 = x116 & x206;
  assign n22353 = n22351 & n22352;
  assign n22354 = n22351 | n22352;
  assign n22355 = ~n22353 & n22354;
  assign n22356 = n51811 & n22355;
  assign n22357 = n51811 | n22355;
  assign n22358 = ~n22356 & n22357;
  assign n22359 = x115 & x207;
  assign n22360 = n22358 & n22359;
  assign n22361 = n22358 | n22359;
  assign n22362 = ~n22360 & n22361;
  assign n22363 = n51809 & n22362;
  assign n22364 = n51809 | n22362;
  assign n22365 = ~n22363 & n22364;
  assign n22366 = x114 & x208;
  assign n22367 = n22365 & n22366;
  assign n22368 = n22365 | n22366;
  assign n22369 = ~n22367 & n22368;
  assign n22370 = n51807 & n22369;
  assign n22371 = n51807 | n22369;
  assign n22372 = ~n22370 & n22371;
  assign n22373 = x113 & x209;
  assign n22374 = n22372 & n22373;
  assign n22375 = n22372 | n22373;
  assign n22376 = ~n22374 & n22375;
  assign n22377 = n22113 & n22376;
  assign n22378 = n22113 | n22376;
  assign n22379 = ~n22377 & n22378;
  assign n22380 = x112 & x210;
  assign n22381 = n22379 & n22380;
  assign n22382 = n22379 | n22380;
  assign n22383 = ~n22381 & n22382;
  assign n67634 = n22113 | n22373;
  assign n67635 = (n22113 & n22372) | (n22113 & n67634) | (n22372 & n67634);
  assign n51929 = (n22374 & n22376) | (n22374 & n67635) | (n22376 & n67635);
  assign n51930 = n22367 | n51807;
  assign n51931 = (n22367 & n22369) | (n22367 & n51930) | (n22369 & n51930);
  assign n51932 = n22360 | n51809;
  assign n51933 = (n22360 & n22362) | (n22360 & n51932) | (n22362 & n51932);
  assign n51934 = n22353 | n51811;
  assign n51935 = (n22353 & n22355) | (n22353 & n51934) | (n22355 & n51934);
  assign n51936 = n22346 | n51813;
  assign n51937 = (n22346 & n22348) | (n22346 & n51936) | (n22348 & n51936);
  assign n51938 = n22339 | n51815;
  assign n51939 = (n22339 & n22341) | (n22339 & n51938) | (n22341 & n51938);
  assign n67636 = n22332 | n67553;
  assign n67637 = (n22332 & n22334) | (n22332 & n67636) | (n22334 & n67636);
  assign n51940 = n22325 | n22327;
  assign n51941 = (n22122 & n22325) | (n22122 & n51940) | (n22325 & n51940);
  assign n51942 = n22318 | n22320;
  assign n51943 = (n22318 & n51817) | (n22318 & n51942) | (n51817 & n51942);
  assign n51944 = n22311 | n22313;
  assign n51945 = (n22311 & n51819) | (n22311 & n51944) | (n51819 & n51944);
  assign n51946 = n22304 | n22306;
  assign n51947 = (n22304 & n51821) | (n22304 & n51946) | (n51821 & n51946);
  assign n51948 = n22297 | n22299;
  assign n51949 = (n22297 & n51823) | (n22297 & n51948) | (n51823 & n51948);
  assign n51950 = n22290 | n22292;
  assign n51951 = (n22290 & n51825) | (n22290 & n51950) | (n51825 & n51950);
  assign n51829 = (n22015 & n51710) | (n22015 & n51828) | (n51710 & n51828);
  assign n51831 = (n22008 & n51712) | (n22008 & n51830) | (n51712 & n51830);
  assign n51836 = (n67459 & n67555) | (n67459 & n51835) | (n67555 & n51835);
  assign n51961 = n22220 | n22222;
  assign n67638 = n21959 | n22220;
  assign n67639 = (n22220 & n22222) | (n22220 & n67638) | (n22222 & n67638);
  assign n67640 = (n51778 & n51961) | (n51778 & n67639) | (n51961 & n67639);
  assign n67641 = (n51779 & n51961) | (n51779 & n67639) | (n51961 & n67639);
  assign n67642 = (n51617 & n67640) | (n51617 & n67641) | (n67640 & n67641);
  assign n51729 = (n51513 & n67484) | (n51513 & n51728) | (n67484 & n51728);
  assign n22417 = x147 & x176;
  assign n22418 = x146 & x177;
  assign n22419 = n22417 & n22418;
  assign n22420 = n22417 | n22418;
  assign n22421 = ~n22419 & n22420;
  assign n67649 = n22150 | n67568;
  assign n67652 = n22421 & n67649;
  assign n67650 = n22150 | n22152;
  assign n67653 = n22421 & n67650;
  assign n67654 = (n67489 & n67652) | (n67489 & n67653) | (n67652 & n67653);
  assign n67655 = n22150 & n22421;
  assign n67656 = (n22421 & n67573) | (n22421 & n67655) | (n67573 & n67655);
  assign n67657 = (n51436 & n67654) | (n51436 & n67656) | (n67654 & n67656);
  assign n67658 = (n67253 & n67654) | (n67253 & n67656) | (n67654 & n67656);
  assign n67659 = (n66988 & n67657) | (n66988 & n67658) | (n67657 & n67658);
  assign n67660 = n22421 | n67649;
  assign n67661 = n22421 | n67650;
  assign n67662 = (n67489 & n67660) | (n67489 & n67661) | (n67660 & n67661);
  assign n67663 = n22150 | n22421;
  assign n67664 = n67573 | n67663;
  assign n67665 = (n51436 & n67662) | (n51436 & n67664) | (n67662 & n67664);
  assign n67666 = (n67253 & n67662) | (n67253 & n67664) | (n67662 & n67664);
  assign n67667 = (n66988 & n67665) | (n66988 & n67666) | (n67665 & n67666);
  assign n22424 = ~n67659 & n67667;
  assign n22425 = x145 & x178;
  assign n22426 = n22424 & n22425;
  assign n22427 = n22424 | n22425;
  assign n22428 = ~n22426 & n22427;
  assign n67668 = n22157 | n22159;
  assign n67669 = (n22157 & n67585) | (n22157 & n67668) | (n67585 & n67668);
  assign n51991 = n22428 & n67669;
  assign n67670 = (n22157 & n51853) | (n22157 & n67668) | (n51853 & n67668);
  assign n51992 = n22428 & n67670;
  assign n51993 = (n67426 & n51991) | (n67426 & n51992) | (n51991 & n51992);
  assign n51994 = n22428 | n67669;
  assign n51995 = n22428 | n67670;
  assign n51996 = (n67426 & n51994) | (n67426 & n51995) | (n51994 & n51995);
  assign n22431 = ~n51993 & n51996;
  assign n22432 = x144 & x179;
  assign n22433 = n22431 & n22432;
  assign n22434 = n22431 | n22432;
  assign n22435 = ~n22433 & n22434;
  assign n51977 = n22164 | n67587;
  assign n67671 = n22435 & n51977;
  assign n67647 = n22164 | n22166;
  assign n67648 = (n22164 & n67589) | (n22164 & n67647) | (n67589 & n67647);
  assign n67672 = n22435 & n67648;
  assign n67673 = (n67407 & n67671) | (n67407 & n67672) | (n67671 & n67672);
  assign n67674 = n22435 | n51977;
  assign n67675 = n22435 | n67648;
  assign n67676 = (n67407 & n67674) | (n67407 & n67675) | (n67674 & n67675);
  assign n22438 = ~n67673 & n67676;
  assign n22439 = x143 & x180;
  assign n22440 = n22438 & n22439;
  assign n22441 = n22438 | n22439;
  assign n22442 = ~n22440 & n22441;
  assign n67677 = n21910 | n22171;
  assign n67678 = (n22171 & n22173) | (n22171 & n67677) | (n22173 & n67677);
  assign n51997 = n22442 & n67678;
  assign n51974 = n22171 | n22173;
  assign n51998 = n22442 & n51974;
  assign n51999 = (n67504 & n51997) | (n67504 & n51998) | (n51997 & n51998);
  assign n52000 = n22442 | n67678;
  assign n52001 = n22442 | n51974;
  assign n52002 = (n67504 & n52000) | (n67504 & n52001) | (n52000 & n52001);
  assign n22445 = ~n51999 & n52002;
  assign n22446 = x142 & x181;
  assign n22447 = n22445 & n22446;
  assign n22448 = n22445 | n22446;
  assign n22449 = ~n22447 & n22448;
  assign n51971 = n22178 | n22180;
  assign n52003 = n22449 & n51971;
  assign n52004 = n22178 & n22449;
  assign n52005 = (n67567 & n52003) | (n67567 & n52004) | (n52003 & n52004);
  assign n52006 = n22449 | n51971;
  assign n52007 = n22178 | n22449;
  assign n52008 = (n67567 & n52006) | (n67567 & n52007) | (n52006 & n52007);
  assign n22452 = ~n52005 & n52008;
  assign n22453 = x141 & x182;
  assign n22454 = n22452 & n22453;
  assign n22455 = n22452 | n22453;
  assign n22456 = ~n22454 & n22455;
  assign n51969 = n22185 | n51880;
  assign n67679 = n22456 & n51969;
  assign n67645 = n21924 | n22185;
  assign n67646 = (n22185 & n22187) | (n22185 & n67645) | (n22187 & n67645);
  assign n67680 = n22456 & n67646;
  assign n67681 = (n51729 & n67679) | (n51729 & n67680) | (n67679 & n67680);
  assign n67682 = n22456 | n51969;
  assign n67683 = n22456 | n67646;
  assign n67684 = (n51729 & n67682) | (n51729 & n67683) | (n67682 & n67683);
  assign n22459 = ~n67681 & n67684;
  assign n22460 = x140 & x183;
  assign n22461 = n22459 & n22460;
  assign n22462 = n22459 | n22460;
  assign n22463 = ~n22461 & n22462;
  assign n52009 = n22192 & n22463;
  assign n67685 = (n22463 & n51886) | (n22463 & n52009) | (n51886 & n52009);
  assign n67686 = (n22463 & n51887) | (n22463 & n52009) | (n51887 & n52009);
  assign n67687 = (n51726 & n67685) | (n51726 & n67686) | (n67685 & n67686);
  assign n52011 = n22192 | n22463;
  assign n67688 = n51886 | n52011;
  assign n67689 = n51887 | n52011;
  assign n67690 = (n51726 & n67688) | (n51726 & n67689) | (n67688 & n67689);
  assign n22466 = ~n67687 & n67690;
  assign n22467 = x139 & x184;
  assign n22468 = n22466 & n22467;
  assign n22469 = n22466 | n22467;
  assign n22470 = ~n22468 & n22469;
  assign n51966 = n22199 | n22201;
  assign n67691 = n22470 & n51966;
  assign n67643 = n21938 | n22199;
  assign n67644 = (n22199 & n22201) | (n22199 & n67643) | (n22201 & n67643);
  assign n67692 = n22470 & n67644;
  assign n67693 = (n51770 & n67691) | (n51770 & n67692) | (n67691 & n67692);
  assign n67694 = n22470 | n51966;
  assign n67695 = n22470 | n67644;
  assign n67696 = (n51770 & n67694) | (n51770 & n67695) | (n67694 & n67695);
  assign n22473 = ~n67693 & n67696;
  assign n22474 = x138 & x185;
  assign n22475 = n22473 & n22474;
  assign n22476 = n22473 | n22474;
  assign n22477 = ~n22475 & n22476;
  assign n51963 = n22206 | n22208;
  assign n52013 = n22477 & n51963;
  assign n52014 = n22206 & n22477;
  assign n52015 = (n67560 & n52013) | (n67560 & n52014) | (n52013 & n52014);
  assign n52016 = n22477 | n51963;
  assign n52017 = n22206 | n22477;
  assign n52018 = (n67560 & n52016) | (n67560 & n52017) | (n52016 & n52017);
  assign n22480 = ~n52015 & n52018;
  assign n22481 = x137 & x186;
  assign n22482 = n22480 & n22481;
  assign n22483 = n22480 | n22481;
  assign n22484 = ~n22482 & n22483;
  assign n52019 = n22213 & n22484;
  assign n52020 = (n22484 & n67600) | (n22484 & n52019) | (n67600 & n52019);
  assign n52021 = n22213 | n22484;
  assign n52022 = n67600 | n52021;
  assign n22487 = ~n52020 & n52022;
  assign n22488 = x136 & x187;
  assign n22489 = n22487 & n22488;
  assign n22490 = n22487 | n22488;
  assign n22491 = ~n22489 & n22490;
  assign n22492 = n67642 & n22491;
  assign n22493 = n67642 | n22491;
  assign n22494 = ~n22492 & n22493;
  assign n22495 = x135 & x188;
  assign n22496 = n22494 & n22495;
  assign n22497 = n22494 | n22495;
  assign n22498 = ~n22496 & n22497;
  assign n51958 = n22227 | n22229;
  assign n52023 = n22498 & n51958;
  assign n52024 = n22227 & n22498;
  assign n52025 = (n51836 & n52023) | (n51836 & n52024) | (n52023 & n52024);
  assign n52026 = n22498 | n51958;
  assign n52027 = n22227 | n22498;
  assign n52028 = (n51836 & n52026) | (n51836 & n52027) | (n52026 & n52027);
  assign n22501 = ~n52025 & n52028;
  assign n22502 = x134 & x189;
  assign n22503 = n22501 & n22502;
  assign n22504 = n22501 | n22502;
  assign n22505 = ~n22503 & n22504;
  assign n52029 = n22234 & n22505;
  assign n52030 = (n22505 & n67618) | (n22505 & n52029) | (n67618 & n52029);
  assign n52031 = n22234 | n22505;
  assign n52032 = n67618 | n52031;
  assign n22508 = ~n52030 & n52032;
  assign n22509 = x133 & x190;
  assign n22510 = n22508 & n22509;
  assign n22511 = n22508 | n22509;
  assign n22512 = ~n22510 & n22511;
  assign n52033 = n22241 & n22512;
  assign n52034 = (n22512 & n51911) | (n22512 & n52033) | (n51911 & n52033);
  assign n52035 = n22241 | n22512;
  assign n52036 = n51911 | n52035;
  assign n22515 = ~n52034 & n52036;
  assign n22516 = x132 & x191;
  assign n22517 = n22515 & n22516;
  assign n22518 = n22515 | n22516;
  assign n22519 = ~n22517 & n22518;
  assign n52037 = n22248 & n22519;
  assign n52038 = (n22519 & n51915) | (n22519 & n52037) | (n51915 & n52037);
  assign n52039 = n22248 | n22519;
  assign n52040 = n51915 | n52039;
  assign n22522 = ~n52038 & n52040;
  assign n22523 = x131 & x192;
  assign n22524 = n22522 & n22523;
  assign n22525 = n22522 | n22523;
  assign n22526 = ~n22524 & n22525;
  assign n52041 = n22255 & n22526;
  assign n52042 = (n22526 & n51919) | (n22526 & n52041) | (n51919 & n52041);
  assign n52043 = n22255 | n22526;
  assign n52044 = n51919 | n52043;
  assign n22529 = ~n52042 & n52044;
  assign n22530 = x130 & x193;
  assign n22531 = n22529 & n22530;
  assign n22532 = n22529 | n22530;
  assign n22533 = ~n22531 & n22532;
  assign n52045 = n22262 & n22533;
  assign n52046 = (n22533 & n51924) | (n22533 & n52045) | (n51924 & n52045);
  assign n52047 = n22262 | n22533;
  assign n52048 = n51924 | n52047;
  assign n22536 = ~n52046 & n52048;
  assign n22537 = x129 & x194;
  assign n22538 = n22536 & n22537;
  assign n22539 = n22536 | n22537;
  assign n22540 = ~n22538 & n22539;
  assign n51956 = n22269 | n22271;
  assign n52049 = n22540 & n51956;
  assign n52050 = n22269 & n22540;
  assign n52051 = (n51831 & n52049) | (n51831 & n52050) | (n52049 & n52050);
  assign n52052 = n22540 | n51956;
  assign n52053 = n22269 | n22540;
  assign n52054 = (n51831 & n52052) | (n51831 & n52053) | (n52052 & n52053);
  assign n22543 = ~n52051 & n52054;
  assign n22544 = x128 & x195;
  assign n22545 = n22543 & n22544;
  assign n22546 = n22543 | n22544;
  assign n22547 = ~n22545 & n22546;
  assign n51954 = n22276 | n22278;
  assign n67697 = n22547 & n51954;
  assign n67698 = n22276 & n22547;
  assign n67699 = (n51829 & n67697) | (n51829 & n67698) | (n67697 & n67698);
  assign n67700 = n22547 | n51954;
  assign n67701 = n22276 | n22547;
  assign n67702 = (n51829 & n67700) | (n51829 & n67701) | (n67700 & n67701);
  assign n22550 = ~n67699 & n67702;
  assign n22551 = x127 & x196;
  assign n22552 = n22550 & n22551;
  assign n22553 = n22550 | n22551;
  assign n22554 = ~n22552 & n22553;
  assign n51952 = n22283 | n22285;
  assign n67703 = n22554 & n51952;
  assign n67704 = n22283 & n22554;
  assign n67705 = (n51827 & n67703) | (n51827 & n67704) | (n67703 & n67704);
  assign n67706 = n22554 | n51952;
  assign n67707 = n22283 | n22554;
  assign n67708 = (n51827 & n67706) | (n51827 & n67707) | (n67706 & n67707);
  assign n22557 = ~n67705 & n67708;
  assign n22558 = x126 & x197;
  assign n22559 = n22557 & n22558;
  assign n22560 = n22557 | n22558;
  assign n22561 = ~n22559 & n22560;
  assign n22562 = n51951 & n22561;
  assign n22563 = n51951 | n22561;
  assign n22564 = ~n22562 & n22563;
  assign n22565 = x125 & x198;
  assign n22566 = n22564 & n22565;
  assign n22567 = n22564 | n22565;
  assign n22568 = ~n22566 & n22567;
  assign n22569 = n51949 & n22568;
  assign n22570 = n51949 | n22568;
  assign n22571 = ~n22569 & n22570;
  assign n22572 = x124 & x199;
  assign n22573 = n22571 & n22572;
  assign n22574 = n22571 | n22572;
  assign n22575 = ~n22573 & n22574;
  assign n22576 = n51947 & n22575;
  assign n22577 = n51947 | n22575;
  assign n22578 = ~n22576 & n22577;
  assign n22579 = x123 & x200;
  assign n22580 = n22578 & n22579;
  assign n22581 = n22578 | n22579;
  assign n22582 = ~n22580 & n22581;
  assign n22583 = n51945 & n22582;
  assign n22584 = n51945 | n22582;
  assign n22585 = ~n22583 & n22584;
  assign n22586 = x122 & x201;
  assign n22587 = n22585 & n22586;
  assign n22588 = n22585 | n22586;
  assign n22589 = ~n22587 & n22588;
  assign n22590 = n51943 & n22589;
  assign n22591 = n51943 | n22589;
  assign n22592 = ~n22590 & n22591;
  assign n22593 = x121 & x202;
  assign n22594 = n22592 & n22593;
  assign n22595 = n22592 | n22593;
  assign n22596 = ~n22594 & n22595;
  assign n22597 = n51941 & n22596;
  assign n22598 = n51941 | n22596;
  assign n22599 = ~n22597 & n22598;
  assign n22600 = x120 & x203;
  assign n22601 = n22599 & n22600;
  assign n22602 = n22599 | n22600;
  assign n22603 = ~n22601 & n22602;
  assign n22604 = n67637 & n22603;
  assign n22605 = n67637 | n22603;
  assign n22606 = ~n22604 & n22605;
  assign n22607 = x119 & x204;
  assign n22608 = n22606 & n22607;
  assign n22609 = n22606 | n22607;
  assign n22610 = ~n22608 & n22609;
  assign n22611 = n51939 & n22610;
  assign n22612 = n51939 | n22610;
  assign n22613 = ~n22611 & n22612;
  assign n22614 = x118 & x205;
  assign n22615 = n22613 & n22614;
  assign n22616 = n22613 | n22614;
  assign n22617 = ~n22615 & n22616;
  assign n22618 = n51937 & n22617;
  assign n22619 = n51937 | n22617;
  assign n22620 = ~n22618 & n22619;
  assign n22621 = x117 & x206;
  assign n22622 = n22620 & n22621;
  assign n22623 = n22620 | n22621;
  assign n22624 = ~n22622 & n22623;
  assign n22625 = n51935 & n22624;
  assign n22626 = n51935 | n22624;
  assign n22627 = ~n22625 & n22626;
  assign n22628 = x116 & x207;
  assign n22629 = n22627 & n22628;
  assign n22630 = n22627 | n22628;
  assign n22631 = ~n22629 & n22630;
  assign n22632 = n51933 & n22631;
  assign n22633 = n51933 | n22631;
  assign n22634 = ~n22632 & n22633;
  assign n22635 = x115 & x208;
  assign n22636 = n22634 & n22635;
  assign n22637 = n22634 | n22635;
  assign n22638 = ~n22636 & n22637;
  assign n22639 = n51931 & n22638;
  assign n22640 = n51931 | n22638;
  assign n22641 = ~n22639 & n22640;
  assign n22642 = x114 & x209;
  assign n22643 = n22641 & n22642;
  assign n22644 = n22641 | n22642;
  assign n22645 = ~n22643 & n22644;
  assign n22646 = n51929 & n22645;
  assign n22647 = n51929 | n22645;
  assign n22648 = ~n22646 & n22647;
  assign n22649 = x113 & x210;
  assign n22650 = n22648 & n22649;
  assign n22651 = n22648 | n22649;
  assign n22652 = ~n22650 & n22651;
  assign n22653 = n22381 & n22652;
  assign n22654 = n22381 | n22652;
  assign n22655 = ~n22653 & n22654;
  assign n22656 = x112 & x211;
  assign n22657 = n22655 & n22656;
  assign n22658 = n22655 | n22656;
  assign n22659 = ~n22657 & n22658;
  assign n52055 = n22381 | n22650;
  assign n52056 = (n22650 & n22652) | (n22650 & n52055) | (n22652 & n52055);
  assign n52057 = n22643 | n51929;
  assign n52058 = (n22643 & n22645) | (n22643 & n52057) | (n22645 & n52057);
  assign n52059 = n22636 | n51931;
  assign n52060 = (n22636 & n22638) | (n22636 & n52059) | (n22638 & n52059);
  assign n52061 = n22629 | n51933;
  assign n52062 = (n22629 & n22631) | (n22629 & n52061) | (n22631 & n52061);
  assign n52063 = n22622 | n51935;
  assign n52064 = (n22622 & n22624) | (n22622 & n52063) | (n22624 & n52063);
  assign n52065 = n22615 | n51937;
  assign n52066 = (n22615 & n22617) | (n22615 & n52065) | (n22617 & n52065);
  assign n52067 = n22608 | n51939;
  assign n52068 = (n22608 & n22610) | (n22608 & n52067) | (n22610 & n52067);
  assign n52069 = n22601 | n22603;
  assign n52070 = (n67637 & n22601) | (n67637 & n52069) | (n22601 & n52069);
  assign n52071 = n22594 | n22596;
  assign n52072 = (n22594 & n51941) | (n22594 & n52071) | (n51941 & n52071);
  assign n52073 = n22587 | n22589;
  assign n52074 = (n22587 & n51943) | (n22587 & n52073) | (n51943 & n52073);
  assign n52075 = n22580 | n22582;
  assign n52076 = (n22580 & n51945) | (n22580 & n52075) | (n51945 & n52075);
  assign n52077 = n22573 | n22575;
  assign n52078 = (n22573 & n51947) | (n22573 & n52077) | (n51947 & n52077);
  assign n52079 = n22566 | n22568;
  assign n52080 = (n22566 & n51949) | (n22566 & n52079) | (n51949 & n52079);
  assign n51953 = (n22283 & n51827) | (n22283 & n51952) | (n51827 & n51952);
  assign n51955 = (n22276 & n51829) | (n22276 & n51954) | (n51829 & n51954);
  assign n51967 = (n51770 & n67644) | (n51770 & n51966) | (n67644 & n51966);
  assign n52098 = n22461 | n22463;
  assign n67713 = n22192 | n22461;
  assign n67714 = (n22461 & n22463) | (n22461 & n67713) | (n22463 & n67713);
  assign n67715 = (n51886 & n52098) | (n51886 & n67714) | (n52098 & n67714);
  assign n67716 = (n51887 & n52098) | (n51887 & n67714) | (n52098 & n67714);
  assign n67717 = (n51726 & n67715) | (n51726 & n67716) | (n67715 & n67716);
  assign n22694 = x148 & x176;
  assign n22695 = x147 & x177;
  assign n22696 = n22694 & n22695;
  assign n22697 = n22694 | n22695;
  assign n22698 = ~n22696 & n22697;
  assign n52113 = n22419 & n22698;
  assign n67728 = (n22698 & n52113) | (n22698 & n67658) | (n52113 & n67658);
  assign n67729 = (n22698 & n52113) | (n22698 & n67657) | (n52113 & n67657);
  assign n67730 = (n66988 & n67728) | (n66988 & n67729) | (n67728 & n67729);
  assign n52115 = n22419 | n22698;
  assign n67731 = n52115 | n67658;
  assign n67732 = n52115 | n67657;
  assign n67733 = (n66988 & n67731) | (n66988 & n67732) | (n67731 & n67732);
  assign n22701 = ~n67730 & n67733;
  assign n22702 = x146 & x178;
  assign n22703 = n22701 & n22702;
  assign n22704 = n22701 | n22702;
  assign n22705 = ~n22703 & n22704;
  assign n67725 = n22426 | n22428;
  assign n67727 = (n22426 & n67670) | (n22426 & n67725) | (n67670 & n67725);
  assign n67734 = n22705 & n67727;
  assign n67726 = (n22426 & n67669) | (n22426 & n67725) | (n67669 & n67725);
  assign n67735 = n22705 & n67726;
  assign n67736 = (n67426 & n67734) | (n67426 & n67735) | (n67734 & n67735);
  assign n67737 = n22705 | n67727;
  assign n67738 = n22705 | n67726;
  assign n67739 = (n67426 & n67737) | (n67426 & n67738) | (n67737 & n67738);
  assign n22708 = ~n67736 & n67739;
  assign n22709 = x145 & x179;
  assign n22710 = n22708 & n22709;
  assign n22711 = n22708 | n22709;
  assign n22712 = ~n22710 & n22711;
  assign n52108 = n22433 | n22435;
  assign n52117 = n22712 & n52108;
  assign n52118 = n22433 & n22712;
  assign n67740 = (n51977 & n52117) | (n51977 & n52118) | (n52117 & n52118);
  assign n67741 = (n52117 & n52118) | (n52117 & n67648) | (n52118 & n67648);
  assign n67742 = (n67407 & n67740) | (n67407 & n67741) | (n67740 & n67741);
  assign n52120 = n22712 | n52108;
  assign n52121 = n22433 | n22712;
  assign n67743 = (n51977 & n52120) | (n51977 & n52121) | (n52120 & n52121);
  assign n67744 = (n52120 & n52121) | (n52120 & n67648) | (n52121 & n67648);
  assign n67745 = (n67407 & n67743) | (n67407 & n67744) | (n67743 & n67744);
  assign n22715 = ~n67742 & n67745;
  assign n22716 = x144 & x180;
  assign n22717 = n22715 & n22716;
  assign n22718 = n22715 | n22716;
  assign n22719 = ~n22717 & n22718;
  assign n67722 = n22440 | n22442;
  assign n67724 = (n22440 & n51974) | (n22440 & n67722) | (n51974 & n67722);
  assign n67746 = n22719 & n67724;
  assign n67723 = (n22440 & n67678) | (n22440 & n67722) | (n67678 & n67722);
  assign n67747 = n22719 & n67723;
  assign n67748 = (n67504 & n67746) | (n67504 & n67747) | (n67746 & n67747);
  assign n67749 = n22719 | n67724;
  assign n67750 = n22719 | n67723;
  assign n67751 = (n67504 & n67749) | (n67504 & n67750) | (n67749 & n67750);
  assign n22722 = ~n67748 & n67751;
  assign n22723 = x143 & x181;
  assign n22724 = n22722 & n22723;
  assign n22725 = n22722 | n22723;
  assign n22726 = ~n22724 & n22725;
  assign n67718 = n22447 | n22449;
  assign n67719 = (n22447 & n51971) | (n22447 & n67718) | (n51971 & n67718);
  assign n67752 = n22726 & n67719;
  assign n67720 = n22178 | n22447;
  assign n67721 = (n22447 & n22449) | (n22447 & n67720) | (n22449 & n67720);
  assign n67753 = n22726 & n67721;
  assign n67754 = (n67567 & n67752) | (n67567 & n67753) | (n67752 & n67753);
  assign n67755 = n22726 | n67719;
  assign n67756 = n22726 | n67721;
  assign n67757 = (n67567 & n67755) | (n67567 & n67756) | (n67755 & n67756);
  assign n22729 = ~n67754 & n67757;
  assign n22730 = x142 & x182;
  assign n22731 = n22729 & n22730;
  assign n22732 = n22729 | n22730;
  assign n22733 = ~n22731 & n22732;
  assign n52100 = n22454 | n22456;
  assign n52123 = n22733 & n52100;
  assign n52124 = n22454 & n22733;
  assign n67758 = (n51969 & n52123) | (n51969 & n52124) | (n52123 & n52124);
  assign n67759 = (n52123 & n52124) | (n52123 & n67646) | (n52124 & n67646);
  assign n67760 = (n51729 & n67758) | (n51729 & n67759) | (n67758 & n67759);
  assign n52126 = n22733 | n52100;
  assign n52127 = n22454 | n22733;
  assign n67761 = (n51969 & n52126) | (n51969 & n52127) | (n52126 & n52127);
  assign n67762 = (n52126 & n52127) | (n52126 & n67646) | (n52127 & n67646);
  assign n67763 = (n51729 & n67761) | (n51729 & n67762) | (n67761 & n67762);
  assign n22736 = ~n67760 & n67763;
  assign n22737 = x141 & x183;
  assign n22738 = n22736 & n22737;
  assign n22739 = n22736 | n22737;
  assign n22740 = ~n22738 & n22739;
  assign n22741 = n67717 & n22740;
  assign n22742 = n67717 | n22740;
  assign n22743 = ~n22741 & n22742;
  assign n22744 = x140 & x184;
  assign n22745 = n22743 & n22744;
  assign n22746 = n22743 | n22744;
  assign n22747 = ~n22745 & n22746;
  assign n52095 = n22468 | n22470;
  assign n52129 = n22747 & n52095;
  assign n52130 = n22468 & n22747;
  assign n52131 = (n51967 & n52129) | (n51967 & n52130) | (n52129 & n52130);
  assign n52132 = n22747 | n52095;
  assign n52133 = n22468 | n22747;
  assign n52134 = (n51967 & n52132) | (n51967 & n52133) | (n52132 & n52133);
  assign n22750 = ~n52131 & n52134;
  assign n22751 = x139 & x185;
  assign n22752 = n22750 & n22751;
  assign n22753 = n22750 | n22751;
  assign n22754 = ~n22752 & n22753;
  assign n52135 = n22475 & n22754;
  assign n52136 = (n22754 & n52015) | (n22754 & n52135) | (n52015 & n52135);
  assign n52137 = n22475 | n22754;
  assign n52138 = n52015 | n52137;
  assign n22757 = ~n52136 & n52138;
  assign n22758 = x138 & x186;
  assign n22759 = n22757 & n22758;
  assign n22760 = n22757 | n22758;
  assign n22761 = ~n22759 & n22760;
  assign n52093 = n22482 | n22484;
  assign n67764 = n22761 & n52093;
  assign n67711 = n22213 | n22482;
  assign n67712 = (n22482 & n22484) | (n22482 & n67711) | (n22484 & n67711);
  assign n67765 = n22761 & n67712;
  assign n67766 = (n67600 & n67764) | (n67600 & n67765) | (n67764 & n67765);
  assign n67767 = n22761 | n52093;
  assign n67768 = n22761 | n67712;
  assign n67769 = (n67600 & n67767) | (n67600 & n67768) | (n67767 & n67768);
  assign n22764 = ~n67766 & n67769;
  assign n22765 = x137 & x187;
  assign n22766 = n22764 & n22765;
  assign n22767 = n22764 | n22765;
  assign n22768 = ~n22766 & n22767;
  assign n52090 = n22489 | n22491;
  assign n52139 = n22768 & n52090;
  assign n52140 = n22489 & n22768;
  assign n52141 = (n67642 & n52139) | (n67642 & n52140) | (n52139 & n52140);
  assign n52142 = n22768 | n52090;
  assign n52143 = n22489 | n22768;
  assign n52144 = (n67642 & n52142) | (n67642 & n52143) | (n52142 & n52143);
  assign n22771 = ~n52141 & n52144;
  assign n22772 = x136 & x188;
  assign n22773 = n22771 & n22772;
  assign n22774 = n22771 | n22772;
  assign n22775 = ~n22773 & n22774;
  assign n52145 = n22496 & n22775;
  assign n67770 = (n22775 & n52024) | (n22775 & n52145) | (n52024 & n52145);
  assign n67771 = (n22775 & n52023) | (n22775 & n52145) | (n52023 & n52145);
  assign n67772 = (n51836 & n67770) | (n51836 & n67771) | (n67770 & n67771);
  assign n52147 = n22496 | n22775;
  assign n67773 = n52024 | n52147;
  assign n67774 = n52023 | n52147;
  assign n67775 = (n51836 & n67773) | (n51836 & n67774) | (n67773 & n67774);
  assign n22778 = ~n67772 & n67775;
  assign n22779 = x135 & x189;
  assign n22780 = n22778 & n22779;
  assign n22781 = n22778 | n22779;
  assign n22782 = ~n22780 & n22781;
  assign n52088 = n22503 | n22505;
  assign n67776 = n22782 & n52088;
  assign n67709 = n22234 | n22503;
  assign n67710 = (n22503 & n22505) | (n22503 & n67709) | (n22505 & n67709);
  assign n67777 = n22782 & n67710;
  assign n67778 = (n67618 & n67776) | (n67618 & n67777) | (n67776 & n67777);
  assign n67779 = n22782 | n52088;
  assign n67780 = n22782 | n67710;
  assign n67781 = (n67618 & n67779) | (n67618 & n67780) | (n67779 & n67780);
  assign n22785 = ~n67778 & n67781;
  assign n22786 = x134 & x190;
  assign n22787 = n22785 & n22786;
  assign n22788 = n22785 | n22786;
  assign n22789 = ~n22787 & n22788;
  assign n52149 = n22510 & n22789;
  assign n67782 = (n22789 & n52033) | (n22789 & n52149) | (n52033 & n52149);
  assign n67783 = (n22512 & n22789) | (n22512 & n52149) | (n22789 & n52149);
  assign n67784 = (n51911 & n67782) | (n51911 & n67783) | (n67782 & n67783);
  assign n52151 = n22510 | n22789;
  assign n67785 = n52033 | n52151;
  assign n67786 = n22512 | n52151;
  assign n67787 = (n51911 & n67785) | (n51911 & n67786) | (n67785 & n67786);
  assign n22792 = ~n67784 & n67787;
  assign n22793 = x133 & x191;
  assign n22794 = n22792 & n22793;
  assign n22795 = n22792 | n22793;
  assign n22796 = ~n22794 & n22795;
  assign n52153 = n22517 & n22796;
  assign n52154 = (n22796 & n52038) | (n22796 & n52153) | (n52038 & n52153);
  assign n52155 = n22517 | n22796;
  assign n52156 = n52038 | n52155;
  assign n22799 = ~n52154 & n52156;
  assign n22800 = x132 & x192;
  assign n22801 = n22799 & n22800;
  assign n22802 = n22799 | n22800;
  assign n22803 = ~n22801 & n22802;
  assign n52157 = n22524 & n22803;
  assign n52158 = (n22803 & n52042) | (n22803 & n52157) | (n52042 & n52157);
  assign n52159 = n22524 | n22803;
  assign n52160 = n52042 | n52159;
  assign n22806 = ~n52158 & n52160;
  assign n22807 = x131 & x193;
  assign n22808 = n22806 & n22807;
  assign n22809 = n22806 | n22807;
  assign n22810 = ~n22808 & n22809;
  assign n52161 = n22531 & n22810;
  assign n52162 = (n22810 & n52046) | (n22810 & n52161) | (n52046 & n52161);
  assign n52163 = n22531 | n22810;
  assign n52164 = n52046 | n52163;
  assign n22813 = ~n52162 & n52164;
  assign n22814 = x130 & x194;
  assign n22815 = n22813 & n22814;
  assign n22816 = n22813 | n22814;
  assign n22817 = ~n22815 & n22816;
  assign n52165 = n22538 & n22817;
  assign n52166 = (n22817 & n52051) | (n22817 & n52165) | (n52051 & n52165);
  assign n52167 = n22538 | n22817;
  assign n52168 = n52051 | n52167;
  assign n22820 = ~n52166 & n52168;
  assign n22821 = x129 & x195;
  assign n22822 = n22820 & n22821;
  assign n22823 = n22820 | n22821;
  assign n22824 = ~n22822 & n22823;
  assign n52085 = n22545 | n22547;
  assign n52169 = n22824 & n52085;
  assign n52170 = n22545 & n22824;
  assign n52171 = (n51955 & n52169) | (n51955 & n52170) | (n52169 & n52170);
  assign n52172 = n22824 | n52085;
  assign n52173 = n22545 | n22824;
  assign n52174 = (n51955 & n52172) | (n51955 & n52173) | (n52172 & n52173);
  assign n22827 = ~n52171 & n52174;
  assign n22828 = x128 & x196;
  assign n22829 = n22827 & n22828;
  assign n22830 = n22827 | n22828;
  assign n22831 = ~n22829 & n22830;
  assign n52083 = n22552 | n22554;
  assign n67788 = n22831 & n52083;
  assign n67789 = n22552 & n22831;
  assign n67790 = (n51953 & n67788) | (n51953 & n67789) | (n67788 & n67789);
  assign n67791 = n22831 | n52083;
  assign n67792 = n22552 | n22831;
  assign n67793 = (n51953 & n67791) | (n51953 & n67792) | (n67791 & n67792);
  assign n22834 = ~n67790 & n67793;
  assign n22835 = x127 & x197;
  assign n22836 = n22834 & n22835;
  assign n22837 = n22834 | n22835;
  assign n22838 = ~n22836 & n22837;
  assign n52081 = n22559 | n22561;
  assign n67794 = n22838 & n52081;
  assign n67795 = n22559 & n22838;
  assign n67796 = (n51951 & n67794) | (n51951 & n67795) | (n67794 & n67795);
  assign n67797 = n22838 | n52081;
  assign n67798 = n22559 | n22838;
  assign n67799 = (n51951 & n67797) | (n51951 & n67798) | (n67797 & n67798);
  assign n22841 = ~n67796 & n67799;
  assign n22842 = x126 & x198;
  assign n22843 = n22841 & n22842;
  assign n22844 = n22841 | n22842;
  assign n22845 = ~n22843 & n22844;
  assign n22846 = n52080 & n22845;
  assign n22847 = n52080 | n22845;
  assign n22848 = ~n22846 & n22847;
  assign n22849 = x125 & x199;
  assign n22850 = n22848 & n22849;
  assign n22851 = n22848 | n22849;
  assign n22852 = ~n22850 & n22851;
  assign n22853 = n52078 & n22852;
  assign n22854 = n52078 | n22852;
  assign n22855 = ~n22853 & n22854;
  assign n22856 = x124 & x200;
  assign n22857 = n22855 & n22856;
  assign n22858 = n22855 | n22856;
  assign n22859 = ~n22857 & n22858;
  assign n22860 = n52076 & n22859;
  assign n22861 = n52076 | n22859;
  assign n22862 = ~n22860 & n22861;
  assign n22863 = x123 & x201;
  assign n22864 = n22862 & n22863;
  assign n22865 = n22862 | n22863;
  assign n22866 = ~n22864 & n22865;
  assign n22867 = n52074 & n22866;
  assign n22868 = n52074 | n22866;
  assign n22869 = ~n22867 & n22868;
  assign n22870 = x122 & x202;
  assign n22871 = n22869 & n22870;
  assign n22872 = n22869 | n22870;
  assign n22873 = ~n22871 & n22872;
  assign n22874 = n52072 & n22873;
  assign n22875 = n52072 | n22873;
  assign n22876 = ~n22874 & n22875;
  assign n22877 = x121 & x203;
  assign n22878 = n22876 & n22877;
  assign n22879 = n22876 | n22877;
  assign n22880 = ~n22878 & n22879;
  assign n22881 = n52070 & n22880;
  assign n22882 = n52070 | n22880;
  assign n22883 = ~n22881 & n22882;
  assign n22884 = x120 & x204;
  assign n22885 = n22883 & n22884;
  assign n22886 = n22883 | n22884;
  assign n22887 = ~n22885 & n22886;
  assign n22888 = n52068 & n22887;
  assign n22889 = n52068 | n22887;
  assign n22890 = ~n22888 & n22889;
  assign n22891 = x119 & x205;
  assign n22892 = n22890 & n22891;
  assign n22893 = n22890 | n22891;
  assign n22894 = ~n22892 & n22893;
  assign n22895 = n52066 & n22894;
  assign n22896 = n52066 | n22894;
  assign n22897 = ~n22895 & n22896;
  assign n22898 = x118 & x206;
  assign n22899 = n22897 & n22898;
  assign n22900 = n22897 | n22898;
  assign n22901 = ~n22899 & n22900;
  assign n22902 = n52064 & n22901;
  assign n22903 = n52064 | n22901;
  assign n22904 = ~n22902 & n22903;
  assign n22905 = x117 & x207;
  assign n22906 = n22904 & n22905;
  assign n22907 = n22904 | n22905;
  assign n22908 = ~n22906 & n22907;
  assign n22909 = n52062 & n22908;
  assign n22910 = n52062 | n22908;
  assign n22911 = ~n22909 & n22910;
  assign n22912 = x116 & x208;
  assign n22913 = n22911 & n22912;
  assign n22914 = n22911 | n22912;
  assign n22915 = ~n22913 & n22914;
  assign n22916 = n52060 & n22915;
  assign n22917 = n52060 | n22915;
  assign n22918 = ~n22916 & n22917;
  assign n22919 = x115 & x209;
  assign n22920 = n22918 & n22919;
  assign n22921 = n22918 | n22919;
  assign n22922 = ~n22920 & n22921;
  assign n22923 = n52058 & n22922;
  assign n22924 = n52058 | n22922;
  assign n22925 = ~n22923 & n22924;
  assign n22926 = x114 & x210;
  assign n22927 = n22925 & n22926;
  assign n22928 = n22925 | n22926;
  assign n22929 = ~n22927 & n22928;
  assign n22930 = n52056 & n22929;
  assign n22931 = n52056 | n22929;
  assign n22932 = ~n22930 & n22931;
  assign n22933 = x113 & x211;
  assign n22934 = n22932 & n22933;
  assign n22935 = n22932 | n22933;
  assign n22936 = ~n22934 & n22935;
  assign n22937 = n22657 & n22936;
  assign n22938 = n22657 | n22936;
  assign n22939 = ~n22937 & n22938;
  assign n22940 = x112 & x212;
  assign n22941 = n22939 & n22940;
  assign n22942 = n22939 | n22940;
  assign n22943 = ~n22941 & n22942;
  assign n67800 = n22657 | n22933;
  assign n67801 = (n22657 & n22932) | (n22657 & n67800) | (n22932 & n67800);
  assign n52176 = (n22934 & n22936) | (n22934 & n67801) | (n22936 & n67801);
  assign n67802 = n22927 | n52056;
  assign n67803 = (n22927 & n22929) | (n22927 & n67802) | (n22929 & n67802);
  assign n22946 = n22920 | n22923;
  assign n22947 = n22913 | n22916;
  assign n22948 = n22906 | n22909;
  assign n22949 = n22899 | n22902;
  assign n22950 = n22892 | n22895;
  assign n22951 = n22885 | n22888;
  assign n52177 = n22878 | n22880;
  assign n52178 = (n22878 & n52070) | (n22878 & n52177) | (n52070 & n52177);
  assign n52179 = n22871 | n22873;
  assign n52180 = (n22871 & n52072) | (n22871 & n52179) | (n52072 & n52179);
  assign n52181 = n22864 | n22866;
  assign n52182 = (n22864 & n52074) | (n22864 & n52181) | (n52074 & n52181);
  assign n52183 = n22857 | n22859;
  assign n52184 = (n22857 & n52076) | (n22857 & n52183) | (n52076 & n52183);
  assign n52185 = n22850 | n22852;
  assign n52186 = (n22850 & n52078) | (n22850 & n52185) | (n52078 & n52185);
  assign n52082 = (n22559 & n51951) | (n22559 & n52081) | (n51951 & n52081);
  assign n52084 = (n22552 & n51953) | (n22552 & n52083) | (n51953 & n52083);
  assign n52089 = (n67618 & n67710) | (n67618 & n52088) | (n67710 & n52088);
  assign n52196 = n22773 | n22775;
  assign n67804 = n22496 | n22773;
  assign n67805 = (n22773 & n22775) | (n22773 & n67804) | (n22775 & n67804);
  assign n67806 = (n52024 & n52196) | (n52024 & n67805) | (n52196 & n67805);
  assign n67807 = (n52023 & n52196) | (n52023 & n67805) | (n52196 & n67805);
  assign n67808 = (n51836 & n67806) | (n51836 & n67807) | (n67806 & n67807);
  assign n52094 = (n67600 & n67712) | (n67600 & n52093) | (n67712 & n52093);
  assign n67811 = n22454 | n22731;
  assign n67812 = (n22731 & n22733) | (n22731 & n67811) | (n22733 & n67811);
  assign n67813 = n22731 | n22733;
  assign n67814 = (n22731 & n52100) | (n22731 & n67813) | (n52100 & n67813);
  assign n67815 = (n51969 & n67812) | (n51969 & n67814) | (n67812 & n67814);
  assign n67816 = (n67646 & n67812) | (n67646 & n67814) | (n67812 & n67814);
  assign n67817 = (n51729 & n67815) | (n51729 & n67816) | (n67815 & n67816);
  assign n22979 = x149 & x176;
  assign n22980 = x148 & x177;
  assign n22981 = n22979 & n22980;
  assign n22982 = n22979 | n22980;
  assign n22983 = ~n22981 & n22982;
  assign n67818 = n22419 | n22696;
  assign n67819 = (n22696 & n22698) | (n22696 & n67818) | (n22698 & n67818);
  assign n52220 = n22983 & n67819;
  assign n52218 = n22696 | n22698;
  assign n52221 = n22983 & n52218;
  assign n67820 = (n52220 & n52221) | (n52220 & n67658) | (n52221 & n67658);
  assign n67821 = (n52220 & n52221) | (n52220 & n67657) | (n52221 & n67657);
  assign n67822 = (n66988 & n67820) | (n66988 & n67821) | (n67820 & n67821);
  assign n52223 = n22983 | n67819;
  assign n52224 = n22983 | n52218;
  assign n67823 = (n52223 & n52224) | (n52223 & n67658) | (n52224 & n67658);
  assign n67824 = (n52223 & n52224) | (n52223 & n67657) | (n52224 & n67657);
  assign n67825 = (n66988 & n67823) | (n66988 & n67824) | (n67823 & n67824);
  assign n22986 = ~n67822 & n67825;
  assign n22987 = x147 & x178;
  assign n22988 = n22986 & n22987;
  assign n22989 = n22986 | n22987;
  assign n22990 = ~n22988 & n22989;
  assign n52215 = n22703 | n22705;
  assign n52226 = n22990 & n52215;
  assign n52227 = n22703 & n22990;
  assign n67826 = (n52226 & n52227) | (n52226 & n67727) | (n52227 & n67727);
  assign n67827 = (n52226 & n52227) | (n52226 & n67726) | (n52227 & n67726);
  assign n67828 = (n67426 & n67826) | (n67426 & n67827) | (n67826 & n67827);
  assign n52229 = n22990 | n52215;
  assign n52230 = n22703 | n22990;
  assign n67829 = (n52229 & n52230) | (n52229 & n67727) | (n52230 & n67727);
  assign n67830 = (n52229 & n52230) | (n52229 & n67726) | (n52230 & n67726);
  assign n67831 = (n67426 & n67829) | (n67426 & n67830) | (n67829 & n67830);
  assign n22993 = ~n67828 & n67831;
  assign n22994 = x146 & x179;
  assign n22995 = n22993 & n22994;
  assign n22996 = n22993 | n22994;
  assign n22997 = ~n22995 & n22996;
  assign n67832 = n22710 | n22712;
  assign n67833 = (n22710 & n52108) | (n22710 & n67832) | (n52108 & n67832);
  assign n52232 = n22997 & n67833;
  assign n67834 = n22433 | n22710;
  assign n67835 = (n22710 & n22712) | (n22710 & n67834) | (n22712 & n67834);
  assign n52233 = n22997 & n67835;
  assign n67836 = (n51977 & n52232) | (n51977 & n52233) | (n52232 & n52233);
  assign n67837 = (n52232 & n52233) | (n52232 & n67648) | (n52233 & n67648);
  assign n67838 = (n67407 & n67836) | (n67407 & n67837) | (n67836 & n67837);
  assign n52235 = n22997 | n67833;
  assign n52236 = n22997 | n67835;
  assign n67839 = (n51977 & n52235) | (n51977 & n52236) | (n52235 & n52236);
  assign n67840 = (n52235 & n52236) | (n52235 & n67648) | (n52236 & n67648);
  assign n67841 = (n67407 & n67839) | (n67407 & n67840) | (n67839 & n67840);
  assign n23000 = ~n67838 & n67841;
  assign n23001 = x145 & x180;
  assign n23002 = n23000 & n23001;
  assign n23003 = n23000 | n23001;
  assign n23004 = ~n23002 & n23003;
  assign n52210 = n22717 | n22719;
  assign n52238 = n23004 & n52210;
  assign n52239 = n22717 & n23004;
  assign n67842 = (n52238 & n52239) | (n52238 & n67724) | (n52239 & n67724);
  assign n67843 = (n52238 & n52239) | (n52238 & n67723) | (n52239 & n67723);
  assign n67844 = (n67504 & n67842) | (n67504 & n67843) | (n67842 & n67843);
  assign n52241 = n23004 | n52210;
  assign n52242 = n22717 | n23004;
  assign n67845 = (n52241 & n52242) | (n52241 & n67724) | (n52242 & n67724);
  assign n67846 = (n52241 & n52242) | (n52241 & n67723) | (n52242 & n67723);
  assign n67847 = (n67504 & n67845) | (n67504 & n67846) | (n67845 & n67846);
  assign n23007 = ~n67844 & n67847;
  assign n23008 = x144 & x181;
  assign n23009 = n23007 & n23008;
  assign n23010 = n23007 | n23008;
  assign n23011 = ~n23009 & n23010;
  assign n52208 = n22724 | n22726;
  assign n52244 = n23011 & n52208;
  assign n52245 = n22724 & n23011;
  assign n67848 = (n52244 & n52245) | (n52244 & n67719) | (n52245 & n67719);
  assign n67849 = (n52244 & n52245) | (n52244 & n67721) | (n52245 & n67721);
  assign n67850 = (n67567 & n67848) | (n67567 & n67849) | (n67848 & n67849);
  assign n52247 = n23011 | n52208;
  assign n52248 = n22724 | n23011;
  assign n67851 = (n52247 & n52248) | (n52247 & n67719) | (n52248 & n67719);
  assign n67852 = (n52247 & n52248) | (n52247 & n67721) | (n52248 & n67721);
  assign n67853 = (n67567 & n67851) | (n67567 & n67852) | (n67851 & n67852);
  assign n23014 = ~n67850 & n67853;
  assign n23015 = x143 & x182;
  assign n23016 = n23014 & n23015;
  assign n23017 = n23014 | n23015;
  assign n23018 = ~n23016 & n23017;
  assign n23019 = n67817 & n23018;
  assign n23020 = n67817 | n23018;
  assign n23021 = ~n23019 & n23020;
  assign n23022 = x142 & x183;
  assign n23023 = n23021 & n23022;
  assign n23024 = n23021 | n23022;
  assign n23025 = ~n23023 & n23024;
  assign n52203 = n22738 | n22740;
  assign n52250 = n23025 & n52203;
  assign n52251 = n22738 & n23025;
  assign n52252 = (n67717 & n52250) | (n67717 & n52251) | (n52250 & n52251);
  assign n52253 = n23025 | n52203;
  assign n52254 = n22738 | n23025;
  assign n52255 = (n67717 & n52253) | (n67717 & n52254) | (n52253 & n52254);
  assign n23028 = ~n52252 & n52255;
  assign n23029 = x141 & x184;
  assign n23030 = n23028 & n23029;
  assign n23031 = n23028 | n23029;
  assign n23032 = ~n23030 & n23031;
  assign n52256 = n22745 & n23032;
  assign n67854 = (n23032 & n52130) | (n23032 & n52256) | (n52130 & n52256);
  assign n67855 = (n23032 & n52129) | (n23032 & n52256) | (n52129 & n52256);
  assign n67856 = (n51967 & n67854) | (n51967 & n67855) | (n67854 & n67855);
  assign n52258 = n22745 | n23032;
  assign n67857 = n52130 | n52258;
  assign n67858 = n52129 | n52258;
  assign n67859 = (n51967 & n67857) | (n51967 & n67858) | (n67857 & n67858);
  assign n23035 = ~n67856 & n67859;
  assign n23036 = x140 & x185;
  assign n23037 = n23035 & n23036;
  assign n23038 = n23035 | n23036;
  assign n23039 = ~n23037 & n23038;
  assign n52201 = n22752 | n22754;
  assign n67860 = n23039 & n52201;
  assign n67809 = n22475 | n22752;
  assign n67810 = (n22752 & n22754) | (n22752 & n67809) | (n22754 & n67809);
  assign n67861 = n23039 & n67810;
  assign n67862 = (n52015 & n67860) | (n52015 & n67861) | (n67860 & n67861);
  assign n67863 = n23039 | n52201;
  assign n67864 = n23039 | n67810;
  assign n67865 = (n52015 & n67863) | (n52015 & n67864) | (n67863 & n67864);
  assign n23042 = ~n67862 & n67865;
  assign n23043 = x139 & x186;
  assign n23044 = n23042 & n23043;
  assign n23045 = n23042 | n23043;
  assign n23046 = ~n23044 & n23045;
  assign n52198 = n22759 | n22761;
  assign n52260 = n23046 & n52198;
  assign n52261 = n22759 & n23046;
  assign n52262 = (n52094 & n52260) | (n52094 & n52261) | (n52260 & n52261);
  assign n52263 = n23046 | n52198;
  assign n52264 = n22759 | n23046;
  assign n52265 = (n52094 & n52263) | (n52094 & n52264) | (n52263 & n52264);
  assign n23049 = ~n52262 & n52265;
  assign n23050 = x138 & x187;
  assign n23051 = n23049 & n23050;
  assign n23052 = n23049 | n23050;
  assign n23053 = ~n23051 & n23052;
  assign n52266 = n22766 & n23053;
  assign n67866 = (n23053 & n52139) | (n23053 & n52266) | (n52139 & n52266);
  assign n67867 = (n23053 & n52140) | (n23053 & n52266) | (n52140 & n52266);
  assign n67868 = (n67642 & n67866) | (n67642 & n67867) | (n67866 & n67867);
  assign n52268 = n22766 | n23053;
  assign n67869 = n52139 | n52268;
  assign n67870 = n52140 | n52268;
  assign n67871 = (n67642 & n67869) | (n67642 & n67870) | (n67869 & n67870);
  assign n23056 = ~n67868 & n67871;
  assign n23057 = x137 & x188;
  assign n23058 = n23056 & n23057;
  assign n23059 = n23056 | n23057;
  assign n23060 = ~n23058 & n23059;
  assign n23061 = n67808 & n23060;
  assign n23062 = n67808 | n23060;
  assign n23063 = ~n23061 & n23062;
  assign n23064 = x136 & x189;
  assign n23065 = n23063 & n23064;
  assign n23066 = n23063 | n23064;
  assign n23067 = ~n23065 & n23066;
  assign n52193 = n22780 | n22782;
  assign n52270 = n23067 & n52193;
  assign n52271 = n22780 & n23067;
  assign n52272 = (n52089 & n52270) | (n52089 & n52271) | (n52270 & n52271);
  assign n52273 = n23067 | n52193;
  assign n52274 = n22780 | n23067;
  assign n52275 = (n52089 & n52273) | (n52089 & n52274) | (n52273 & n52274);
  assign n23070 = ~n52272 & n52275;
  assign n23071 = x135 & x190;
  assign n23072 = n23070 & n23071;
  assign n23073 = n23070 | n23071;
  assign n23074 = ~n23072 & n23073;
  assign n52276 = n22787 & n23074;
  assign n52277 = (n23074 & n67784) | (n23074 & n52276) | (n67784 & n52276);
  assign n52278 = n22787 | n23074;
  assign n52279 = n67784 | n52278;
  assign n23077 = ~n52277 & n52279;
  assign n23078 = x134 & x191;
  assign n23079 = n23077 & n23078;
  assign n23080 = n23077 | n23078;
  assign n23081 = ~n23079 & n23080;
  assign n52280 = n22794 & n23081;
  assign n52281 = (n23081 & n52154) | (n23081 & n52280) | (n52154 & n52280);
  assign n52282 = n22794 | n23081;
  assign n52283 = n52154 | n52282;
  assign n23084 = ~n52281 & n52283;
  assign n23085 = x133 & x192;
  assign n23086 = n23084 & n23085;
  assign n23087 = n23084 | n23085;
  assign n23088 = ~n23086 & n23087;
  assign n52284 = n22801 & n23088;
  assign n52285 = (n23088 & n52158) | (n23088 & n52284) | (n52158 & n52284);
  assign n52286 = n22801 | n23088;
  assign n52287 = n52158 | n52286;
  assign n23091 = ~n52285 & n52287;
  assign n23092 = x132 & x193;
  assign n23093 = n23091 & n23092;
  assign n23094 = n23091 | n23092;
  assign n23095 = ~n23093 & n23094;
  assign n52288 = n22808 & n23095;
  assign n52289 = (n23095 & n52162) | (n23095 & n52288) | (n52162 & n52288);
  assign n52290 = n22808 | n23095;
  assign n52291 = n52162 | n52290;
  assign n23098 = ~n52289 & n52291;
  assign n23099 = x131 & x194;
  assign n23100 = n23098 & n23099;
  assign n23101 = n23098 | n23099;
  assign n23102 = ~n23100 & n23101;
  assign n52292 = n22815 & n23102;
  assign n52293 = (n23102 & n52166) | (n23102 & n52292) | (n52166 & n52292);
  assign n52294 = n22815 | n23102;
  assign n52295 = n52166 | n52294;
  assign n23105 = ~n52293 & n52295;
  assign n23106 = x130 & x195;
  assign n23107 = n23105 & n23106;
  assign n23108 = n23105 | n23106;
  assign n23109 = ~n23107 & n23108;
  assign n52296 = n22822 & n23109;
  assign n52297 = (n23109 & n52171) | (n23109 & n52296) | (n52171 & n52296);
  assign n52298 = n22822 | n23109;
  assign n52299 = n52171 | n52298;
  assign n23112 = ~n52297 & n52299;
  assign n23113 = x129 & x196;
  assign n23114 = n23112 & n23113;
  assign n23115 = n23112 | n23113;
  assign n23116 = ~n23114 & n23115;
  assign n52191 = n22829 | n22831;
  assign n52300 = n23116 & n52191;
  assign n52301 = n22829 & n23116;
  assign n52302 = (n52084 & n52300) | (n52084 & n52301) | (n52300 & n52301);
  assign n52303 = n23116 | n52191;
  assign n52304 = n22829 | n23116;
  assign n52305 = (n52084 & n52303) | (n52084 & n52304) | (n52303 & n52304);
  assign n23119 = ~n52302 & n52305;
  assign n23120 = x128 & x197;
  assign n23121 = n23119 & n23120;
  assign n23122 = n23119 | n23120;
  assign n23123 = ~n23121 & n23122;
  assign n52189 = n22836 | n22838;
  assign n67872 = n23123 & n52189;
  assign n67873 = n22836 & n23123;
  assign n67874 = (n52082 & n67872) | (n52082 & n67873) | (n67872 & n67873);
  assign n67875 = n23123 | n52189;
  assign n67876 = n22836 | n23123;
  assign n67877 = (n52082 & n67875) | (n52082 & n67876) | (n67875 & n67876);
  assign n23126 = ~n67874 & n67877;
  assign n23127 = x127 & x198;
  assign n23128 = n23126 & n23127;
  assign n23129 = n23126 | n23127;
  assign n23130 = ~n23128 & n23129;
  assign n52187 = n22843 | n22845;
  assign n67878 = n23130 & n52187;
  assign n67879 = n22843 & n23130;
  assign n67880 = (n52080 & n67878) | (n52080 & n67879) | (n67878 & n67879);
  assign n67881 = n23130 | n52187;
  assign n67882 = n22843 | n23130;
  assign n67883 = (n52080 & n67881) | (n52080 & n67882) | (n67881 & n67882);
  assign n23133 = ~n67880 & n67883;
  assign n23134 = x126 & x199;
  assign n23135 = n23133 & n23134;
  assign n23136 = n23133 | n23134;
  assign n23137 = ~n23135 & n23136;
  assign n23138 = n52186 & n23137;
  assign n23139 = n52186 | n23137;
  assign n23140 = ~n23138 & n23139;
  assign n23141 = x125 & x200;
  assign n23142 = n23140 & n23141;
  assign n23143 = n23140 | n23141;
  assign n23144 = ~n23142 & n23143;
  assign n23145 = n52184 & n23144;
  assign n23146 = n52184 | n23144;
  assign n23147 = ~n23145 & n23146;
  assign n23148 = x124 & x201;
  assign n23149 = n23147 & n23148;
  assign n23150 = n23147 | n23148;
  assign n23151 = ~n23149 & n23150;
  assign n23152 = n52182 & n23151;
  assign n23153 = n52182 | n23151;
  assign n23154 = ~n23152 & n23153;
  assign n23155 = x123 & x202;
  assign n23156 = n23154 & n23155;
  assign n23157 = n23154 | n23155;
  assign n23158 = ~n23156 & n23157;
  assign n23159 = n52180 & n23158;
  assign n23160 = n52180 | n23158;
  assign n23161 = ~n23159 & n23160;
  assign n23162 = x122 & x203;
  assign n23163 = n23161 & n23162;
  assign n23164 = n23161 | n23162;
  assign n23165 = ~n23163 & n23164;
  assign n23166 = n52178 & n23165;
  assign n23167 = n52178 | n23165;
  assign n23168 = ~n23166 & n23167;
  assign n23169 = x121 & x204;
  assign n23170 = n23168 & n23169;
  assign n23171 = n23168 | n23169;
  assign n23172 = ~n23170 & n23171;
  assign n23173 = n22951 & n23172;
  assign n23174 = n22951 | n23172;
  assign n23175 = ~n23173 & n23174;
  assign n23176 = x120 & x205;
  assign n23177 = n23175 & n23176;
  assign n23178 = n23175 | n23176;
  assign n23179 = ~n23177 & n23178;
  assign n23180 = n22950 & n23179;
  assign n23181 = n22950 | n23179;
  assign n23182 = ~n23180 & n23181;
  assign n23183 = x119 & x206;
  assign n23184 = n23182 & n23183;
  assign n23185 = n23182 | n23183;
  assign n23186 = ~n23184 & n23185;
  assign n23187 = n22949 & n23186;
  assign n23188 = n22949 | n23186;
  assign n23189 = ~n23187 & n23188;
  assign n23190 = x118 & x207;
  assign n23191 = n23189 & n23190;
  assign n23192 = n23189 | n23190;
  assign n23193 = ~n23191 & n23192;
  assign n23194 = n22948 & n23193;
  assign n23195 = n22948 | n23193;
  assign n23196 = ~n23194 & n23195;
  assign n23197 = x117 & x208;
  assign n23198 = n23196 & n23197;
  assign n23199 = n23196 | n23197;
  assign n23200 = ~n23198 & n23199;
  assign n23201 = n22947 & n23200;
  assign n23202 = n22947 | n23200;
  assign n23203 = ~n23201 & n23202;
  assign n23204 = x116 & x209;
  assign n23205 = n23203 & n23204;
  assign n23206 = n23203 | n23204;
  assign n23207 = ~n23205 & n23206;
  assign n23208 = n22946 & n23207;
  assign n23209 = n22946 | n23207;
  assign n23210 = ~n23208 & n23209;
  assign n23211 = x115 & x210;
  assign n23212 = n23210 & n23211;
  assign n23213 = n23210 | n23211;
  assign n23214 = ~n23212 & n23213;
  assign n23215 = n67803 & n23214;
  assign n23216 = n67803 | n23214;
  assign n23217 = ~n23215 & n23216;
  assign n23218 = x114 & x211;
  assign n23219 = n23217 & n23218;
  assign n23220 = n23217 | n23218;
  assign n23221 = ~n23219 & n23220;
  assign n23222 = n52176 & n23221;
  assign n23223 = n52176 | n23221;
  assign n23224 = ~n23222 & n23223;
  assign n23225 = x113 & x212;
  assign n23226 = n23224 & n23225;
  assign n23227 = n23224 | n23225;
  assign n23228 = ~n23226 & n23227;
  assign n23229 = n22941 & n23228;
  assign n23230 = n22941 | n23228;
  assign n23231 = ~n23229 & n23230;
  assign n23232 = x112 & x213;
  assign n23233 = n23231 & n23232;
  assign n23234 = n23231 | n23232;
  assign n23235 = ~n23233 & n23234;
  assign n67884 = n22941 | n23225;
  assign n67885 = (n22941 & n23224) | (n22941 & n67884) | (n23224 & n67884);
  assign n52307 = (n23226 & n23228) | (n23226 & n67885) | (n23228 & n67885);
  assign n52308 = n23219 | n52176;
  assign n52309 = (n23219 & n23221) | (n23219 & n52308) | (n23221 & n52308);
  assign n67886 = n23212 | n67803;
  assign n67887 = (n23212 & n23214) | (n23212 & n67886) | (n23214 & n67886);
  assign n23239 = n23205 | n23208;
  assign n23240 = n23198 | n23201;
  assign n23241 = n23191 | n23194;
  assign n23242 = n23184 | n23187;
  assign n23243 = n23177 | n23180;
  assign n52310 = n23170 | n23172;
  assign n52311 = (n22951 & n23170) | (n22951 & n52310) | (n23170 & n52310);
  assign n52312 = n23163 | n23165;
  assign n52313 = (n23163 & n52178) | (n23163 & n52312) | (n52178 & n52312);
  assign n52314 = n23156 | n23158;
  assign n52315 = (n23156 & n52180) | (n23156 & n52314) | (n52180 & n52314);
  assign n52316 = n23149 | n23151;
  assign n52317 = (n23149 & n52182) | (n23149 & n52316) | (n52182 & n52316);
  assign n52318 = n23142 | n23144;
  assign n52319 = (n23142 & n52184) | (n23142 & n52318) | (n52184 & n52318);
  assign n52188 = (n22843 & n52080) | (n22843 & n52187) | (n52080 & n52187);
  assign n52190 = (n22836 & n52082) | (n22836 & n52189) | (n52082 & n52189);
  assign n52332 = n23051 | n23053;
  assign n67890 = n22766 | n23051;
  assign n67891 = (n23051 & n23053) | (n23051 & n67890) | (n23053 & n67890);
  assign n67892 = (n52139 & n52332) | (n52139 & n67891) | (n52332 & n67891);
  assign n67893 = (n52140 & n52332) | (n52140 & n67891) | (n52332 & n67891);
  assign n67894 = (n67642 & n67892) | (n67642 & n67893) | (n67892 & n67893);
  assign n52202 = (n52015 & n67810) | (n52015 & n52201) | (n67810 & n52201);
  assign n52337 = n23030 | n23032;
  assign n67895 = n22745 | n23030;
  assign n67896 = (n23030 & n23032) | (n23030 & n67895) | (n23032 & n67895);
  assign n67897 = (n52130 & n52337) | (n52130 & n67896) | (n52337 & n67896);
  assign n67898 = (n52129 & n52337) | (n52129 & n67896) | (n52337 & n67896);
  assign n67899 = (n51967 & n67897) | (n51967 & n67898) | (n67897 & n67898);
  assign n67900 = n22738 | n23023;
  assign n67901 = (n23023 & n23025) | (n23023 & n67900) | (n23025 & n67900);
  assign n52340 = n23023 | n52250;
  assign n52341 = (n67717 & n67901) | (n67717 & n52340) | (n67901 & n52340);
  assign n67902 = n23009 | n23011;
  assign n67903 = (n23009 & n52208) | (n23009 & n67902) | (n52208 & n67902);
  assign n67904 = n22724 | n23009;
  assign n67905 = (n23009 & n23011) | (n23009 & n67904) | (n23011 & n67904);
  assign n67906 = (n67719 & n67903) | (n67719 & n67905) | (n67903 & n67905);
  assign n67907 = (n67721 & n67903) | (n67721 & n67905) | (n67903 & n67905);
  assign n67908 = (n67567 & n67906) | (n67567 & n67907) | (n67906 & n67907);
  assign n67909 = n22995 | n22997;
  assign n67910 = (n22995 & n67835) | (n22995 & n67909) | (n67835 & n67909);
  assign n67911 = (n22995 & n67833) | (n22995 & n67909) | (n67833 & n67909);
  assign n67912 = (n51977 & n67910) | (n51977 & n67911) | (n67910 & n67911);
  assign n67913 = (n67648 & n67910) | (n67648 & n67911) | (n67910 & n67911);
  assign n67914 = (n67407 & n67912) | (n67407 & n67913) | (n67912 & n67913);
  assign n23272 = x150 & x176;
  assign n23273 = x149 & x177;
  assign n23274 = n23272 & n23273;
  assign n23275 = n23272 | n23273;
  assign n23276 = ~n23274 & n23275;
  assign n67915 = n22981 | n22983;
  assign n67916 = (n22981 & n67819) | (n22981 & n67915) | (n67819 & n67915);
  assign n52359 = n23276 & n67916;
  assign n67917 = (n22981 & n52218) | (n22981 & n67915) | (n52218 & n67915);
  assign n52360 = n23276 & n67917;
  assign n67918 = (n52359 & n52360) | (n52359 & n67658) | (n52360 & n67658);
  assign n67919 = (n52359 & n52360) | (n52359 & n67657) | (n52360 & n67657);
  assign n67920 = (n66988 & n67918) | (n66988 & n67919) | (n67918 & n67919);
  assign n52362 = n23276 | n67916;
  assign n52363 = n23276 | n67917;
  assign n67921 = (n52362 & n52363) | (n52362 & n67658) | (n52363 & n67658);
  assign n67922 = (n52362 & n52363) | (n52362 & n67657) | (n52363 & n67657);
  assign n67923 = (n66988 & n67921) | (n66988 & n67922) | (n67921 & n67922);
  assign n23279 = ~n67920 & n67923;
  assign n23280 = x148 & x178;
  assign n23281 = n23279 & n23280;
  assign n23282 = n23279 | n23280;
  assign n23283 = ~n23281 & n23282;
  assign n67924 = n22988 | n22990;
  assign n67925 = (n22988 & n52215) | (n22988 & n67924) | (n52215 & n67924);
  assign n52365 = n23283 & n67925;
  assign n67926 = n22703 | n22988;
  assign n67927 = (n22988 & n22990) | (n22988 & n67926) | (n22990 & n67926);
  assign n52366 = n23283 & n67927;
  assign n67928 = (n52365 & n52366) | (n52365 & n67727) | (n52366 & n67727);
  assign n67929 = (n52365 & n52366) | (n52365 & n67726) | (n52366 & n67726);
  assign n67930 = (n67426 & n67928) | (n67426 & n67929) | (n67928 & n67929);
  assign n52368 = n23283 | n67925;
  assign n52369 = n23283 | n67927;
  assign n67931 = (n52368 & n52369) | (n52368 & n67727) | (n52369 & n67727);
  assign n67932 = (n52368 & n52369) | (n52368 & n67726) | (n52369 & n67726);
  assign n67933 = (n67426 & n67931) | (n67426 & n67932) | (n67931 & n67932);
  assign n23286 = ~n67930 & n67933;
  assign n23287 = x147 & x179;
  assign n23288 = n23286 & n23287;
  assign n23289 = n23286 | n23287;
  assign n23290 = ~n23288 & n23289;
  assign n23291 = n67914 & n23290;
  assign n23292 = n67914 | n23290;
  assign n23293 = ~n23291 & n23292;
  assign n23294 = x146 & x180;
  assign n23295 = n23293 & n23294;
  assign n23296 = n23293 | n23294;
  assign n23297 = ~n23295 & n23296;
  assign n67934 = n23002 | n23004;
  assign n67935 = (n23002 & n52210) | (n23002 & n67934) | (n52210 & n67934);
  assign n52371 = n23297 & n67935;
  assign n67936 = n22717 | n23002;
  assign n67937 = (n23002 & n23004) | (n23002 & n67936) | (n23004 & n67936);
  assign n52372 = n23297 & n67937;
  assign n67938 = (n52371 & n52372) | (n52371 & n67724) | (n52372 & n67724);
  assign n67939 = (n52371 & n52372) | (n52371 & n67723) | (n52372 & n67723);
  assign n67940 = (n67504 & n67938) | (n67504 & n67939) | (n67938 & n67939);
  assign n52374 = n23297 | n67935;
  assign n52375 = n23297 | n67937;
  assign n67941 = (n52374 & n52375) | (n52374 & n67724) | (n52375 & n67724);
  assign n67942 = (n52374 & n52375) | (n52374 & n67723) | (n52375 & n67723);
  assign n67943 = (n67504 & n67941) | (n67504 & n67942) | (n67941 & n67942);
  assign n23300 = ~n67940 & n67943;
  assign n23301 = x145 & x181;
  assign n23302 = n23300 & n23301;
  assign n23303 = n23300 | n23301;
  assign n23304 = ~n23302 & n23303;
  assign n23305 = n67908 & n23304;
  assign n23306 = n67908 | n23304;
  assign n23307 = ~n23305 & n23306;
  assign n23308 = x144 & x182;
  assign n23309 = n23307 & n23308;
  assign n23310 = n23307 | n23308;
  assign n23311 = ~n23309 & n23310;
  assign n52342 = n23016 | n23018;
  assign n52377 = n23311 & n52342;
  assign n52378 = n23016 & n23311;
  assign n52379 = (n67817 & n52377) | (n67817 & n52378) | (n52377 & n52378);
  assign n52380 = n23311 | n52342;
  assign n52381 = n23016 | n23311;
  assign n52382 = (n67817 & n52380) | (n67817 & n52381) | (n52380 & n52381);
  assign n23314 = ~n52379 & n52382;
  assign n23315 = x143 & x183;
  assign n23316 = n23314 & n23315;
  assign n23317 = n23314 | n23315;
  assign n23318 = ~n23316 & n23317;
  assign n23319 = n52341 & n23318;
  assign n23320 = n52341 | n23318;
  assign n23321 = ~n23319 & n23320;
  assign n23322 = x142 & x184;
  assign n23323 = n23321 & n23322;
  assign n23324 = n23321 | n23322;
  assign n23325 = ~n23323 & n23324;
  assign n23326 = n67899 & n23325;
  assign n23327 = n67899 | n23325;
  assign n23328 = ~n23326 & n23327;
  assign n23329 = x141 & x185;
  assign n23330 = n23328 & n23329;
  assign n23331 = n23328 | n23329;
  assign n23332 = ~n23330 & n23331;
  assign n52334 = n23037 | n23039;
  assign n52383 = n23332 & n52334;
  assign n52384 = n23037 & n23332;
  assign n52385 = (n52202 & n52383) | (n52202 & n52384) | (n52383 & n52384);
  assign n52386 = n23332 | n52334;
  assign n52387 = n23037 | n23332;
  assign n52388 = (n52202 & n52386) | (n52202 & n52387) | (n52386 & n52387);
  assign n23335 = ~n52385 & n52388;
  assign n23336 = x140 & x186;
  assign n23337 = n23335 & n23336;
  assign n23338 = n23335 | n23336;
  assign n23339 = ~n23337 & n23338;
  assign n52389 = n23044 & n23339;
  assign n67944 = (n23339 & n52260) | (n23339 & n52389) | (n52260 & n52389);
  assign n67945 = (n23339 & n52261) | (n23339 & n52389) | (n52261 & n52389);
  assign n67946 = (n52094 & n67944) | (n52094 & n67945) | (n67944 & n67945);
  assign n52391 = n23044 | n23339;
  assign n67947 = n52260 | n52391;
  assign n67948 = n52261 | n52391;
  assign n67949 = (n52094 & n67947) | (n52094 & n67948) | (n67947 & n67948);
  assign n23342 = ~n67946 & n67949;
  assign n23343 = x139 & x187;
  assign n23344 = n23342 & n23343;
  assign n23345 = n23342 | n23343;
  assign n23346 = ~n23344 & n23345;
  assign n23347 = n67894 & n23346;
  assign n23348 = n67894 | n23346;
  assign n23349 = ~n23347 & n23348;
  assign n23350 = x138 & x188;
  assign n23351 = n23349 & n23350;
  assign n23352 = n23349 | n23350;
  assign n23353 = ~n23351 & n23352;
  assign n52329 = n23058 | n23060;
  assign n52393 = n23353 & n52329;
  assign n52394 = n23058 & n23353;
  assign n52395 = (n67808 & n52393) | (n67808 & n52394) | (n52393 & n52394);
  assign n52396 = n23353 | n52329;
  assign n52397 = n23058 | n23353;
  assign n52398 = (n67808 & n52396) | (n67808 & n52397) | (n52396 & n52397);
  assign n23356 = ~n52395 & n52398;
  assign n23357 = x137 & x189;
  assign n23358 = n23356 & n23357;
  assign n23359 = n23356 | n23357;
  assign n23360 = ~n23358 & n23359;
  assign n52399 = n23065 & n23360;
  assign n67950 = (n23360 & n52271) | (n23360 & n52399) | (n52271 & n52399);
  assign n67951 = (n23360 & n52270) | (n23360 & n52399) | (n52270 & n52399);
  assign n67952 = (n52089 & n67950) | (n52089 & n67951) | (n67950 & n67951);
  assign n52401 = n23065 | n23360;
  assign n67953 = n52271 | n52401;
  assign n67954 = n52270 | n52401;
  assign n67955 = (n52089 & n67953) | (n52089 & n67954) | (n67953 & n67954);
  assign n23363 = ~n67952 & n67955;
  assign n23364 = x136 & x190;
  assign n23365 = n23363 & n23364;
  assign n23366 = n23363 | n23364;
  assign n23367 = ~n23365 & n23366;
  assign n52327 = n23072 | n23074;
  assign n67956 = n23367 & n52327;
  assign n67888 = n22787 | n23072;
  assign n67889 = (n23072 & n23074) | (n23072 & n67888) | (n23074 & n67888);
  assign n67957 = n23367 & n67889;
  assign n67958 = (n67784 & n67956) | (n67784 & n67957) | (n67956 & n67957);
  assign n67959 = n23367 | n52327;
  assign n67960 = n23367 | n67889;
  assign n67961 = (n67784 & n67959) | (n67784 & n67960) | (n67959 & n67960);
  assign n23370 = ~n67958 & n67961;
  assign n23371 = x135 & x191;
  assign n23372 = n23370 & n23371;
  assign n23373 = n23370 | n23371;
  assign n23374 = ~n23372 & n23373;
  assign n52403 = n23079 & n23374;
  assign n67962 = (n23374 & n52280) | (n23374 & n52403) | (n52280 & n52403);
  assign n67963 = (n23081 & n23374) | (n23081 & n52403) | (n23374 & n52403);
  assign n67964 = (n52154 & n67962) | (n52154 & n67963) | (n67962 & n67963);
  assign n52405 = n23079 | n23374;
  assign n67965 = n52280 | n52405;
  assign n67966 = n23081 | n52405;
  assign n67967 = (n52154 & n67965) | (n52154 & n67966) | (n67965 & n67966);
  assign n23377 = ~n67964 & n67967;
  assign n23378 = x134 & x192;
  assign n23379 = n23377 & n23378;
  assign n23380 = n23377 | n23378;
  assign n23381 = ~n23379 & n23380;
  assign n52407 = n23086 & n23381;
  assign n52408 = (n23381 & n52285) | (n23381 & n52407) | (n52285 & n52407);
  assign n52409 = n23086 | n23381;
  assign n52410 = n52285 | n52409;
  assign n23384 = ~n52408 & n52410;
  assign n23385 = x133 & x193;
  assign n23386 = n23384 & n23385;
  assign n23387 = n23384 | n23385;
  assign n23388 = ~n23386 & n23387;
  assign n52411 = n23093 & n23388;
  assign n52412 = (n23388 & n52289) | (n23388 & n52411) | (n52289 & n52411);
  assign n52413 = n23093 | n23388;
  assign n52414 = n52289 | n52413;
  assign n23391 = ~n52412 & n52414;
  assign n23392 = x132 & x194;
  assign n23393 = n23391 & n23392;
  assign n23394 = n23391 | n23392;
  assign n23395 = ~n23393 & n23394;
  assign n52415 = n23100 & n23395;
  assign n52416 = (n23395 & n52293) | (n23395 & n52415) | (n52293 & n52415);
  assign n52417 = n23100 | n23395;
  assign n52418 = n52293 | n52417;
  assign n23398 = ~n52416 & n52418;
  assign n23399 = x131 & x195;
  assign n23400 = n23398 & n23399;
  assign n23401 = n23398 | n23399;
  assign n23402 = ~n23400 & n23401;
  assign n52419 = n23107 & n23402;
  assign n52420 = (n23402 & n52297) | (n23402 & n52419) | (n52297 & n52419);
  assign n52421 = n23107 | n23402;
  assign n52422 = n52297 | n52421;
  assign n23405 = ~n52420 & n52422;
  assign n23406 = x130 & x196;
  assign n23407 = n23405 & n23406;
  assign n23408 = n23405 | n23406;
  assign n23409 = ~n23407 & n23408;
  assign n52423 = n23114 & n23409;
  assign n52424 = (n23409 & n52302) | (n23409 & n52423) | (n52302 & n52423);
  assign n52425 = n23114 | n23409;
  assign n52426 = n52302 | n52425;
  assign n23412 = ~n52424 & n52426;
  assign n23413 = x129 & x197;
  assign n23414 = n23412 & n23413;
  assign n23415 = n23412 | n23413;
  assign n23416 = ~n23414 & n23415;
  assign n52324 = n23121 | n23123;
  assign n52427 = n23416 & n52324;
  assign n52428 = n23121 & n23416;
  assign n52429 = (n52190 & n52427) | (n52190 & n52428) | (n52427 & n52428);
  assign n52430 = n23416 | n52324;
  assign n52431 = n23121 | n23416;
  assign n52432 = (n52190 & n52430) | (n52190 & n52431) | (n52430 & n52431);
  assign n23419 = ~n52429 & n52432;
  assign n23420 = x128 & x198;
  assign n23421 = n23419 & n23420;
  assign n23422 = n23419 | n23420;
  assign n23423 = ~n23421 & n23422;
  assign n52322 = n23128 | n23130;
  assign n67968 = n23423 & n52322;
  assign n67969 = n23128 & n23423;
  assign n67970 = (n52188 & n67968) | (n52188 & n67969) | (n67968 & n67969);
  assign n67971 = n23423 | n52322;
  assign n67972 = n23128 | n23423;
  assign n67973 = (n52188 & n67971) | (n52188 & n67972) | (n67971 & n67972);
  assign n23426 = ~n67970 & n67973;
  assign n23427 = x127 & x199;
  assign n23428 = n23426 & n23427;
  assign n23429 = n23426 | n23427;
  assign n23430 = ~n23428 & n23429;
  assign n52320 = n23135 | n23137;
  assign n67974 = n23430 & n52320;
  assign n67975 = n23135 & n23430;
  assign n67976 = (n52186 & n67974) | (n52186 & n67975) | (n67974 & n67975);
  assign n67977 = n23430 | n52320;
  assign n67978 = n23135 | n23430;
  assign n67979 = (n52186 & n67977) | (n52186 & n67978) | (n67977 & n67978);
  assign n23433 = ~n67976 & n67979;
  assign n23434 = x126 & x200;
  assign n23435 = n23433 & n23434;
  assign n23436 = n23433 | n23434;
  assign n23437 = ~n23435 & n23436;
  assign n23438 = n52319 & n23437;
  assign n23439 = n52319 | n23437;
  assign n23440 = ~n23438 & n23439;
  assign n23441 = x125 & x201;
  assign n23442 = n23440 & n23441;
  assign n23443 = n23440 | n23441;
  assign n23444 = ~n23442 & n23443;
  assign n23445 = n52317 & n23444;
  assign n23446 = n52317 | n23444;
  assign n23447 = ~n23445 & n23446;
  assign n23448 = x124 & x202;
  assign n23449 = n23447 & n23448;
  assign n23450 = n23447 | n23448;
  assign n23451 = ~n23449 & n23450;
  assign n23452 = n52315 & n23451;
  assign n23453 = n52315 | n23451;
  assign n23454 = ~n23452 & n23453;
  assign n23455 = x123 & x203;
  assign n23456 = n23454 & n23455;
  assign n23457 = n23454 | n23455;
  assign n23458 = ~n23456 & n23457;
  assign n23459 = n52313 & n23458;
  assign n23460 = n52313 | n23458;
  assign n23461 = ~n23459 & n23460;
  assign n23462 = x122 & x204;
  assign n23463 = n23461 & n23462;
  assign n23464 = n23461 | n23462;
  assign n23465 = ~n23463 & n23464;
  assign n23466 = n52311 & n23465;
  assign n23467 = n52311 | n23465;
  assign n23468 = ~n23466 & n23467;
  assign n23469 = x121 & x205;
  assign n23470 = n23468 & n23469;
  assign n23471 = n23468 | n23469;
  assign n23472 = ~n23470 & n23471;
  assign n23473 = n23243 & n23472;
  assign n23474 = n23243 | n23472;
  assign n23475 = ~n23473 & n23474;
  assign n23476 = x120 & x206;
  assign n23477 = n23475 & n23476;
  assign n23478 = n23475 | n23476;
  assign n23479 = ~n23477 & n23478;
  assign n23480 = n23242 & n23479;
  assign n23481 = n23242 | n23479;
  assign n23482 = ~n23480 & n23481;
  assign n23483 = x119 & x207;
  assign n23484 = n23482 & n23483;
  assign n23485 = n23482 | n23483;
  assign n23486 = ~n23484 & n23485;
  assign n23487 = n23241 & n23486;
  assign n23488 = n23241 | n23486;
  assign n23489 = ~n23487 & n23488;
  assign n23490 = x118 & x208;
  assign n23491 = n23489 & n23490;
  assign n23492 = n23489 | n23490;
  assign n23493 = ~n23491 & n23492;
  assign n23494 = n23240 & n23493;
  assign n23495 = n23240 | n23493;
  assign n23496 = ~n23494 & n23495;
  assign n23497 = x117 & x209;
  assign n23498 = n23496 & n23497;
  assign n23499 = n23496 | n23497;
  assign n23500 = ~n23498 & n23499;
  assign n23501 = n23239 & n23500;
  assign n23502 = n23239 | n23500;
  assign n23503 = ~n23501 & n23502;
  assign n23504 = x116 & x210;
  assign n23505 = n23503 & n23504;
  assign n23506 = n23503 | n23504;
  assign n23507 = ~n23505 & n23506;
  assign n23508 = n67887 & n23507;
  assign n23509 = n67887 | n23507;
  assign n23510 = ~n23508 & n23509;
  assign n23511 = x115 & x211;
  assign n23512 = n23510 & n23511;
  assign n23513 = n23510 | n23511;
  assign n23514 = ~n23512 & n23513;
  assign n23515 = n52309 & n23514;
  assign n23516 = n52309 | n23514;
  assign n23517 = ~n23515 & n23516;
  assign n23518 = x114 & x212;
  assign n23519 = n23517 & n23518;
  assign n23520 = n23517 | n23518;
  assign n23521 = ~n23519 & n23520;
  assign n23522 = n52307 & n23521;
  assign n23523 = n52307 | n23521;
  assign n23524 = ~n23522 & n23523;
  assign n23525 = x113 & x213;
  assign n23526 = n23524 & n23525;
  assign n23527 = n23524 | n23525;
  assign n23528 = ~n23526 & n23527;
  assign n23529 = n23233 & n23528;
  assign n23530 = n23233 | n23528;
  assign n23531 = ~n23529 & n23530;
  assign n23532 = x112 & x214;
  assign n23533 = n23531 & n23532;
  assign n23534 = n23531 | n23532;
  assign n23535 = ~n23533 & n23534;
  assign n67980 = n23233 | n23525;
  assign n67981 = (n23233 & n23524) | (n23233 & n67980) | (n23524 & n67980);
  assign n52434 = (n23526 & n23528) | (n23526 & n67981) | (n23528 & n67981);
  assign n52435 = n23519 | n52307;
  assign n52436 = (n23519 & n23521) | (n23519 & n52435) | (n23521 & n52435);
  assign n52437 = n23512 | n52309;
  assign n52438 = (n23512 & n23514) | (n23512 & n52437) | (n23514 & n52437);
  assign n67982 = n23505 | n67887;
  assign n67983 = (n23505 & n23507) | (n23505 & n67982) | (n23507 & n67982);
  assign n23540 = n23498 | n23501;
  assign n23541 = n23491 | n23494;
  assign n23542 = n23484 | n23487;
  assign n23543 = n23477 | n23480;
  assign n52439 = n23470 | n23472;
  assign n52440 = (n23243 & n23470) | (n23243 & n52439) | (n23470 & n52439);
  assign n52441 = n23463 | n23465;
  assign n52442 = (n23463 & n52311) | (n23463 & n52441) | (n52311 & n52441);
  assign n52443 = n23456 | n23458;
  assign n52444 = (n23456 & n52313) | (n23456 & n52443) | (n52313 & n52443);
  assign n52445 = n23449 | n23451;
  assign n52446 = (n23449 & n52315) | (n23449 & n52445) | (n52315 & n52445);
  assign n52447 = n23442 | n23444;
  assign n52448 = (n23442 & n52317) | (n23442 & n52447) | (n52317 & n52447);
  assign n52321 = (n23135 & n52186) | (n23135 & n52320) | (n52186 & n52320);
  assign n52323 = (n23128 & n52188) | (n23128 & n52322) | (n52188 & n52322);
  assign n52328 = (n67784 & n67889) | (n67784 & n52327) | (n67889 & n52327);
  assign n52458 = n23358 | n23360;
  assign n67984 = n23065 | n23358;
  assign n67985 = (n23358 & n23360) | (n23358 & n67984) | (n23360 & n67984);
  assign n67986 = (n52271 & n52458) | (n52271 & n67985) | (n52458 & n67985);
  assign n67987 = (n52270 & n52458) | (n52270 & n67985) | (n52458 & n67985);
  assign n67988 = (n52089 & n67986) | (n52089 & n67987) | (n67986 & n67987);
  assign n52463 = n23337 | n23339;
  assign n67989 = n23044 | n23337;
  assign n67990 = (n23337 & n23339) | (n23337 & n67989) | (n23339 & n67989);
  assign n67991 = (n52260 & n52463) | (n52260 & n67990) | (n52463 & n67990);
  assign n67992 = (n52261 & n52463) | (n52261 & n67990) | (n52463 & n67990);
  assign n67993 = (n52094 & n67991) | (n52094 & n67992) | (n67991 & n67992);
  assign n23573 = x151 & x176;
  assign n23574 = x150 & x177;
  assign n23575 = n23573 & n23574;
  assign n23576 = n23573 | n23574;
  assign n23577 = ~n23575 & n23576;
  assign n67996 = n23274 | n23276;
  assign n67998 = n23577 & n67996;
  assign n67999 = n23274 & n23577;
  assign n68000 = (n67916 & n67998) | (n67916 & n67999) | (n67998 & n67999);
  assign n68002 = (n67917 & n67998) | (n67917 & n67999) | (n67998 & n67999);
  assign n68003 = (n67658 & n68000) | (n67658 & n68002) | (n68000 & n68002);
  assign n68004 = (n67657 & n68000) | (n67657 & n68002) | (n68000 & n68002);
  assign n68005 = (n66988 & n68003) | (n66988 & n68004) | (n68003 & n68004);
  assign n68006 = n23577 | n67996;
  assign n68007 = n23274 | n23577;
  assign n68008 = (n67916 & n68006) | (n67916 & n68007) | (n68006 & n68007);
  assign n68009 = (n67917 & n68006) | (n67917 & n68007) | (n68006 & n68007);
  assign n68010 = (n67658 & n68008) | (n67658 & n68009) | (n68008 & n68009);
  assign n68011 = (n67657 & n68008) | (n67657 & n68009) | (n68008 & n68009);
  assign n68012 = (n66988 & n68010) | (n66988 & n68011) | (n68010 & n68011);
  assign n23580 = ~n68005 & n68012;
  assign n23581 = x149 & x178;
  assign n23582 = n23580 & n23581;
  assign n23583 = n23580 | n23581;
  assign n23584 = ~n23582 & n23583;
  assign n68013 = n23281 | n23283;
  assign n68018 = (n23281 & n67927) | (n23281 & n68013) | (n67927 & n68013);
  assign n52489 = n23584 & n68018;
  assign n68015 = n23584 & n68013;
  assign n68016 = n23281 & n23584;
  assign n68017 = (n67925 & n68015) | (n67925 & n68016) | (n68015 & n68016);
  assign n68019 = (n52489 & n67727) | (n52489 & n68017) | (n67727 & n68017);
  assign n68020 = (n52489 & n67726) | (n52489 & n68017) | (n67726 & n68017);
  assign n68021 = (n67426 & n68019) | (n67426 & n68020) | (n68019 & n68020);
  assign n52492 = n23584 | n68018;
  assign n68022 = n23584 | n68013;
  assign n68023 = n23281 | n23584;
  assign n68024 = (n67925 & n68022) | (n67925 & n68023) | (n68022 & n68023);
  assign n68025 = (n52492 & n67727) | (n52492 & n68024) | (n67727 & n68024);
  assign n68026 = (n52492 & n67726) | (n52492 & n68024) | (n67726 & n68024);
  assign n68027 = (n67426 & n68025) | (n67426 & n68026) | (n68025 & n68026);
  assign n23587 = ~n68021 & n68027;
  assign n23588 = x148 & x179;
  assign n23589 = n23587 & n23588;
  assign n23590 = n23587 | n23588;
  assign n23591 = ~n23589 & n23590;
  assign n52474 = n23288 | n23290;
  assign n52494 = n23591 & n52474;
  assign n52495 = n23288 & n23591;
  assign n52496 = (n67914 & n52494) | (n67914 & n52495) | (n52494 & n52495);
  assign n52497 = n23591 | n52474;
  assign n52498 = n23288 | n23591;
  assign n52499 = (n67914 & n52497) | (n67914 & n52498) | (n52497 & n52498);
  assign n23594 = ~n52496 & n52499;
  assign n23595 = x147 & x180;
  assign n23596 = n23594 & n23595;
  assign n23597 = n23594 | n23595;
  assign n23598 = ~n23596 & n23597;
  assign n52500 = n23295 & n23598;
  assign n52501 = (n23598 & n67940) | (n23598 & n52500) | (n67940 & n52500);
  assign n52502 = n23295 | n23598;
  assign n52503 = n67940 | n52502;
  assign n23601 = ~n52501 & n52503;
  assign n23602 = x146 & x181;
  assign n23603 = n23601 & n23602;
  assign n23604 = n23601 | n23602;
  assign n23605 = ~n23603 & n23604;
  assign n52472 = n23302 | n23304;
  assign n52504 = n23605 & n52472;
  assign n52505 = n23302 & n23605;
  assign n52506 = (n67908 & n52504) | (n67908 & n52505) | (n52504 & n52505);
  assign n52507 = n23605 | n52472;
  assign n52508 = n23302 | n23605;
  assign n52509 = (n67908 & n52507) | (n67908 & n52508) | (n52507 & n52508);
  assign n23608 = ~n52506 & n52509;
  assign n23609 = x145 & x182;
  assign n23610 = n23608 & n23609;
  assign n23611 = n23608 | n23609;
  assign n23612 = ~n23610 & n23611;
  assign n52470 = n23309 | n52377;
  assign n68028 = n23612 & n52470;
  assign n67994 = n23016 | n23309;
  assign n67995 = (n23309 & n23311) | (n23309 & n67994) | (n23311 & n67994);
  assign n68029 = n23612 & n67995;
  assign n68030 = (n67817 & n68028) | (n67817 & n68029) | (n68028 & n68029);
  assign n68031 = n23612 | n52470;
  assign n68032 = n23612 | n67995;
  assign n68033 = (n67817 & n68031) | (n67817 & n68032) | (n68031 & n68032);
  assign n23615 = ~n68030 & n68033;
  assign n23616 = x144 & x183;
  assign n23617 = n23615 & n23616;
  assign n23618 = n23615 | n23616;
  assign n23619 = ~n23617 & n23618;
  assign n52467 = n23316 | n23318;
  assign n52510 = n23619 & n52467;
  assign n52511 = n23316 & n23619;
  assign n52512 = (n52341 & n52510) | (n52341 & n52511) | (n52510 & n52511);
  assign n52513 = n23619 | n52467;
  assign n52514 = n23316 | n23619;
  assign n52515 = (n52341 & n52513) | (n52341 & n52514) | (n52513 & n52514);
  assign n23622 = ~n52512 & n52515;
  assign n23623 = x143 & x184;
  assign n23624 = n23622 & n23623;
  assign n23625 = n23622 | n23623;
  assign n23626 = ~n23624 & n23625;
  assign n52465 = n23323 | n23325;
  assign n52516 = n23626 & n52465;
  assign n52517 = n23323 & n23626;
  assign n52518 = (n67899 & n52516) | (n67899 & n52517) | (n52516 & n52517);
  assign n52519 = n23626 | n52465;
  assign n52520 = n23323 | n23626;
  assign n52521 = (n67899 & n52519) | (n67899 & n52520) | (n52519 & n52520);
  assign n23629 = ~n52518 & n52521;
  assign n23630 = x142 & x185;
  assign n23631 = n23629 & n23630;
  assign n23632 = n23629 | n23630;
  assign n23633 = ~n23631 & n23632;
  assign n52522 = n23330 & n23633;
  assign n68034 = (n23633 & n52384) | (n23633 & n52522) | (n52384 & n52522);
  assign n68035 = (n23633 & n52383) | (n23633 & n52522) | (n52383 & n52522);
  assign n68036 = (n52202 & n68034) | (n52202 & n68035) | (n68034 & n68035);
  assign n52524 = n23330 | n23633;
  assign n68037 = n52384 | n52524;
  assign n68038 = n52383 | n52524;
  assign n68039 = (n52202 & n68037) | (n52202 & n68038) | (n68037 & n68038);
  assign n23636 = ~n68036 & n68039;
  assign n23637 = x141 & x186;
  assign n23638 = n23636 & n23637;
  assign n23639 = n23636 | n23637;
  assign n23640 = ~n23638 & n23639;
  assign n23641 = n67993 & n23640;
  assign n23642 = n67993 | n23640;
  assign n23643 = ~n23641 & n23642;
  assign n23644 = x140 & x187;
  assign n23645 = n23643 & n23644;
  assign n23646 = n23643 | n23644;
  assign n23647 = ~n23645 & n23646;
  assign n52460 = n23344 | n23346;
  assign n52526 = n23647 & n52460;
  assign n52527 = n23344 & n23647;
  assign n52528 = (n67894 & n52526) | (n67894 & n52527) | (n52526 & n52527);
  assign n52529 = n23647 | n52460;
  assign n52530 = n23344 | n23647;
  assign n52531 = (n67894 & n52529) | (n67894 & n52530) | (n52529 & n52530);
  assign n23650 = ~n52528 & n52531;
  assign n23651 = x139 & x188;
  assign n23652 = n23650 & n23651;
  assign n23653 = n23650 | n23651;
  assign n23654 = ~n23652 & n23653;
  assign n52532 = n23351 & n23654;
  assign n68040 = (n23654 & n52394) | (n23654 & n52532) | (n52394 & n52532);
  assign n68041 = (n23654 & n52393) | (n23654 & n52532) | (n52393 & n52532);
  assign n68042 = (n67808 & n68040) | (n67808 & n68041) | (n68040 & n68041);
  assign n52534 = n23351 | n23654;
  assign n68043 = n52394 | n52534;
  assign n68044 = n52393 | n52534;
  assign n68045 = (n67808 & n68043) | (n67808 & n68044) | (n68043 & n68044);
  assign n23657 = ~n68042 & n68045;
  assign n23658 = x138 & x189;
  assign n23659 = n23657 & n23658;
  assign n23660 = n23657 | n23658;
  assign n23661 = ~n23659 & n23660;
  assign n23662 = n67988 & n23661;
  assign n23663 = n67988 | n23661;
  assign n23664 = ~n23662 & n23663;
  assign n23665 = x137 & x190;
  assign n23666 = n23664 & n23665;
  assign n23667 = n23664 | n23665;
  assign n23668 = ~n23666 & n23667;
  assign n52455 = n23365 | n23367;
  assign n52536 = n23668 & n52455;
  assign n52537 = n23365 & n23668;
  assign n52538 = (n52328 & n52536) | (n52328 & n52537) | (n52536 & n52537);
  assign n52539 = n23668 | n52455;
  assign n52540 = n23365 | n23668;
  assign n52541 = (n52328 & n52539) | (n52328 & n52540) | (n52539 & n52540);
  assign n23671 = ~n52538 & n52541;
  assign n23672 = x136 & x191;
  assign n23673 = n23671 & n23672;
  assign n23674 = n23671 | n23672;
  assign n23675 = ~n23673 & n23674;
  assign n52542 = n23372 & n23675;
  assign n52543 = (n23675 & n67964) | (n23675 & n52542) | (n67964 & n52542);
  assign n52544 = n23372 | n23675;
  assign n52545 = n67964 | n52544;
  assign n23678 = ~n52543 & n52545;
  assign n23679 = x135 & x192;
  assign n23680 = n23678 & n23679;
  assign n23681 = n23678 | n23679;
  assign n23682 = ~n23680 & n23681;
  assign n52546 = n23379 & n23682;
  assign n52547 = (n23682 & n52408) | (n23682 & n52546) | (n52408 & n52546);
  assign n52548 = n23379 | n23682;
  assign n52549 = n52408 | n52548;
  assign n23685 = ~n52547 & n52549;
  assign n23686 = x134 & x193;
  assign n23687 = n23685 & n23686;
  assign n23688 = n23685 | n23686;
  assign n23689 = ~n23687 & n23688;
  assign n52550 = n23386 & n23689;
  assign n52551 = (n23689 & n52412) | (n23689 & n52550) | (n52412 & n52550);
  assign n52552 = n23386 | n23689;
  assign n52553 = n52412 | n52552;
  assign n23692 = ~n52551 & n52553;
  assign n23693 = x133 & x194;
  assign n23694 = n23692 & n23693;
  assign n23695 = n23692 | n23693;
  assign n23696 = ~n23694 & n23695;
  assign n52554 = n23393 & n23696;
  assign n52555 = (n23696 & n52416) | (n23696 & n52554) | (n52416 & n52554);
  assign n52556 = n23393 | n23696;
  assign n52557 = n52416 | n52556;
  assign n23699 = ~n52555 & n52557;
  assign n23700 = x132 & x195;
  assign n23701 = n23699 & n23700;
  assign n23702 = n23699 | n23700;
  assign n23703 = ~n23701 & n23702;
  assign n52558 = n23400 & n23703;
  assign n52559 = (n23703 & n52420) | (n23703 & n52558) | (n52420 & n52558);
  assign n52560 = n23400 | n23703;
  assign n52561 = n52420 | n52560;
  assign n23706 = ~n52559 & n52561;
  assign n23707 = x131 & x196;
  assign n23708 = n23706 & n23707;
  assign n23709 = n23706 | n23707;
  assign n23710 = ~n23708 & n23709;
  assign n52562 = n23407 & n23710;
  assign n52563 = (n23710 & n52424) | (n23710 & n52562) | (n52424 & n52562);
  assign n52564 = n23407 | n23710;
  assign n52565 = n52424 | n52564;
  assign n23713 = ~n52563 & n52565;
  assign n23714 = x130 & x197;
  assign n23715 = n23713 & n23714;
  assign n23716 = n23713 | n23714;
  assign n23717 = ~n23715 & n23716;
  assign n52566 = n23414 & n23717;
  assign n52567 = (n23717 & n52429) | (n23717 & n52566) | (n52429 & n52566);
  assign n52568 = n23414 | n23717;
  assign n52569 = n52429 | n52568;
  assign n23720 = ~n52567 & n52569;
  assign n23721 = x129 & x198;
  assign n23722 = n23720 & n23721;
  assign n23723 = n23720 | n23721;
  assign n23724 = ~n23722 & n23723;
  assign n52453 = n23421 | n23423;
  assign n52570 = n23724 & n52453;
  assign n52571 = n23421 & n23724;
  assign n52572 = (n52323 & n52570) | (n52323 & n52571) | (n52570 & n52571);
  assign n52573 = n23724 | n52453;
  assign n52574 = n23421 | n23724;
  assign n52575 = (n52323 & n52573) | (n52323 & n52574) | (n52573 & n52574);
  assign n23727 = ~n52572 & n52575;
  assign n23728 = x128 & x199;
  assign n23729 = n23727 & n23728;
  assign n23730 = n23727 | n23728;
  assign n23731 = ~n23729 & n23730;
  assign n52451 = n23428 | n23430;
  assign n68046 = n23731 & n52451;
  assign n68047 = n23428 & n23731;
  assign n68048 = (n52321 & n68046) | (n52321 & n68047) | (n68046 & n68047);
  assign n68049 = n23731 | n52451;
  assign n68050 = n23428 | n23731;
  assign n68051 = (n52321 & n68049) | (n52321 & n68050) | (n68049 & n68050);
  assign n23734 = ~n68048 & n68051;
  assign n23735 = x127 & x200;
  assign n23736 = n23734 & n23735;
  assign n23737 = n23734 | n23735;
  assign n23738 = ~n23736 & n23737;
  assign n52449 = n23435 | n23437;
  assign n68052 = n23738 & n52449;
  assign n68053 = n23435 & n23738;
  assign n68054 = (n52319 & n68052) | (n52319 & n68053) | (n68052 & n68053);
  assign n68055 = n23738 | n52449;
  assign n68056 = n23435 | n23738;
  assign n68057 = (n52319 & n68055) | (n52319 & n68056) | (n68055 & n68056);
  assign n23741 = ~n68054 & n68057;
  assign n23742 = x126 & x201;
  assign n23743 = n23741 & n23742;
  assign n23744 = n23741 | n23742;
  assign n23745 = ~n23743 & n23744;
  assign n23746 = n52448 & n23745;
  assign n23747 = n52448 | n23745;
  assign n23748 = ~n23746 & n23747;
  assign n23749 = x125 & x202;
  assign n23750 = n23748 & n23749;
  assign n23751 = n23748 | n23749;
  assign n23752 = ~n23750 & n23751;
  assign n23753 = n52446 & n23752;
  assign n23754 = n52446 | n23752;
  assign n23755 = ~n23753 & n23754;
  assign n23756 = x124 & x203;
  assign n23757 = n23755 & n23756;
  assign n23758 = n23755 | n23756;
  assign n23759 = ~n23757 & n23758;
  assign n23760 = n52444 & n23759;
  assign n23761 = n52444 | n23759;
  assign n23762 = ~n23760 & n23761;
  assign n23763 = x123 & x204;
  assign n23764 = n23762 & n23763;
  assign n23765 = n23762 | n23763;
  assign n23766 = ~n23764 & n23765;
  assign n23767 = n52442 & n23766;
  assign n23768 = n52442 | n23766;
  assign n23769 = ~n23767 & n23768;
  assign n23770 = x122 & x205;
  assign n23771 = n23769 & n23770;
  assign n23772 = n23769 | n23770;
  assign n23773 = ~n23771 & n23772;
  assign n23774 = n52440 & n23773;
  assign n23775 = n52440 | n23773;
  assign n23776 = ~n23774 & n23775;
  assign n23777 = x121 & x206;
  assign n23778 = n23776 & n23777;
  assign n23779 = n23776 | n23777;
  assign n23780 = ~n23778 & n23779;
  assign n23781 = n23543 & n23780;
  assign n23782 = n23543 | n23780;
  assign n23783 = ~n23781 & n23782;
  assign n23784 = x120 & x207;
  assign n23785 = n23783 & n23784;
  assign n23786 = n23783 | n23784;
  assign n23787 = ~n23785 & n23786;
  assign n23788 = n23542 & n23787;
  assign n23789 = n23542 | n23787;
  assign n23790 = ~n23788 & n23789;
  assign n23791 = x119 & x208;
  assign n23792 = n23790 & n23791;
  assign n23793 = n23790 | n23791;
  assign n23794 = ~n23792 & n23793;
  assign n23795 = n23541 & n23794;
  assign n23796 = n23541 | n23794;
  assign n23797 = ~n23795 & n23796;
  assign n23798 = x118 & x209;
  assign n23799 = n23797 & n23798;
  assign n23800 = n23797 | n23798;
  assign n23801 = ~n23799 & n23800;
  assign n23802 = n23540 & n23801;
  assign n23803 = n23540 | n23801;
  assign n23804 = ~n23802 & n23803;
  assign n23805 = x117 & x210;
  assign n23806 = n23804 & n23805;
  assign n23807 = n23804 | n23805;
  assign n23808 = ~n23806 & n23807;
  assign n23809 = n67983 & n23808;
  assign n23810 = n67983 | n23808;
  assign n23811 = ~n23809 & n23810;
  assign n23812 = x116 & x211;
  assign n23813 = n23811 & n23812;
  assign n23814 = n23811 | n23812;
  assign n23815 = ~n23813 & n23814;
  assign n23816 = n52438 & n23815;
  assign n23817 = n52438 | n23815;
  assign n23818 = ~n23816 & n23817;
  assign n23819 = x115 & x212;
  assign n23820 = n23818 & n23819;
  assign n23821 = n23818 | n23819;
  assign n23822 = ~n23820 & n23821;
  assign n23823 = n52436 & n23822;
  assign n23824 = n52436 | n23822;
  assign n23825 = ~n23823 & n23824;
  assign n23826 = x114 & x213;
  assign n23827 = n23825 & n23826;
  assign n23828 = n23825 | n23826;
  assign n23829 = ~n23827 & n23828;
  assign n23830 = n52434 & n23829;
  assign n23831 = n52434 | n23829;
  assign n23832 = ~n23830 & n23831;
  assign n23833 = x113 & x214;
  assign n23834 = n23832 & n23833;
  assign n23835 = n23832 | n23833;
  assign n23836 = ~n23834 & n23835;
  assign n23837 = n23533 & n23836;
  assign n23838 = n23533 | n23836;
  assign n23839 = ~n23837 & n23838;
  assign n23840 = x112 & x215;
  assign n23841 = n23839 & n23840;
  assign n23842 = n23839 | n23840;
  assign n23843 = ~n23841 & n23842;
  assign n68058 = n23533 | n23833;
  assign n68059 = (n23533 & n23832) | (n23533 & n68058) | (n23832 & n68058);
  assign n52577 = (n23834 & n23836) | (n23834 & n68059) | (n23836 & n68059);
  assign n52578 = n23827 | n52434;
  assign n52579 = (n23827 & n23829) | (n23827 & n52578) | (n23829 & n52578);
  assign n52580 = n23820 | n52436;
  assign n52581 = (n23820 & n23822) | (n23820 & n52580) | (n23822 & n52580);
  assign n52582 = n23813 | n52438;
  assign n52583 = (n23813 & n23815) | (n23813 & n52582) | (n23815 & n52582);
  assign n68060 = n23806 | n67983;
  assign n68061 = (n23806 & n23808) | (n23806 & n68060) | (n23808 & n68060);
  assign n23849 = n23799 | n23802;
  assign n23850 = n23792 | n23795;
  assign n23851 = n23785 | n23788;
  assign n52584 = n23778 | n23780;
  assign n52585 = (n23543 & n23778) | (n23543 & n52584) | (n23778 & n52584);
  assign n52586 = n23771 | n23773;
  assign n52587 = (n23771 & n52440) | (n23771 & n52586) | (n52440 & n52586);
  assign n52588 = n23764 | n23766;
  assign n52589 = (n23764 & n52442) | (n23764 & n52588) | (n52442 & n52588);
  assign n52590 = n23757 | n23759;
  assign n52591 = (n23757 & n52444) | (n23757 & n52590) | (n52444 & n52590);
  assign n52592 = n23750 | n23752;
  assign n52593 = (n23750 & n52446) | (n23750 & n52592) | (n52446 & n52592);
  assign n52450 = (n23435 & n52319) | (n23435 & n52449) | (n52319 & n52449);
  assign n52452 = (n23428 & n52321) | (n23428 & n52451) | (n52321 & n52451);
  assign n52606 = n23652 | n23654;
  assign n68064 = n23351 | n23652;
  assign n68065 = (n23652 & n23654) | (n23652 & n68064) | (n23654 & n68064);
  assign n68066 = (n52394 & n52606) | (n52394 & n68065) | (n52606 & n68065);
  assign n68067 = (n52393 & n52606) | (n52393 & n68065) | (n52606 & n68065);
  assign n68068 = (n67808 & n68066) | (n67808 & n68067) | (n68066 & n68067);
  assign n52611 = n23631 | n23633;
  assign n68069 = n23330 | n23631;
  assign n68070 = (n23631 & n23633) | (n23631 & n68069) | (n23633 & n68069);
  assign n68071 = (n52384 & n52611) | (n52384 & n68070) | (n52611 & n68070);
  assign n68072 = (n52383 & n52611) | (n52383 & n68070) | (n52611 & n68070);
  assign n68073 = (n52202 & n68071) | (n52202 & n68072) | (n68071 & n68072);
  assign n23882 = x152 & x176;
  assign n23883 = x151 & x177;
  assign n23884 = n23882 & n23883;
  assign n23885 = n23882 | n23883;
  assign n23886 = ~n23884 & n23885;
  assign n68078 = n23575 & n23886;
  assign n68079 = (n23886 & n68000) | (n23886 & n68078) | (n68000 & n68078);
  assign n68080 = (n23886 & n68002) | (n23886 & n68078) | (n68002 & n68078);
  assign n68081 = (n67658 & n68079) | (n67658 & n68080) | (n68079 & n68080);
  assign n68082 = (n67657 & n68079) | (n67657 & n68080) | (n68079 & n68080);
  assign n68083 = (n66988 & n68081) | (n66988 & n68082) | (n68081 & n68082);
  assign n68084 = n23575 | n23886;
  assign n68085 = n68000 | n68084;
  assign n68086 = n68002 | n68084;
  assign n68087 = (n67658 & n68085) | (n67658 & n68086) | (n68085 & n68086);
  assign n68088 = (n67657 & n68085) | (n67657 & n68086) | (n68085 & n68086);
  assign n68089 = (n66988 & n68087) | (n66988 & n68088) | (n68087 & n68088);
  assign n23889 = ~n68083 & n68089;
  assign n23890 = x150 & x178;
  assign n23891 = n23889 & n23890;
  assign n23892 = n23889 | n23890;
  assign n23893 = ~n23891 & n23892;
  assign n52636 = n23582 & n23893;
  assign n68090 = (n23893 & n52636) | (n23893 & n68020) | (n52636 & n68020);
  assign n68091 = (n23893 & n52636) | (n23893 & n68019) | (n52636 & n68019);
  assign n68092 = (n67426 & n68090) | (n67426 & n68091) | (n68090 & n68091);
  assign n52638 = n23582 | n23893;
  assign n68093 = n52638 | n68020;
  assign n68094 = n52638 | n68019;
  assign n68095 = (n67426 & n68093) | (n67426 & n68094) | (n68093 & n68094);
  assign n23896 = ~n68092 & n68095;
  assign n23897 = x149 & x179;
  assign n23898 = n23896 & n23897;
  assign n23899 = n23896 | n23897;
  assign n23900 = ~n23898 & n23899;
  assign n68096 = n23589 | n23591;
  assign n68097 = (n23589 & n52474) | (n23589 & n68096) | (n52474 & n68096);
  assign n52640 = n23900 & n68097;
  assign n68098 = n23288 | n23589;
  assign n68099 = (n23589 & n23591) | (n23589 & n68098) | (n23591 & n68098);
  assign n52641 = n23900 & n68099;
  assign n52642 = (n67914 & n52640) | (n67914 & n52641) | (n52640 & n52641);
  assign n52643 = n23900 | n68097;
  assign n52644 = n23900 | n68099;
  assign n52645 = (n67914 & n52643) | (n67914 & n52644) | (n52643 & n52644);
  assign n23903 = ~n52642 & n52645;
  assign n23904 = x148 & x180;
  assign n23905 = n23903 & n23904;
  assign n23906 = n23903 | n23904;
  assign n23907 = ~n23905 & n23906;
  assign n68100 = n23295 | n23596;
  assign n68101 = (n23596 & n23598) | (n23596 & n68100) | (n23598 & n68100);
  assign n52646 = n23907 & n68101;
  assign n52622 = n23596 | n23598;
  assign n52647 = n23907 & n52622;
  assign n52648 = (n67940 & n52646) | (n67940 & n52647) | (n52646 & n52647);
  assign n52649 = n23907 | n68101;
  assign n52650 = n23907 | n52622;
  assign n52651 = (n67940 & n52649) | (n67940 & n52650) | (n52649 & n52650);
  assign n23910 = ~n52648 & n52651;
  assign n23911 = x147 & x181;
  assign n23912 = n23910 & n23911;
  assign n23913 = n23910 | n23911;
  assign n23914 = ~n23912 & n23913;
  assign n68102 = n23603 & n23914;
  assign n68103 = (n23914 & n52504) | (n23914 & n68102) | (n52504 & n68102);
  assign n68104 = n23302 | n23603;
  assign n68105 = (n23603 & n23605) | (n23603 & n68104) | (n23605 & n68104);
  assign n52653 = n23914 & n68105;
  assign n52654 = (n67908 & n68103) | (n67908 & n52653) | (n68103 & n52653);
  assign n68106 = n23603 | n23914;
  assign n68107 = n52504 | n68106;
  assign n52656 = n23914 | n68105;
  assign n52657 = (n67908 & n68107) | (n67908 & n52656) | (n68107 & n52656);
  assign n23917 = ~n52654 & n52657;
  assign n23918 = x146 & x182;
  assign n23919 = n23917 & n23918;
  assign n23920 = n23917 | n23918;
  assign n23921 = ~n23919 & n23920;
  assign n52616 = n23610 | n23612;
  assign n52658 = n23921 & n52616;
  assign n52659 = n23610 & n23921;
  assign n68108 = (n52470 & n52658) | (n52470 & n52659) | (n52658 & n52659);
  assign n68109 = (n52658 & n52659) | (n52658 & n67995) | (n52659 & n67995);
  assign n68110 = (n67817 & n68108) | (n67817 & n68109) | (n68108 & n68109);
  assign n52661 = n23921 | n52616;
  assign n52662 = n23610 | n23921;
  assign n68111 = (n52470 & n52661) | (n52470 & n52662) | (n52661 & n52662);
  assign n68112 = (n52661 & n52662) | (n52661 & n67995) | (n52662 & n67995);
  assign n68113 = (n67817 & n68111) | (n67817 & n68112) | (n68111 & n68112);
  assign n23924 = ~n68110 & n68113;
  assign n23925 = x145 & x183;
  assign n23926 = n23924 & n23925;
  assign n23927 = n23924 | n23925;
  assign n23928 = ~n23926 & n23927;
  assign n68076 = n23617 | n23619;
  assign n68077 = (n23617 & n52467) | (n23617 & n68076) | (n52467 & n68076);
  assign n68114 = n23928 & n68077;
  assign n68074 = n23316 | n23617;
  assign n68075 = (n23617 & n23619) | (n23617 & n68074) | (n23619 & n68074);
  assign n68115 = n23928 & n68075;
  assign n68116 = (n52341 & n68114) | (n52341 & n68115) | (n68114 & n68115);
  assign n68117 = n23928 | n68077;
  assign n68118 = n23928 | n68075;
  assign n68119 = (n52341 & n68117) | (n52341 & n68118) | (n68117 & n68118);
  assign n23931 = ~n68116 & n68119;
  assign n23932 = x144 & x184;
  assign n23933 = n23931 & n23932;
  assign n23934 = n23931 | n23932;
  assign n23935 = ~n23933 & n23934;
  assign n52664 = n23624 & n23935;
  assign n52665 = (n23935 & n52518) | (n23935 & n52664) | (n52518 & n52664);
  assign n52666 = n23624 | n23935;
  assign n52667 = n52518 | n52666;
  assign n23938 = ~n52665 & n52667;
  assign n23939 = x143 & x185;
  assign n23940 = n23938 & n23939;
  assign n23941 = n23938 | n23939;
  assign n23942 = ~n23940 & n23941;
  assign n23943 = n68073 & n23942;
  assign n23944 = n68073 | n23942;
  assign n23945 = ~n23943 & n23944;
  assign n23946 = x142 & x186;
  assign n23947 = n23945 & n23946;
  assign n23948 = n23945 | n23946;
  assign n23949 = ~n23947 & n23948;
  assign n52608 = n23638 | n23640;
  assign n52668 = n23949 & n52608;
  assign n52669 = n23638 & n23949;
  assign n52670 = (n67993 & n52668) | (n67993 & n52669) | (n52668 & n52669);
  assign n52671 = n23949 | n52608;
  assign n52672 = n23638 | n23949;
  assign n52673 = (n67993 & n52671) | (n67993 & n52672) | (n52671 & n52672);
  assign n23952 = ~n52670 & n52673;
  assign n23953 = x141 & x187;
  assign n23954 = n23952 & n23953;
  assign n23955 = n23952 | n23953;
  assign n23956 = ~n23954 & n23955;
  assign n52674 = n23645 & n23956;
  assign n68120 = (n23956 & n52527) | (n23956 & n52674) | (n52527 & n52674);
  assign n68121 = (n23956 & n52526) | (n23956 & n52674) | (n52526 & n52674);
  assign n68122 = (n67894 & n68120) | (n67894 & n68121) | (n68120 & n68121);
  assign n52676 = n23645 | n23956;
  assign n68123 = n52527 | n52676;
  assign n68124 = n52526 | n52676;
  assign n68125 = (n67894 & n68123) | (n67894 & n68124) | (n68123 & n68124);
  assign n23959 = ~n68122 & n68125;
  assign n23960 = x140 & x188;
  assign n23961 = n23959 & n23960;
  assign n23962 = n23959 | n23960;
  assign n23963 = ~n23961 & n23962;
  assign n23964 = n68068 & n23963;
  assign n23965 = n68068 | n23963;
  assign n23966 = ~n23964 & n23965;
  assign n23967 = x139 & x189;
  assign n23968 = n23966 & n23967;
  assign n23969 = n23966 | n23967;
  assign n23970 = ~n23968 & n23969;
  assign n52603 = n23659 | n23661;
  assign n52678 = n23970 & n52603;
  assign n52679 = n23659 & n23970;
  assign n52680 = (n67988 & n52678) | (n67988 & n52679) | (n52678 & n52679);
  assign n52681 = n23970 | n52603;
  assign n52682 = n23659 | n23970;
  assign n52683 = (n67988 & n52681) | (n67988 & n52682) | (n52681 & n52682);
  assign n23973 = ~n52680 & n52683;
  assign n23974 = x138 & x190;
  assign n23975 = n23973 & n23974;
  assign n23976 = n23973 | n23974;
  assign n23977 = ~n23975 & n23976;
  assign n52684 = n23666 & n23977;
  assign n68126 = (n23977 & n52537) | (n23977 & n52684) | (n52537 & n52684);
  assign n68127 = (n23977 & n52536) | (n23977 & n52684) | (n52536 & n52684);
  assign n68128 = (n52328 & n68126) | (n52328 & n68127) | (n68126 & n68127);
  assign n52686 = n23666 | n23977;
  assign n68129 = n52537 | n52686;
  assign n68130 = n52536 | n52686;
  assign n68131 = (n52328 & n68129) | (n52328 & n68130) | (n68129 & n68130);
  assign n23980 = ~n68128 & n68131;
  assign n23981 = x137 & x191;
  assign n23982 = n23980 & n23981;
  assign n23983 = n23980 | n23981;
  assign n23984 = ~n23982 & n23983;
  assign n52601 = n23673 | n23675;
  assign n68132 = n23984 & n52601;
  assign n68062 = n23372 | n23673;
  assign n68063 = (n23673 & n23675) | (n23673 & n68062) | (n23675 & n68062);
  assign n68133 = n23984 & n68063;
  assign n68134 = (n67964 & n68132) | (n67964 & n68133) | (n68132 & n68133);
  assign n68135 = n23984 | n52601;
  assign n68136 = n23984 | n68063;
  assign n68137 = (n67964 & n68135) | (n67964 & n68136) | (n68135 & n68136);
  assign n23987 = ~n68134 & n68137;
  assign n23988 = x136 & x192;
  assign n23989 = n23987 & n23988;
  assign n23990 = n23987 | n23988;
  assign n23991 = ~n23989 & n23990;
  assign n52688 = n23680 & n23991;
  assign n68138 = (n23991 & n52546) | (n23991 & n52688) | (n52546 & n52688);
  assign n68139 = (n23682 & n23991) | (n23682 & n52688) | (n23991 & n52688);
  assign n68140 = (n52408 & n68138) | (n52408 & n68139) | (n68138 & n68139);
  assign n52690 = n23680 | n23991;
  assign n68141 = n52546 | n52690;
  assign n68142 = n23682 | n52690;
  assign n68143 = (n52408 & n68141) | (n52408 & n68142) | (n68141 & n68142);
  assign n23994 = ~n68140 & n68143;
  assign n23995 = x135 & x193;
  assign n23996 = n23994 & n23995;
  assign n23997 = n23994 | n23995;
  assign n23998 = ~n23996 & n23997;
  assign n52692 = n23687 & n23998;
  assign n52693 = (n23998 & n52551) | (n23998 & n52692) | (n52551 & n52692);
  assign n52694 = n23687 | n23998;
  assign n52695 = n52551 | n52694;
  assign n24001 = ~n52693 & n52695;
  assign n24002 = x134 & x194;
  assign n24003 = n24001 & n24002;
  assign n24004 = n24001 | n24002;
  assign n24005 = ~n24003 & n24004;
  assign n52696 = n23694 & n24005;
  assign n52697 = (n24005 & n52555) | (n24005 & n52696) | (n52555 & n52696);
  assign n52698 = n23694 | n24005;
  assign n52699 = n52555 | n52698;
  assign n24008 = ~n52697 & n52699;
  assign n24009 = x133 & x195;
  assign n24010 = n24008 & n24009;
  assign n24011 = n24008 | n24009;
  assign n24012 = ~n24010 & n24011;
  assign n52700 = n23701 & n24012;
  assign n52701 = (n24012 & n52559) | (n24012 & n52700) | (n52559 & n52700);
  assign n52702 = n23701 | n24012;
  assign n52703 = n52559 | n52702;
  assign n24015 = ~n52701 & n52703;
  assign n24016 = x132 & x196;
  assign n24017 = n24015 & n24016;
  assign n24018 = n24015 | n24016;
  assign n24019 = ~n24017 & n24018;
  assign n52704 = n23708 & n24019;
  assign n52705 = (n24019 & n52563) | (n24019 & n52704) | (n52563 & n52704);
  assign n52706 = n23708 | n24019;
  assign n52707 = n52563 | n52706;
  assign n24022 = ~n52705 & n52707;
  assign n24023 = x131 & x197;
  assign n24024 = n24022 & n24023;
  assign n24025 = n24022 | n24023;
  assign n24026 = ~n24024 & n24025;
  assign n52708 = n23715 & n24026;
  assign n52709 = (n24026 & n52567) | (n24026 & n52708) | (n52567 & n52708);
  assign n52710 = n23715 | n24026;
  assign n52711 = n52567 | n52710;
  assign n24029 = ~n52709 & n52711;
  assign n24030 = x130 & x198;
  assign n24031 = n24029 & n24030;
  assign n24032 = n24029 | n24030;
  assign n24033 = ~n24031 & n24032;
  assign n52712 = n23722 & n24033;
  assign n52713 = (n24033 & n52572) | (n24033 & n52712) | (n52572 & n52712);
  assign n52714 = n23722 | n24033;
  assign n52715 = n52572 | n52714;
  assign n24036 = ~n52713 & n52715;
  assign n24037 = x129 & x199;
  assign n24038 = n24036 & n24037;
  assign n24039 = n24036 | n24037;
  assign n24040 = ~n24038 & n24039;
  assign n52598 = n23729 | n23731;
  assign n52716 = n24040 & n52598;
  assign n52717 = n23729 & n24040;
  assign n52718 = (n52452 & n52716) | (n52452 & n52717) | (n52716 & n52717);
  assign n52719 = n24040 | n52598;
  assign n52720 = n23729 | n24040;
  assign n52721 = (n52452 & n52719) | (n52452 & n52720) | (n52719 & n52720);
  assign n24043 = ~n52718 & n52721;
  assign n24044 = x128 & x200;
  assign n24045 = n24043 & n24044;
  assign n24046 = n24043 | n24044;
  assign n24047 = ~n24045 & n24046;
  assign n52596 = n23736 | n23738;
  assign n68144 = n24047 & n52596;
  assign n68145 = n23736 & n24047;
  assign n68146 = (n52450 & n68144) | (n52450 & n68145) | (n68144 & n68145);
  assign n68147 = n24047 | n52596;
  assign n68148 = n23736 | n24047;
  assign n68149 = (n52450 & n68147) | (n52450 & n68148) | (n68147 & n68148);
  assign n24050 = ~n68146 & n68149;
  assign n24051 = x127 & x201;
  assign n24052 = n24050 & n24051;
  assign n24053 = n24050 | n24051;
  assign n24054 = ~n24052 & n24053;
  assign n52594 = n23743 | n23745;
  assign n68150 = n24054 & n52594;
  assign n68151 = n23743 & n24054;
  assign n68152 = (n52448 & n68150) | (n52448 & n68151) | (n68150 & n68151);
  assign n68153 = n24054 | n52594;
  assign n68154 = n23743 | n24054;
  assign n68155 = (n52448 & n68153) | (n52448 & n68154) | (n68153 & n68154);
  assign n24057 = ~n68152 & n68155;
  assign n24058 = x126 & x202;
  assign n24059 = n24057 & n24058;
  assign n24060 = n24057 | n24058;
  assign n24061 = ~n24059 & n24060;
  assign n24062 = n52593 & n24061;
  assign n24063 = n52593 | n24061;
  assign n24064 = ~n24062 & n24063;
  assign n24065 = x125 & x203;
  assign n24066 = n24064 & n24065;
  assign n24067 = n24064 | n24065;
  assign n24068 = ~n24066 & n24067;
  assign n24069 = n52591 & n24068;
  assign n24070 = n52591 | n24068;
  assign n24071 = ~n24069 & n24070;
  assign n24072 = x124 & x204;
  assign n24073 = n24071 & n24072;
  assign n24074 = n24071 | n24072;
  assign n24075 = ~n24073 & n24074;
  assign n24076 = n52589 & n24075;
  assign n24077 = n52589 | n24075;
  assign n24078 = ~n24076 & n24077;
  assign n24079 = x123 & x205;
  assign n24080 = n24078 & n24079;
  assign n24081 = n24078 | n24079;
  assign n24082 = ~n24080 & n24081;
  assign n24083 = n52587 & n24082;
  assign n24084 = n52587 | n24082;
  assign n24085 = ~n24083 & n24084;
  assign n24086 = x122 & x206;
  assign n24087 = n24085 & n24086;
  assign n24088 = n24085 | n24086;
  assign n24089 = ~n24087 & n24088;
  assign n24090 = n52585 & n24089;
  assign n24091 = n52585 | n24089;
  assign n24092 = ~n24090 & n24091;
  assign n24093 = x121 & x207;
  assign n24094 = n24092 & n24093;
  assign n24095 = n24092 | n24093;
  assign n24096 = ~n24094 & n24095;
  assign n24097 = n23851 & n24096;
  assign n24098 = n23851 | n24096;
  assign n24099 = ~n24097 & n24098;
  assign n24100 = x120 & x208;
  assign n24101 = n24099 & n24100;
  assign n24102 = n24099 | n24100;
  assign n24103 = ~n24101 & n24102;
  assign n24104 = n23850 & n24103;
  assign n24105 = n23850 | n24103;
  assign n24106 = ~n24104 & n24105;
  assign n24107 = x119 & x209;
  assign n24108 = n24106 & n24107;
  assign n24109 = n24106 | n24107;
  assign n24110 = ~n24108 & n24109;
  assign n24111 = n23849 & n24110;
  assign n24112 = n23849 | n24110;
  assign n24113 = ~n24111 & n24112;
  assign n24114 = x118 & x210;
  assign n24115 = n24113 & n24114;
  assign n24116 = n24113 | n24114;
  assign n24117 = ~n24115 & n24116;
  assign n24118 = n68061 & n24117;
  assign n24119 = n68061 | n24117;
  assign n24120 = ~n24118 & n24119;
  assign n24121 = x117 & x211;
  assign n24122 = n24120 & n24121;
  assign n24123 = n24120 | n24121;
  assign n24124 = ~n24122 & n24123;
  assign n24125 = n52583 & n24124;
  assign n24126 = n52583 | n24124;
  assign n24127 = ~n24125 & n24126;
  assign n24128 = x116 & x212;
  assign n24129 = n24127 & n24128;
  assign n24130 = n24127 | n24128;
  assign n24131 = ~n24129 & n24130;
  assign n24132 = n52581 & n24131;
  assign n24133 = n52581 | n24131;
  assign n24134 = ~n24132 & n24133;
  assign n24135 = x115 & x213;
  assign n24136 = n24134 & n24135;
  assign n24137 = n24134 | n24135;
  assign n24138 = ~n24136 & n24137;
  assign n24139 = n52579 & n24138;
  assign n24140 = n52579 | n24138;
  assign n24141 = ~n24139 & n24140;
  assign n24142 = x114 & x214;
  assign n24143 = n24141 & n24142;
  assign n24144 = n24141 | n24142;
  assign n24145 = ~n24143 & n24144;
  assign n24146 = n52577 & n24145;
  assign n24147 = n52577 | n24145;
  assign n24148 = ~n24146 & n24147;
  assign n24149 = x113 & x215;
  assign n24150 = n24148 & n24149;
  assign n24151 = n24148 | n24149;
  assign n24152 = ~n24150 & n24151;
  assign n24153 = n23841 & n24152;
  assign n24154 = n23841 | n24152;
  assign n24155 = ~n24153 & n24154;
  assign n24156 = x112 & x216;
  assign n24157 = n24155 & n24156;
  assign n24158 = n24155 | n24156;
  assign n24159 = ~n24157 & n24158;
  assign n68156 = n23841 | n24149;
  assign n68157 = (n23841 & n24148) | (n23841 & n68156) | (n24148 & n68156);
  assign n52723 = (n24150 & n24152) | (n24150 & n68157) | (n24152 & n68157);
  assign n52724 = n24143 | n52577;
  assign n52725 = (n24143 & n24145) | (n24143 & n52724) | (n24145 & n52724);
  assign n52726 = n24136 | n52579;
  assign n52727 = (n24136 & n24138) | (n24136 & n52726) | (n24138 & n52726);
  assign n52728 = n24129 | n52581;
  assign n52729 = (n24129 & n24131) | (n24129 & n52728) | (n24131 & n52728);
  assign n52730 = n24122 | n52583;
  assign n52731 = (n24122 & n24124) | (n24122 & n52730) | (n24124 & n52730);
  assign n68158 = n24115 | n68061;
  assign n68159 = (n24115 & n24117) | (n24115 & n68158) | (n24117 & n68158);
  assign n24166 = n24108 | n24111;
  assign n24167 = n24101 | n24104;
  assign n52732 = n24094 | n24096;
  assign n52733 = (n23851 & n24094) | (n23851 & n52732) | (n24094 & n52732);
  assign n52734 = n24087 | n24089;
  assign n52735 = (n24087 & n52585) | (n24087 & n52734) | (n52585 & n52734);
  assign n52736 = n24080 | n24082;
  assign n52737 = (n24080 & n52587) | (n24080 & n52736) | (n52587 & n52736);
  assign n52738 = n24073 | n24075;
  assign n52739 = (n24073 & n52589) | (n24073 & n52738) | (n52589 & n52738);
  assign n52740 = n24066 | n24068;
  assign n52741 = (n24066 & n52591) | (n24066 & n52740) | (n52591 & n52740);
  assign n52595 = (n23743 & n52448) | (n23743 & n52594) | (n52448 & n52594);
  assign n52597 = (n23736 & n52450) | (n23736 & n52596) | (n52450 & n52596);
  assign n52602 = (n67964 & n68063) | (n67964 & n52601) | (n68063 & n52601);
  assign n52751 = n23975 | n23977;
  assign n68160 = n23666 | n23975;
  assign n68161 = (n23975 & n23977) | (n23975 & n68160) | (n23977 & n68160);
  assign n68162 = (n52537 & n52751) | (n52537 & n68161) | (n52751 & n68161);
  assign n68163 = (n52536 & n52751) | (n52536 & n68161) | (n52751 & n68161);
  assign n68164 = (n52328 & n68162) | (n52328 & n68163) | (n68162 & n68163);
  assign n52756 = n23954 | n23956;
  assign n68165 = n23645 | n23954;
  assign n68166 = (n23954 & n23956) | (n23954 & n68165) | (n23956 & n68165);
  assign n68167 = (n52527 & n52756) | (n52527 & n68166) | (n52756 & n68166);
  assign n68168 = (n52526 & n52756) | (n52526 & n68166) | (n52756 & n68166);
  assign n68169 = (n67894 & n68167) | (n67894 & n68168) | (n68167 & n68168);
  assign n68172 = n23919 | n23921;
  assign n68173 = (n23919 & n52616) | (n23919 & n68172) | (n52616 & n68172);
  assign n68174 = n23610 | n23919;
  assign n68175 = (n23919 & n23921) | (n23919 & n68174) | (n23921 & n68174);
  assign n68176 = (n52470 & n68173) | (n52470 & n68175) | (n68173 & n68175);
  assign n68177 = (n67995 & n68173) | (n67995 & n68175) | (n68173 & n68175);
  assign n68178 = (n67817 & n68176) | (n67817 & n68177) | (n68176 & n68177);
  assign n24199 = x153 & x176;
  assign n24200 = x152 & x177;
  assign n24201 = n24199 & n24200;
  assign n24202 = n24199 | n24200;
  assign n24203 = ~n24201 & n24202;
  assign n68185 = n23884 | n68078;
  assign n68188 = n24203 & n68185;
  assign n68186 = n23884 | n23886;
  assign n68189 = n24203 & n68186;
  assign n68190 = (n68000 & n68188) | (n68000 & n68189) | (n68188 & n68189);
  assign n68192 = (n68002 & n68188) | (n68002 & n68189) | (n68188 & n68189);
  assign n68193 = (n67658 & n68190) | (n67658 & n68192) | (n68190 & n68192);
  assign n68194 = (n67657 & n68190) | (n67657 & n68192) | (n68190 & n68192);
  assign n68195 = (n66988 & n68193) | (n66988 & n68194) | (n68193 & n68194);
  assign n68196 = n24203 | n68185;
  assign n68197 = n24203 | n68186;
  assign n68198 = (n68000 & n68196) | (n68000 & n68197) | (n68196 & n68197);
  assign n68199 = (n68002 & n68196) | (n68002 & n68197) | (n68196 & n68197);
  assign n68200 = (n67658 & n68198) | (n67658 & n68199) | (n68198 & n68199);
  assign n68201 = (n67657 & n68198) | (n67657 & n68199) | (n68198 & n68199);
  assign n68202 = (n66988 & n68200) | (n66988 & n68201) | (n68200 & n68201);
  assign n24206 = ~n68195 & n68202;
  assign n24207 = x151 & x178;
  assign n24208 = n24206 & n24207;
  assign n24209 = n24206 | n24207;
  assign n24210 = ~n24208 & n24209;
  assign n68203 = n23582 | n23891;
  assign n68204 = (n23891 & n23893) | (n23891 & n68203) | (n23893 & n68203);
  assign n52786 = n24210 & n68204;
  assign n52775 = n23891 | n23893;
  assign n52787 = n24210 & n52775;
  assign n68205 = (n52786 & n52787) | (n52786 & n68020) | (n52787 & n68020);
  assign n68206 = (n52786 & n52787) | (n52786 & n68019) | (n52787 & n68019);
  assign n68207 = (n67426 & n68205) | (n67426 & n68206) | (n68205 & n68206);
  assign n52789 = n24210 | n68204;
  assign n52790 = n24210 | n52775;
  assign n68208 = (n52789 & n52790) | (n52789 & n68020) | (n52790 & n68020);
  assign n68209 = (n52789 & n52790) | (n52789 & n68019) | (n52790 & n68019);
  assign n68210 = (n67426 & n68208) | (n67426 & n68209) | (n68208 & n68209);
  assign n24213 = ~n68207 & n68210;
  assign n24214 = x150 & x179;
  assign n24215 = n24213 & n24214;
  assign n24216 = n24213 | n24214;
  assign n24217 = ~n24215 & n24216;
  assign n68182 = n23898 | n23900;
  assign n68183 = (n23898 & n68097) | (n23898 & n68182) | (n68097 & n68182);
  assign n68211 = n24217 & n68183;
  assign n68184 = (n23898 & n68099) | (n23898 & n68182) | (n68099 & n68182);
  assign n68212 = n24217 & n68184;
  assign n68213 = (n67914 & n68211) | (n67914 & n68212) | (n68211 & n68212);
  assign n68214 = n24217 | n68183;
  assign n68215 = n24217 | n68184;
  assign n68216 = (n67914 & n68214) | (n67914 & n68215) | (n68214 & n68215);
  assign n24220 = ~n68213 & n68216;
  assign n24221 = x149 & x180;
  assign n24222 = n24220 & n24221;
  assign n24223 = n24220 | n24221;
  assign n24224 = ~n24222 & n24223;
  assign n68179 = n23905 | n23907;
  assign n68181 = (n23905 & n52622) | (n23905 & n68179) | (n52622 & n68179);
  assign n68217 = n24224 & n68181;
  assign n68180 = (n23905 & n68101) | (n23905 & n68179) | (n68101 & n68179);
  assign n68218 = n24224 & n68180;
  assign n68219 = (n67940 & n68217) | (n67940 & n68218) | (n68217 & n68218);
  assign n68220 = n24224 | n68181;
  assign n68221 = n24224 | n68180;
  assign n68222 = (n67940 & n68220) | (n67940 & n68221) | (n68220 & n68221);
  assign n24227 = ~n68219 & n68222;
  assign n24228 = x148 & x181;
  assign n24229 = n24227 & n24228;
  assign n24230 = n24227 | n24228;
  assign n24231 = ~n24229 & n24230;
  assign n52792 = n23912 & n24231;
  assign n68223 = (n24231 & n52653) | (n24231 & n52792) | (n52653 & n52792);
  assign n68224 = (n24231 & n52792) | (n24231 & n68103) | (n52792 & n68103);
  assign n68225 = (n67908 & n68223) | (n67908 & n68224) | (n68223 & n68224);
  assign n52794 = n23912 | n24231;
  assign n68226 = n52653 | n52794;
  assign n68227 = n52794 | n68103;
  assign n68228 = (n67908 & n68226) | (n67908 & n68227) | (n68226 & n68227);
  assign n24234 = ~n68225 & n68228;
  assign n24235 = x147 & x182;
  assign n24236 = n24234 & n24235;
  assign n24237 = n24234 | n24235;
  assign n24238 = ~n24236 & n24237;
  assign n24239 = n68178 & n24238;
  assign n24240 = n68178 | n24238;
  assign n24241 = ~n24239 & n24240;
  assign n24242 = x146 & x183;
  assign n24243 = n24241 & n24242;
  assign n24244 = n24241 | n24242;
  assign n24245 = ~n24243 & n24244;
  assign n52763 = n23926 | n23928;
  assign n52796 = n24245 & n52763;
  assign n52797 = n23926 & n24245;
  assign n68229 = (n52796 & n52797) | (n52796 & n68077) | (n52797 & n68077);
  assign n68230 = (n52796 & n52797) | (n52796 & n68075) | (n52797 & n68075);
  assign n68231 = (n52341 & n68229) | (n52341 & n68230) | (n68229 & n68230);
  assign n52799 = n24245 | n52763;
  assign n52800 = n23926 | n24245;
  assign n68232 = (n52799 & n52800) | (n52799 & n68077) | (n52800 & n68077);
  assign n68233 = (n52799 & n52800) | (n52799 & n68075) | (n52800 & n68075);
  assign n68234 = (n52341 & n68232) | (n52341 & n68233) | (n68232 & n68233);
  assign n24248 = ~n68231 & n68234;
  assign n24249 = x145 & x184;
  assign n24250 = n24248 & n24249;
  assign n24251 = n24248 | n24249;
  assign n24252 = ~n24250 & n24251;
  assign n52761 = n23933 | n23935;
  assign n68235 = n24252 & n52761;
  assign n68170 = n23624 | n23933;
  assign n68171 = (n23933 & n23935) | (n23933 & n68170) | (n23935 & n68170);
  assign n68236 = n24252 & n68171;
  assign n68237 = (n52518 & n68235) | (n52518 & n68236) | (n68235 & n68236);
  assign n68238 = n24252 | n52761;
  assign n68239 = n24252 | n68171;
  assign n68240 = (n52518 & n68238) | (n52518 & n68239) | (n68238 & n68239);
  assign n24255 = ~n68237 & n68240;
  assign n24256 = x144 & x185;
  assign n24257 = n24255 & n24256;
  assign n24258 = n24255 | n24256;
  assign n24259 = ~n24257 & n24258;
  assign n52758 = n23940 | n23942;
  assign n52802 = n24259 & n52758;
  assign n52803 = n23940 & n24259;
  assign n52804 = (n68073 & n52802) | (n68073 & n52803) | (n52802 & n52803);
  assign n52805 = n24259 | n52758;
  assign n52806 = n23940 | n24259;
  assign n52807 = (n68073 & n52805) | (n68073 & n52806) | (n52805 & n52806);
  assign n24262 = ~n52804 & n52807;
  assign n24263 = x143 & x186;
  assign n24264 = n24262 & n24263;
  assign n24265 = n24262 | n24263;
  assign n24266 = ~n24264 & n24265;
  assign n52808 = n23947 & n24266;
  assign n68241 = (n24266 & n52669) | (n24266 & n52808) | (n52669 & n52808);
  assign n68242 = (n24266 & n52668) | (n24266 & n52808) | (n52668 & n52808);
  assign n68243 = (n67993 & n68241) | (n67993 & n68242) | (n68241 & n68242);
  assign n52810 = n23947 | n24266;
  assign n68244 = n52669 | n52810;
  assign n68245 = n52668 | n52810;
  assign n68246 = (n67993 & n68244) | (n67993 & n68245) | (n68244 & n68245);
  assign n24269 = ~n68243 & n68246;
  assign n24270 = x142 & x187;
  assign n24271 = n24269 & n24270;
  assign n24272 = n24269 | n24270;
  assign n24273 = ~n24271 & n24272;
  assign n24274 = n68169 & n24273;
  assign n24275 = n68169 | n24273;
  assign n24276 = ~n24274 & n24275;
  assign n24277 = x141 & x188;
  assign n24278 = n24276 & n24277;
  assign n24279 = n24276 | n24277;
  assign n24280 = ~n24278 & n24279;
  assign n52753 = n23961 | n23963;
  assign n52812 = n24280 & n52753;
  assign n52813 = n23961 & n24280;
  assign n52814 = (n68068 & n52812) | (n68068 & n52813) | (n52812 & n52813);
  assign n52815 = n24280 | n52753;
  assign n52816 = n23961 | n24280;
  assign n52817 = (n68068 & n52815) | (n68068 & n52816) | (n52815 & n52816);
  assign n24283 = ~n52814 & n52817;
  assign n24284 = x140 & x189;
  assign n24285 = n24283 & n24284;
  assign n24286 = n24283 | n24284;
  assign n24287 = ~n24285 & n24286;
  assign n52818 = n23968 & n24287;
  assign n68247 = (n24287 & n52679) | (n24287 & n52818) | (n52679 & n52818);
  assign n68248 = (n24287 & n52678) | (n24287 & n52818) | (n52678 & n52818);
  assign n68249 = (n67988 & n68247) | (n67988 & n68248) | (n68247 & n68248);
  assign n52820 = n23968 | n24287;
  assign n68250 = n52679 | n52820;
  assign n68251 = n52678 | n52820;
  assign n68252 = (n67988 & n68250) | (n67988 & n68251) | (n68250 & n68251);
  assign n24290 = ~n68249 & n68252;
  assign n24291 = x139 & x190;
  assign n24292 = n24290 & n24291;
  assign n24293 = n24290 | n24291;
  assign n24294 = ~n24292 & n24293;
  assign n24295 = n68164 & n24294;
  assign n24296 = n68164 | n24294;
  assign n24297 = ~n24295 & n24296;
  assign n24298 = x138 & x191;
  assign n24299 = n24297 & n24298;
  assign n24300 = n24297 | n24298;
  assign n24301 = ~n24299 & n24300;
  assign n52748 = n23982 | n23984;
  assign n52822 = n24301 & n52748;
  assign n52823 = n23982 & n24301;
  assign n52824 = (n52602 & n52822) | (n52602 & n52823) | (n52822 & n52823);
  assign n52825 = n24301 | n52748;
  assign n52826 = n23982 | n24301;
  assign n52827 = (n52602 & n52825) | (n52602 & n52826) | (n52825 & n52826);
  assign n24304 = ~n52824 & n52827;
  assign n24305 = x137 & x192;
  assign n24306 = n24304 & n24305;
  assign n24307 = n24304 | n24305;
  assign n24308 = ~n24306 & n24307;
  assign n52828 = n23989 & n24308;
  assign n52829 = (n24308 & n68140) | (n24308 & n52828) | (n68140 & n52828);
  assign n52830 = n23989 | n24308;
  assign n52831 = n68140 | n52830;
  assign n24311 = ~n52829 & n52831;
  assign n24312 = x136 & x193;
  assign n24313 = n24311 & n24312;
  assign n24314 = n24311 | n24312;
  assign n24315 = ~n24313 & n24314;
  assign n52832 = n23996 & n24315;
  assign n52833 = (n24315 & n52693) | (n24315 & n52832) | (n52693 & n52832);
  assign n52834 = n23996 | n24315;
  assign n52835 = n52693 | n52834;
  assign n24318 = ~n52833 & n52835;
  assign n24319 = x135 & x194;
  assign n24320 = n24318 & n24319;
  assign n24321 = n24318 | n24319;
  assign n24322 = ~n24320 & n24321;
  assign n52836 = n24003 & n24322;
  assign n52837 = (n24322 & n52697) | (n24322 & n52836) | (n52697 & n52836);
  assign n52838 = n24003 | n24322;
  assign n52839 = n52697 | n52838;
  assign n24325 = ~n52837 & n52839;
  assign n24326 = x134 & x195;
  assign n24327 = n24325 & n24326;
  assign n24328 = n24325 | n24326;
  assign n24329 = ~n24327 & n24328;
  assign n52840 = n24010 & n24329;
  assign n52841 = (n24329 & n52701) | (n24329 & n52840) | (n52701 & n52840);
  assign n52842 = n24010 | n24329;
  assign n52843 = n52701 | n52842;
  assign n24332 = ~n52841 & n52843;
  assign n24333 = x133 & x196;
  assign n24334 = n24332 & n24333;
  assign n24335 = n24332 | n24333;
  assign n24336 = ~n24334 & n24335;
  assign n52844 = n24017 & n24336;
  assign n52845 = (n24336 & n52705) | (n24336 & n52844) | (n52705 & n52844);
  assign n52846 = n24017 | n24336;
  assign n52847 = n52705 | n52846;
  assign n24339 = ~n52845 & n52847;
  assign n24340 = x132 & x197;
  assign n24341 = n24339 & n24340;
  assign n24342 = n24339 | n24340;
  assign n24343 = ~n24341 & n24342;
  assign n52848 = n24024 & n24343;
  assign n52849 = (n24343 & n52709) | (n24343 & n52848) | (n52709 & n52848);
  assign n52850 = n24024 | n24343;
  assign n52851 = n52709 | n52850;
  assign n24346 = ~n52849 & n52851;
  assign n24347 = x131 & x198;
  assign n24348 = n24346 & n24347;
  assign n24349 = n24346 | n24347;
  assign n24350 = ~n24348 & n24349;
  assign n52852 = n24031 & n24350;
  assign n52853 = (n24350 & n52713) | (n24350 & n52852) | (n52713 & n52852);
  assign n52854 = n24031 | n24350;
  assign n52855 = n52713 | n52854;
  assign n24353 = ~n52853 & n52855;
  assign n24354 = x130 & x199;
  assign n24355 = n24353 & n24354;
  assign n24356 = n24353 | n24354;
  assign n24357 = ~n24355 & n24356;
  assign n52856 = n24038 & n24357;
  assign n52857 = (n24357 & n52718) | (n24357 & n52856) | (n52718 & n52856);
  assign n52858 = n24038 | n24357;
  assign n52859 = n52718 | n52858;
  assign n24360 = ~n52857 & n52859;
  assign n24361 = x129 & x200;
  assign n24362 = n24360 & n24361;
  assign n24363 = n24360 | n24361;
  assign n24364 = ~n24362 & n24363;
  assign n52746 = n24045 | n24047;
  assign n52860 = n24364 & n52746;
  assign n52861 = n24045 & n24364;
  assign n52862 = (n52597 & n52860) | (n52597 & n52861) | (n52860 & n52861);
  assign n52863 = n24364 | n52746;
  assign n52864 = n24045 | n24364;
  assign n52865 = (n52597 & n52863) | (n52597 & n52864) | (n52863 & n52864);
  assign n24367 = ~n52862 & n52865;
  assign n24368 = x128 & x201;
  assign n24369 = n24367 & n24368;
  assign n24370 = n24367 | n24368;
  assign n24371 = ~n24369 & n24370;
  assign n52744 = n24052 | n24054;
  assign n68253 = n24371 & n52744;
  assign n68254 = n24052 & n24371;
  assign n68255 = (n52595 & n68253) | (n52595 & n68254) | (n68253 & n68254);
  assign n68256 = n24371 | n52744;
  assign n68257 = n24052 | n24371;
  assign n68258 = (n52595 & n68256) | (n52595 & n68257) | (n68256 & n68257);
  assign n24374 = ~n68255 & n68258;
  assign n24375 = x127 & x202;
  assign n24376 = n24374 & n24375;
  assign n24377 = n24374 | n24375;
  assign n24378 = ~n24376 & n24377;
  assign n52742 = n24059 | n24061;
  assign n68259 = n24378 & n52742;
  assign n68260 = n24059 & n24378;
  assign n68261 = (n52593 & n68259) | (n52593 & n68260) | (n68259 & n68260);
  assign n68262 = n24378 | n52742;
  assign n68263 = n24059 | n24378;
  assign n68264 = (n52593 & n68262) | (n52593 & n68263) | (n68262 & n68263);
  assign n24381 = ~n68261 & n68264;
  assign n24382 = x126 & x203;
  assign n24383 = n24381 & n24382;
  assign n24384 = n24381 | n24382;
  assign n24385 = ~n24383 & n24384;
  assign n24386 = n52741 & n24385;
  assign n24387 = n52741 | n24385;
  assign n24388 = ~n24386 & n24387;
  assign n24389 = x125 & x204;
  assign n24390 = n24388 & n24389;
  assign n24391 = n24388 | n24389;
  assign n24392 = ~n24390 & n24391;
  assign n24393 = n52739 & n24392;
  assign n24394 = n52739 | n24392;
  assign n24395 = ~n24393 & n24394;
  assign n24396 = x124 & x205;
  assign n24397 = n24395 & n24396;
  assign n24398 = n24395 | n24396;
  assign n24399 = ~n24397 & n24398;
  assign n24400 = n52737 & n24399;
  assign n24401 = n52737 | n24399;
  assign n24402 = ~n24400 & n24401;
  assign n24403 = x123 & x206;
  assign n24404 = n24402 & n24403;
  assign n24405 = n24402 | n24403;
  assign n24406 = ~n24404 & n24405;
  assign n24407 = n52735 & n24406;
  assign n24408 = n52735 | n24406;
  assign n24409 = ~n24407 & n24408;
  assign n24410 = x122 & x207;
  assign n24411 = n24409 & n24410;
  assign n24412 = n24409 | n24410;
  assign n24413 = ~n24411 & n24412;
  assign n24414 = n52733 & n24413;
  assign n24415 = n52733 | n24413;
  assign n24416 = ~n24414 & n24415;
  assign n24417 = x121 & x208;
  assign n24418 = n24416 & n24417;
  assign n24419 = n24416 | n24417;
  assign n24420 = ~n24418 & n24419;
  assign n24421 = n24167 & n24420;
  assign n24422 = n24167 | n24420;
  assign n24423 = ~n24421 & n24422;
  assign n24424 = x120 & x209;
  assign n24425 = n24423 & n24424;
  assign n24426 = n24423 | n24424;
  assign n24427 = ~n24425 & n24426;
  assign n24428 = n24166 & n24427;
  assign n24429 = n24166 | n24427;
  assign n24430 = ~n24428 & n24429;
  assign n24431 = x119 & x210;
  assign n24432 = n24430 & n24431;
  assign n24433 = n24430 | n24431;
  assign n24434 = ~n24432 & n24433;
  assign n24435 = n68159 & n24434;
  assign n24436 = n68159 | n24434;
  assign n24437 = ~n24435 & n24436;
  assign n24438 = x118 & x211;
  assign n24439 = n24437 & n24438;
  assign n24440 = n24437 | n24438;
  assign n24441 = ~n24439 & n24440;
  assign n24442 = n52731 & n24441;
  assign n24443 = n52731 | n24441;
  assign n24444 = ~n24442 & n24443;
  assign n24445 = x117 & x212;
  assign n24446 = n24444 & n24445;
  assign n24447 = n24444 | n24445;
  assign n24448 = ~n24446 & n24447;
  assign n24449 = n52729 & n24448;
  assign n24450 = n52729 | n24448;
  assign n24451 = ~n24449 & n24450;
  assign n24452 = x116 & x213;
  assign n24453 = n24451 & n24452;
  assign n24454 = n24451 | n24452;
  assign n24455 = ~n24453 & n24454;
  assign n24456 = n52727 & n24455;
  assign n24457 = n52727 | n24455;
  assign n24458 = ~n24456 & n24457;
  assign n24459 = x115 & x214;
  assign n24460 = n24458 & n24459;
  assign n24461 = n24458 | n24459;
  assign n24462 = ~n24460 & n24461;
  assign n24463 = n52725 & n24462;
  assign n24464 = n52725 | n24462;
  assign n24465 = ~n24463 & n24464;
  assign n24466 = x114 & x215;
  assign n24467 = n24465 & n24466;
  assign n24468 = n24465 | n24466;
  assign n24469 = ~n24467 & n24468;
  assign n24470 = n52723 & n24469;
  assign n24471 = n52723 | n24469;
  assign n24472 = ~n24470 & n24471;
  assign n24473 = x113 & x216;
  assign n24474 = n24472 & n24473;
  assign n24475 = n24472 | n24473;
  assign n24476 = ~n24474 & n24475;
  assign n24477 = n24157 & n24476;
  assign n24478 = n24157 | n24476;
  assign n24479 = ~n24477 & n24478;
  assign n24480 = x112 & x217;
  assign n24481 = n24479 & n24480;
  assign n24482 = n24479 | n24480;
  assign n24483 = ~n24481 & n24482;
  assign n68265 = n24157 | n24473;
  assign n68266 = (n24157 & n24472) | (n24157 & n68265) | (n24472 & n68265);
  assign n52867 = (n24474 & n24476) | (n24474 & n68266) | (n24476 & n68266);
  assign n52868 = n24467 | n52723;
  assign n52869 = (n24467 & n24469) | (n24467 & n52868) | (n24469 & n52868);
  assign n52870 = n24460 | n52725;
  assign n52871 = (n24460 & n24462) | (n24460 & n52870) | (n24462 & n52870);
  assign n52872 = n24453 | n52727;
  assign n52873 = (n24453 & n24455) | (n24453 & n52872) | (n24455 & n52872);
  assign n52874 = n24446 | n52729;
  assign n52875 = (n24446 & n24448) | (n24446 & n52874) | (n24448 & n52874);
  assign n52876 = n24439 | n52731;
  assign n52877 = (n24439 & n24441) | (n24439 & n52876) | (n24441 & n52876);
  assign n68267 = n24432 | n68159;
  assign n68268 = (n24432 & n24434) | (n24432 & n68267) | (n24434 & n68267);
  assign n24491 = n24425 | n24428;
  assign n52878 = n24418 | n24420;
  assign n52879 = (n24167 & n24418) | (n24167 & n52878) | (n24418 & n52878);
  assign n52880 = n24411 | n24413;
  assign n52881 = (n24411 & n52733) | (n24411 & n52880) | (n52733 & n52880);
  assign n52882 = n24404 | n24406;
  assign n52883 = (n24404 & n52735) | (n24404 & n52882) | (n52735 & n52882);
  assign n52884 = n24397 | n24399;
  assign n52885 = (n24397 & n52737) | (n24397 & n52884) | (n52737 & n52884);
  assign n52886 = n24390 | n24392;
  assign n52887 = (n24390 & n52739) | (n24390 & n52886) | (n52739 & n52886);
  assign n52743 = (n24059 & n52593) | (n24059 & n52742) | (n52593 & n52742);
  assign n52745 = (n24052 & n52595) | (n24052 & n52744) | (n52595 & n52744);
  assign n52900 = n24285 | n24287;
  assign n68271 = n23968 | n24285;
  assign n68272 = (n24285 & n24287) | (n24285 & n68271) | (n24287 & n68271);
  assign n68273 = (n52679 & n52900) | (n52679 & n68272) | (n52900 & n68272);
  assign n68274 = (n52678 & n52900) | (n52678 & n68272) | (n52900 & n68272);
  assign n68275 = (n67988 & n68273) | (n67988 & n68274) | (n68273 & n68274);
  assign n52905 = n24264 | n24266;
  assign n68276 = n23947 | n24264;
  assign n68277 = (n24264 & n24266) | (n24264 & n68276) | (n24266 & n68276);
  assign n68278 = (n52669 & n52905) | (n52669 & n68277) | (n52905 & n68277);
  assign n68279 = (n52668 & n52905) | (n52668 & n68277) | (n52905 & n68277);
  assign n68280 = (n67993 & n68278) | (n67993 & n68279) | (n68278 & n68279);
  assign n52615 = (n52341 & n68075) | (n52341 & n68077) | (n68075 & n68077);
  assign n24524 = x154 & x176;
  assign n24525 = x153 & x177;
  assign n24526 = n24524 & n24525;
  assign n24527 = n24524 | n24525;
  assign n24528 = ~n24526 & n24527;
  assign n52924 = n24201 & n24528;
  assign n52925 = (n24528 & n68195) | (n24528 & n52924) | (n68195 & n52924);
  assign n52926 = n24201 | n24528;
  assign n52927 = n68195 | n52926;
  assign n24531 = ~n52925 & n52927;
  assign n24532 = x152 & x178;
  assign n24533 = n24531 & n24532;
  assign n24534 = n24531 | n24532;
  assign n24535 = ~n24533 & n24534;
  assign n68283 = n24208 | n24210;
  assign n68284 = (n24208 & n68204) | (n24208 & n68283) | (n68204 & n68283);
  assign n52928 = n24535 & n68284;
  assign n68285 = (n24208 & n52775) | (n24208 & n68283) | (n52775 & n68283);
  assign n52929 = n24535 & n68285;
  assign n68286 = (n52928 & n52929) | (n52928 & n68020) | (n52929 & n68020);
  assign n68287 = (n52928 & n52929) | (n52928 & n68019) | (n52929 & n68019);
  assign n68288 = (n67426 & n68286) | (n67426 & n68287) | (n68286 & n68287);
  assign n52931 = n24535 | n68284;
  assign n52932 = n24535 | n68285;
  assign n68289 = (n52931 & n52932) | (n52931 & n68020) | (n52932 & n68020);
  assign n68290 = (n52931 & n52932) | (n52931 & n68019) | (n52932 & n68019);
  assign n68291 = (n67426 & n68289) | (n67426 & n68290) | (n68289 & n68290);
  assign n24538 = ~n68288 & n68291;
  assign n24539 = x151 & x179;
  assign n24540 = n24538 & n24539;
  assign n24541 = n24538 | n24539;
  assign n24542 = ~n24540 & n24541;
  assign n52919 = n24215 | n24217;
  assign n52934 = n24542 & n52919;
  assign n52935 = n24215 & n24542;
  assign n68292 = (n52934 & n52935) | (n52934 & n68183) | (n52935 & n68183);
  assign n68293 = (n52934 & n52935) | (n52934 & n68184) | (n52935 & n68184);
  assign n68294 = (n67914 & n68292) | (n67914 & n68293) | (n68292 & n68293);
  assign n52937 = n24542 | n52919;
  assign n52938 = n24215 | n24542;
  assign n68295 = (n52937 & n52938) | (n52937 & n68183) | (n52938 & n68183);
  assign n68296 = (n52937 & n52938) | (n52937 & n68184) | (n52938 & n68184);
  assign n68297 = (n67914 & n68295) | (n67914 & n68296) | (n68295 & n68296);
  assign n24545 = ~n68294 & n68297;
  assign n24546 = x150 & x180;
  assign n24547 = n24545 & n24546;
  assign n24548 = n24545 | n24546;
  assign n24549 = ~n24547 & n24548;
  assign n52917 = n24222 | n24224;
  assign n52940 = n24549 & n52917;
  assign n52941 = n24222 & n24549;
  assign n68298 = (n52940 & n52941) | (n52940 & n68181) | (n52941 & n68181);
  assign n68299 = (n52940 & n52941) | (n52940 & n68180) | (n52941 & n68180);
  assign n68300 = (n67940 & n68298) | (n67940 & n68299) | (n68298 & n68299);
  assign n52943 = n24549 | n52917;
  assign n52944 = n24222 | n24549;
  assign n68301 = (n52943 & n52944) | (n52943 & n68181) | (n52944 & n68181);
  assign n68302 = (n52943 & n52944) | (n52943 & n68180) | (n52944 & n68180);
  assign n68303 = (n67940 & n68301) | (n67940 & n68302) | (n68301 & n68302);
  assign n24552 = ~n68300 & n68303;
  assign n24553 = x149 & x181;
  assign n24554 = n24552 & n24553;
  assign n24555 = n24552 | n24553;
  assign n24556 = ~n24554 & n24555;
  assign n68304 = n23912 | n24229;
  assign n68305 = (n24229 & n24231) | (n24229 & n68304) | (n24231 & n68304);
  assign n52946 = n24556 & n68305;
  assign n52915 = n24229 | n24231;
  assign n52947 = n24556 & n52915;
  assign n68306 = (n52653 & n52946) | (n52653 & n52947) | (n52946 & n52947);
  assign n68307 = (n52946 & n52947) | (n52946 & n68103) | (n52947 & n68103);
  assign n68308 = (n67908 & n68306) | (n67908 & n68307) | (n68306 & n68307);
  assign n52949 = n24556 | n68305;
  assign n52950 = n24556 | n52915;
  assign n68309 = (n52653 & n52949) | (n52653 & n52950) | (n52949 & n52950);
  assign n68310 = (n52949 & n52950) | (n52949 & n68103) | (n52950 & n68103);
  assign n68311 = (n67908 & n68309) | (n67908 & n68310) | (n68309 & n68310);
  assign n24559 = ~n68308 & n68311;
  assign n24560 = x148 & x182;
  assign n24561 = n24559 & n24560;
  assign n24562 = n24559 | n24560;
  assign n24563 = ~n24561 & n24562;
  assign n52912 = n24236 | n24238;
  assign n52952 = n24563 & n52912;
  assign n52953 = n24236 & n24563;
  assign n52954 = (n68178 & n52952) | (n68178 & n52953) | (n52952 & n52953);
  assign n52955 = n24563 | n52912;
  assign n52956 = n24236 | n24563;
  assign n52957 = (n68178 & n52955) | (n68178 & n52956) | (n52955 & n52956);
  assign n24566 = ~n52954 & n52957;
  assign n24567 = x147 & x183;
  assign n24568 = n24566 & n24567;
  assign n24569 = n24566 | n24567;
  assign n24570 = ~n24568 & n24569;
  assign n52910 = n24243 | n52796;
  assign n68312 = n24570 & n52910;
  assign n68281 = n23926 | n24243;
  assign n68282 = (n24243 & n24245) | (n24243 & n68281) | (n24245 & n68281);
  assign n68313 = n24570 & n68282;
  assign n68314 = (n52615 & n68312) | (n52615 & n68313) | (n68312 & n68313);
  assign n68315 = n24570 | n52910;
  assign n68316 = n24570 | n68282;
  assign n68317 = (n52615 & n68315) | (n52615 & n68316) | (n68315 & n68316);
  assign n24573 = ~n68314 & n68317;
  assign n24574 = x146 & x184;
  assign n24575 = n24573 & n24574;
  assign n24576 = n24573 | n24574;
  assign n24577 = ~n24575 & n24576;
  assign n52907 = n24250 | n24252;
  assign n52958 = n24577 & n52907;
  assign n52959 = n24250 & n24577;
  assign n68318 = (n52761 & n52958) | (n52761 & n52959) | (n52958 & n52959);
  assign n68319 = (n52958 & n52959) | (n52958 & n68171) | (n52959 & n68171);
  assign n68320 = (n52518 & n68318) | (n52518 & n68319) | (n68318 & n68319);
  assign n52961 = n24577 | n52907;
  assign n52962 = n24250 | n24577;
  assign n68321 = (n52761 & n52961) | (n52761 & n52962) | (n52961 & n52962);
  assign n68322 = (n52961 & n52962) | (n52961 & n68171) | (n52962 & n68171);
  assign n68323 = (n52518 & n68321) | (n52518 & n68322) | (n68321 & n68322);
  assign n24580 = ~n68320 & n68323;
  assign n24581 = x145 & x185;
  assign n24582 = n24580 & n24581;
  assign n24583 = n24580 | n24581;
  assign n24584 = ~n24582 & n24583;
  assign n52964 = n24257 & n24584;
  assign n52965 = (n24584 & n52804) | (n24584 & n52964) | (n52804 & n52964);
  assign n52966 = n24257 | n24584;
  assign n52967 = n52804 | n52966;
  assign n24587 = ~n52965 & n52967;
  assign n24588 = x144 & x186;
  assign n24589 = n24587 & n24588;
  assign n24590 = n24587 | n24588;
  assign n24591 = ~n24589 & n24590;
  assign n24592 = n68280 & n24591;
  assign n24593 = n68280 | n24591;
  assign n24594 = ~n24592 & n24593;
  assign n24595 = x143 & x187;
  assign n24596 = n24594 & n24595;
  assign n24597 = n24594 | n24595;
  assign n24598 = ~n24596 & n24597;
  assign n52902 = n24271 | n24273;
  assign n52968 = n24598 & n52902;
  assign n52969 = n24271 & n24598;
  assign n52970 = (n68169 & n52968) | (n68169 & n52969) | (n52968 & n52969);
  assign n52971 = n24598 | n52902;
  assign n52972 = n24271 | n24598;
  assign n52973 = (n68169 & n52971) | (n68169 & n52972) | (n52971 & n52972);
  assign n24601 = ~n52970 & n52973;
  assign n24602 = x142 & x188;
  assign n24603 = n24601 & n24602;
  assign n24604 = n24601 | n24602;
  assign n24605 = ~n24603 & n24604;
  assign n52974 = n24278 & n24605;
  assign n68324 = (n24605 & n52813) | (n24605 & n52974) | (n52813 & n52974);
  assign n68325 = (n24605 & n52812) | (n24605 & n52974) | (n52812 & n52974);
  assign n68326 = (n68068 & n68324) | (n68068 & n68325) | (n68324 & n68325);
  assign n52976 = n24278 | n24605;
  assign n68327 = n52813 | n52976;
  assign n68328 = n52812 | n52976;
  assign n68329 = (n68068 & n68327) | (n68068 & n68328) | (n68327 & n68328);
  assign n24608 = ~n68326 & n68329;
  assign n24609 = x141 & x189;
  assign n24610 = n24608 & n24609;
  assign n24611 = n24608 | n24609;
  assign n24612 = ~n24610 & n24611;
  assign n24613 = n68275 & n24612;
  assign n24614 = n68275 | n24612;
  assign n24615 = ~n24613 & n24614;
  assign n24616 = x140 & x190;
  assign n24617 = n24615 & n24616;
  assign n24618 = n24615 | n24616;
  assign n24619 = ~n24617 & n24618;
  assign n52897 = n24292 | n24294;
  assign n52978 = n24619 & n52897;
  assign n52979 = n24292 & n24619;
  assign n52980 = (n68164 & n52978) | (n68164 & n52979) | (n52978 & n52979);
  assign n52981 = n24619 | n52897;
  assign n52982 = n24292 | n24619;
  assign n52983 = (n68164 & n52981) | (n68164 & n52982) | (n52981 & n52982);
  assign n24622 = ~n52980 & n52983;
  assign n24623 = x139 & x191;
  assign n24624 = n24622 & n24623;
  assign n24625 = n24622 | n24623;
  assign n24626 = ~n24624 & n24625;
  assign n52984 = n24299 & n24626;
  assign n68330 = (n24626 & n52823) | (n24626 & n52984) | (n52823 & n52984);
  assign n68331 = (n24626 & n52822) | (n24626 & n52984) | (n52822 & n52984);
  assign n68332 = (n52602 & n68330) | (n52602 & n68331) | (n68330 & n68331);
  assign n52986 = n24299 | n24626;
  assign n68333 = n52823 | n52986;
  assign n68334 = n52822 | n52986;
  assign n68335 = (n52602 & n68333) | (n52602 & n68334) | (n68333 & n68334);
  assign n24629 = ~n68332 & n68335;
  assign n24630 = x138 & x192;
  assign n24631 = n24629 & n24630;
  assign n24632 = n24629 | n24630;
  assign n24633 = ~n24631 & n24632;
  assign n52895 = n24306 | n24308;
  assign n68336 = n24633 & n52895;
  assign n68269 = n23989 | n24306;
  assign n68270 = (n24306 & n24308) | (n24306 & n68269) | (n24308 & n68269);
  assign n68337 = n24633 & n68270;
  assign n68338 = (n68140 & n68336) | (n68140 & n68337) | (n68336 & n68337);
  assign n68339 = n24633 | n52895;
  assign n68340 = n24633 | n68270;
  assign n68341 = (n68140 & n68339) | (n68140 & n68340) | (n68339 & n68340);
  assign n24636 = ~n68338 & n68341;
  assign n24637 = x137 & x193;
  assign n24638 = n24636 & n24637;
  assign n24639 = n24636 | n24637;
  assign n24640 = ~n24638 & n24639;
  assign n52988 = n24313 & n24640;
  assign n68342 = (n24640 & n52832) | (n24640 & n52988) | (n52832 & n52988);
  assign n68343 = (n24315 & n24640) | (n24315 & n52988) | (n24640 & n52988);
  assign n68344 = (n52693 & n68342) | (n52693 & n68343) | (n68342 & n68343);
  assign n52990 = n24313 | n24640;
  assign n68345 = n52832 | n52990;
  assign n68346 = n24315 | n52990;
  assign n68347 = (n52693 & n68345) | (n52693 & n68346) | (n68345 & n68346);
  assign n24643 = ~n68344 & n68347;
  assign n24644 = x136 & x194;
  assign n24645 = n24643 & n24644;
  assign n24646 = n24643 | n24644;
  assign n24647 = ~n24645 & n24646;
  assign n52992 = n24320 & n24647;
  assign n52993 = (n24647 & n52837) | (n24647 & n52992) | (n52837 & n52992);
  assign n52994 = n24320 | n24647;
  assign n52995 = n52837 | n52994;
  assign n24650 = ~n52993 & n52995;
  assign n24651 = x135 & x195;
  assign n24652 = n24650 & n24651;
  assign n24653 = n24650 | n24651;
  assign n24654 = ~n24652 & n24653;
  assign n52996 = n24327 & n24654;
  assign n52997 = (n24654 & n52841) | (n24654 & n52996) | (n52841 & n52996);
  assign n52998 = n24327 | n24654;
  assign n52999 = n52841 | n52998;
  assign n24657 = ~n52997 & n52999;
  assign n24658 = x134 & x196;
  assign n24659 = n24657 & n24658;
  assign n24660 = n24657 | n24658;
  assign n24661 = ~n24659 & n24660;
  assign n53000 = n24334 & n24661;
  assign n53001 = (n24661 & n52845) | (n24661 & n53000) | (n52845 & n53000);
  assign n53002 = n24334 | n24661;
  assign n53003 = n52845 | n53002;
  assign n24664 = ~n53001 & n53003;
  assign n24665 = x133 & x197;
  assign n24666 = n24664 & n24665;
  assign n24667 = n24664 | n24665;
  assign n24668 = ~n24666 & n24667;
  assign n53004 = n24341 & n24668;
  assign n53005 = (n24668 & n52849) | (n24668 & n53004) | (n52849 & n53004);
  assign n53006 = n24341 | n24668;
  assign n53007 = n52849 | n53006;
  assign n24671 = ~n53005 & n53007;
  assign n24672 = x132 & x198;
  assign n24673 = n24671 & n24672;
  assign n24674 = n24671 | n24672;
  assign n24675 = ~n24673 & n24674;
  assign n53008 = n24348 & n24675;
  assign n53009 = (n24675 & n52853) | (n24675 & n53008) | (n52853 & n53008);
  assign n53010 = n24348 | n24675;
  assign n53011 = n52853 | n53010;
  assign n24678 = ~n53009 & n53011;
  assign n24679 = x131 & x199;
  assign n24680 = n24678 & n24679;
  assign n24681 = n24678 | n24679;
  assign n24682 = ~n24680 & n24681;
  assign n53012 = n24355 & n24682;
  assign n53013 = (n24682 & n52857) | (n24682 & n53012) | (n52857 & n53012);
  assign n53014 = n24355 | n24682;
  assign n53015 = n52857 | n53014;
  assign n24685 = ~n53013 & n53015;
  assign n24686 = x130 & x200;
  assign n24687 = n24685 & n24686;
  assign n24688 = n24685 | n24686;
  assign n24689 = ~n24687 & n24688;
  assign n53016 = n24362 & n24689;
  assign n53017 = (n24689 & n52862) | (n24689 & n53016) | (n52862 & n53016);
  assign n53018 = n24362 | n24689;
  assign n53019 = n52862 | n53018;
  assign n24692 = ~n53017 & n53019;
  assign n24693 = x129 & x201;
  assign n24694 = n24692 & n24693;
  assign n24695 = n24692 | n24693;
  assign n24696 = ~n24694 & n24695;
  assign n52892 = n24369 | n24371;
  assign n53020 = n24696 & n52892;
  assign n53021 = n24369 & n24696;
  assign n53022 = (n52745 & n53020) | (n52745 & n53021) | (n53020 & n53021);
  assign n53023 = n24696 | n52892;
  assign n53024 = n24369 | n24696;
  assign n53025 = (n52745 & n53023) | (n52745 & n53024) | (n53023 & n53024);
  assign n24699 = ~n53022 & n53025;
  assign n24700 = x128 & x202;
  assign n24701 = n24699 & n24700;
  assign n24702 = n24699 | n24700;
  assign n24703 = ~n24701 & n24702;
  assign n52890 = n24376 | n24378;
  assign n68348 = n24703 & n52890;
  assign n68349 = n24376 & n24703;
  assign n68350 = (n52743 & n68348) | (n52743 & n68349) | (n68348 & n68349);
  assign n68351 = n24703 | n52890;
  assign n68352 = n24376 | n24703;
  assign n68353 = (n52743 & n68351) | (n52743 & n68352) | (n68351 & n68352);
  assign n24706 = ~n68350 & n68353;
  assign n24707 = x127 & x203;
  assign n24708 = n24706 & n24707;
  assign n24709 = n24706 | n24707;
  assign n24710 = ~n24708 & n24709;
  assign n52888 = n24383 | n24385;
  assign n68354 = n24710 & n52888;
  assign n68355 = n24383 & n24710;
  assign n68356 = (n52741 & n68354) | (n52741 & n68355) | (n68354 & n68355);
  assign n68357 = n24710 | n52888;
  assign n68358 = n24383 | n24710;
  assign n68359 = (n52741 & n68357) | (n52741 & n68358) | (n68357 & n68358);
  assign n24713 = ~n68356 & n68359;
  assign n24714 = x126 & x204;
  assign n24715 = n24713 & n24714;
  assign n24716 = n24713 | n24714;
  assign n24717 = ~n24715 & n24716;
  assign n24718 = n52887 & n24717;
  assign n24719 = n52887 | n24717;
  assign n24720 = ~n24718 & n24719;
  assign n24721 = x125 & x205;
  assign n24722 = n24720 & n24721;
  assign n24723 = n24720 | n24721;
  assign n24724 = ~n24722 & n24723;
  assign n24725 = n52885 & n24724;
  assign n24726 = n52885 | n24724;
  assign n24727 = ~n24725 & n24726;
  assign n24728 = x124 & x206;
  assign n24729 = n24727 & n24728;
  assign n24730 = n24727 | n24728;
  assign n24731 = ~n24729 & n24730;
  assign n24732 = n52883 & n24731;
  assign n24733 = n52883 | n24731;
  assign n24734 = ~n24732 & n24733;
  assign n24735 = x123 & x207;
  assign n24736 = n24734 & n24735;
  assign n24737 = n24734 | n24735;
  assign n24738 = ~n24736 & n24737;
  assign n24739 = n52881 & n24738;
  assign n24740 = n52881 | n24738;
  assign n24741 = ~n24739 & n24740;
  assign n24742 = x122 & x208;
  assign n24743 = n24741 & n24742;
  assign n24744 = n24741 | n24742;
  assign n24745 = ~n24743 & n24744;
  assign n24746 = n52879 & n24745;
  assign n24747 = n52879 | n24745;
  assign n24748 = ~n24746 & n24747;
  assign n24749 = x121 & x209;
  assign n24750 = n24748 & n24749;
  assign n24751 = n24748 | n24749;
  assign n24752 = ~n24750 & n24751;
  assign n24753 = n24491 & n24752;
  assign n24754 = n24491 | n24752;
  assign n24755 = ~n24753 & n24754;
  assign n24756 = x120 & x210;
  assign n24757 = n24755 & n24756;
  assign n24758 = n24755 | n24756;
  assign n24759 = ~n24757 & n24758;
  assign n24760 = n68268 & n24759;
  assign n24761 = n68268 | n24759;
  assign n24762 = ~n24760 & n24761;
  assign n24763 = x119 & x211;
  assign n24764 = n24762 & n24763;
  assign n24765 = n24762 | n24763;
  assign n24766 = ~n24764 & n24765;
  assign n24767 = n52877 & n24766;
  assign n24768 = n52877 | n24766;
  assign n24769 = ~n24767 & n24768;
  assign n24770 = x118 & x212;
  assign n24771 = n24769 & n24770;
  assign n24772 = n24769 | n24770;
  assign n24773 = ~n24771 & n24772;
  assign n24774 = n52875 & n24773;
  assign n24775 = n52875 | n24773;
  assign n24776 = ~n24774 & n24775;
  assign n24777 = x117 & x213;
  assign n24778 = n24776 & n24777;
  assign n24779 = n24776 | n24777;
  assign n24780 = ~n24778 & n24779;
  assign n24781 = n52873 & n24780;
  assign n24782 = n52873 | n24780;
  assign n24783 = ~n24781 & n24782;
  assign n24784 = x116 & x214;
  assign n24785 = n24783 & n24784;
  assign n24786 = n24783 | n24784;
  assign n24787 = ~n24785 & n24786;
  assign n24788 = n52871 & n24787;
  assign n24789 = n52871 | n24787;
  assign n24790 = ~n24788 & n24789;
  assign n24791 = x115 & x215;
  assign n24792 = n24790 & n24791;
  assign n24793 = n24790 | n24791;
  assign n24794 = ~n24792 & n24793;
  assign n24795 = n52869 & n24794;
  assign n24796 = n52869 | n24794;
  assign n24797 = ~n24795 & n24796;
  assign n24798 = x114 & x216;
  assign n24799 = n24797 & n24798;
  assign n24800 = n24797 | n24798;
  assign n24801 = ~n24799 & n24800;
  assign n24802 = n52867 & n24801;
  assign n24803 = n52867 | n24801;
  assign n24804 = ~n24802 & n24803;
  assign n24805 = x113 & x217;
  assign n24806 = n24804 & n24805;
  assign n24807 = n24804 | n24805;
  assign n24808 = ~n24806 & n24807;
  assign n24809 = n24481 & n24808;
  assign n24810 = n24481 | n24808;
  assign n24811 = ~n24809 & n24810;
  assign n24812 = x112 & x218;
  assign n24813 = n24811 & n24812;
  assign n24814 = n24811 | n24812;
  assign n24815 = ~n24813 & n24814;
  assign n68360 = n24481 | n24805;
  assign n68361 = (n24481 & n24804) | (n24481 & n68360) | (n24804 & n68360);
  assign n53027 = (n24806 & n24808) | (n24806 & n68361) | (n24808 & n68361);
  assign n53028 = n24799 | n52867;
  assign n53029 = (n24799 & n24801) | (n24799 & n53028) | (n24801 & n53028);
  assign n53030 = n24792 | n52869;
  assign n53031 = (n24792 & n24794) | (n24792 & n53030) | (n24794 & n53030);
  assign n53032 = n24785 | n52871;
  assign n53033 = (n24785 & n24787) | (n24785 & n53032) | (n24787 & n53032);
  assign n53034 = n24778 | n52873;
  assign n53035 = (n24778 & n24780) | (n24778 & n53034) | (n24780 & n53034);
  assign n53036 = n24771 | n52875;
  assign n53037 = (n24771 & n24773) | (n24771 & n53036) | (n24773 & n53036);
  assign n53038 = n24764 | n52877;
  assign n53039 = (n24764 & n24766) | (n24764 & n53038) | (n24766 & n53038);
  assign n68362 = n24757 | n68268;
  assign n68363 = (n24757 & n24759) | (n24757 & n68362) | (n24759 & n68362);
  assign n53040 = n24750 | n24752;
  assign n53041 = (n24491 & n24750) | (n24491 & n53040) | (n24750 & n53040);
  assign n53042 = n24743 | n24745;
  assign n53043 = (n24743 & n52879) | (n24743 & n53042) | (n52879 & n53042);
  assign n53044 = n24736 | n24738;
  assign n53045 = (n24736 & n52881) | (n24736 & n53044) | (n52881 & n53044);
  assign n53046 = n24729 | n24731;
  assign n53047 = (n24729 & n52883) | (n24729 & n53046) | (n52883 & n53046);
  assign n53048 = n24722 | n24724;
  assign n53049 = (n24722 & n52885) | (n24722 & n53048) | (n52885 & n53048);
  assign n52889 = (n24383 & n52741) | (n24383 & n52888) | (n52741 & n52888);
  assign n52891 = (n24376 & n52743) | (n24376 & n52890) | (n52743 & n52890);
  assign n52896 = (n68140 & n68270) | (n68140 & n52895) | (n68270 & n52895);
  assign n53059 = n24624 | n24626;
  assign n68364 = n24299 | n24624;
  assign n68365 = (n24624 & n24626) | (n24624 & n68364) | (n24626 & n68364);
  assign n68366 = (n52823 & n53059) | (n52823 & n68365) | (n53059 & n68365);
  assign n68367 = (n52822 & n53059) | (n52822 & n68365) | (n53059 & n68365);
  assign n68368 = (n52602 & n68366) | (n52602 & n68367) | (n68366 & n68367);
  assign n53064 = n24603 | n24605;
  assign n68369 = n24278 | n24603;
  assign n68370 = (n24603 & n24605) | (n24603 & n68369) | (n24605 & n68369);
  assign n68371 = (n52813 & n53064) | (n52813 & n68370) | (n53064 & n68370);
  assign n68372 = (n52812 & n53064) | (n52812 & n68370) | (n53064 & n68370);
  assign n68373 = (n68068 & n68371) | (n68068 & n68372) | (n68371 & n68372);
  assign n52762 = (n52518 & n68171) | (n52518 & n52761) | (n68171 & n52761);
  assign n24857 = x155 & x176;
  assign n24858 = x154 & x177;
  assign n24859 = n24857 & n24858;
  assign n24860 = n24857 | n24858;
  assign n24861 = ~n24859 & n24860;
  assign n68382 = n24201 | n24526;
  assign n68383 = (n24526 & n24528) | (n24526 & n68382) | (n24528 & n68382);
  assign n53091 = n24861 & n68383;
  assign n53089 = n24526 | n24528;
  assign n53092 = n24861 & n53089;
  assign n53093 = (n68195 & n53091) | (n68195 & n53092) | (n53091 & n53092);
  assign n53094 = n24861 | n68383;
  assign n53095 = n24861 | n53089;
  assign n53096 = (n68195 & n53094) | (n68195 & n53095) | (n53094 & n53095);
  assign n24864 = ~n53093 & n53096;
  assign n24865 = x153 & x178;
  assign n24866 = n24864 & n24865;
  assign n24867 = n24864 | n24865;
  assign n24868 = ~n24866 & n24867;
  assign n68384 = n24533 | n24535;
  assign n68385 = (n24533 & n68284) | (n24533 & n68384) | (n68284 & n68384);
  assign n53097 = n24868 & n68385;
  assign n68386 = (n24533 & n68285) | (n24533 & n68384) | (n68285 & n68384);
  assign n53098 = n24868 & n68386;
  assign n68387 = (n53097 & n53098) | (n53097 & n68020) | (n53098 & n68020);
  assign n68388 = (n53097 & n53098) | (n53097 & n68019) | (n53098 & n68019);
  assign n68389 = (n67426 & n68387) | (n67426 & n68388) | (n68387 & n68388);
  assign n53100 = n24868 | n68385;
  assign n53101 = n24868 | n68386;
  assign n68390 = (n53100 & n53101) | (n53100 & n68020) | (n53101 & n68020);
  assign n68391 = (n53100 & n53101) | (n53100 & n68019) | (n53101 & n68019);
  assign n68392 = (n67426 & n68390) | (n67426 & n68391) | (n68390 & n68391);
  assign n24871 = ~n68389 & n68392;
  assign n24872 = x152 & x179;
  assign n24873 = n24871 & n24872;
  assign n24874 = n24871 | n24872;
  assign n24875 = ~n24873 & n24874;
  assign n68393 = n24540 | n24542;
  assign n68394 = (n24540 & n52919) | (n24540 & n68393) | (n52919 & n68393);
  assign n53103 = n24875 & n68394;
  assign n68395 = n24215 | n24540;
  assign n68396 = (n24540 & n24542) | (n24540 & n68395) | (n24542 & n68395);
  assign n53104 = n24875 & n68396;
  assign n68397 = (n53103 & n53104) | (n53103 & n68183) | (n53104 & n68183);
  assign n68398 = (n53103 & n53104) | (n53103 & n68184) | (n53104 & n68184);
  assign n68399 = (n67914 & n68397) | (n67914 & n68398) | (n68397 & n68398);
  assign n53106 = n24875 | n68394;
  assign n53107 = n24875 | n68396;
  assign n68400 = (n53106 & n53107) | (n53106 & n68183) | (n53107 & n68183);
  assign n68401 = (n53106 & n53107) | (n53106 & n68184) | (n53107 & n68184);
  assign n68402 = (n67914 & n68400) | (n67914 & n68401) | (n68400 & n68401);
  assign n24878 = ~n68399 & n68402;
  assign n24879 = x151 & x180;
  assign n24880 = n24878 & n24879;
  assign n24881 = n24878 | n24879;
  assign n24882 = ~n24880 & n24881;
  assign n68403 = n24547 | n24549;
  assign n68404 = (n24547 & n52917) | (n24547 & n68403) | (n52917 & n68403);
  assign n53109 = n24882 & n68404;
  assign n68405 = n24222 | n24547;
  assign n68406 = (n24547 & n24549) | (n24547 & n68405) | (n24549 & n68405);
  assign n53110 = n24882 & n68406;
  assign n68407 = (n53109 & n53110) | (n53109 & n68181) | (n53110 & n68181);
  assign n68408 = (n53109 & n53110) | (n53109 & n68180) | (n53110 & n68180);
  assign n68409 = (n67940 & n68407) | (n67940 & n68408) | (n68407 & n68408);
  assign n53112 = n24882 | n68404;
  assign n53113 = n24882 | n68406;
  assign n68410 = (n53112 & n53113) | (n53112 & n68181) | (n53113 & n68181);
  assign n68411 = (n53112 & n53113) | (n53112 & n68180) | (n53113 & n68180);
  assign n68412 = (n67940 & n68410) | (n67940 & n68411) | (n68410 & n68411);
  assign n24885 = ~n68409 & n68412;
  assign n24886 = x150 & x181;
  assign n24887 = n24885 & n24886;
  assign n24888 = n24885 | n24886;
  assign n24889 = ~n24887 & n24888;
  assign n53115 = n24554 & n24889;
  assign n53116 = (n24889 & n68308) | (n24889 & n53115) | (n68308 & n53115);
  assign n53117 = n24554 | n24889;
  assign n53118 = n68308 | n53117;
  assign n24892 = ~n53116 & n53118;
  assign n24893 = x149 & x182;
  assign n24894 = n24892 & n24893;
  assign n24895 = n24892 | n24893;
  assign n24896 = ~n24894 & n24895;
  assign n68378 = n24561 | n24563;
  assign n68379 = (n24561 & n52912) | (n24561 & n68378) | (n52912 & n68378);
  assign n68413 = n24896 & n68379;
  assign n68380 = n24236 | n24561;
  assign n68381 = (n24561 & n24563) | (n24561 & n68380) | (n24563 & n68380);
  assign n68414 = n24896 & n68381;
  assign n68415 = (n68178 & n68413) | (n68178 & n68414) | (n68413 & n68414);
  assign n68416 = n24896 | n68379;
  assign n68417 = n24896 | n68381;
  assign n68418 = (n68178 & n68416) | (n68178 & n68417) | (n68416 & n68417);
  assign n24899 = ~n68415 & n68418;
  assign n24900 = x148 & x183;
  assign n24901 = n24899 & n24900;
  assign n24902 = n24899 | n24900;
  assign n24903 = ~n24901 & n24902;
  assign n53074 = n24568 | n24570;
  assign n53119 = n24903 & n53074;
  assign n53120 = n24568 & n24903;
  assign n68419 = (n52910 & n53119) | (n52910 & n53120) | (n53119 & n53120);
  assign n68420 = (n53119 & n53120) | (n53119 & n68282) | (n53120 & n68282);
  assign n68421 = (n52615 & n68419) | (n52615 & n68420) | (n68419 & n68420);
  assign n53122 = n24903 | n53074;
  assign n53123 = n24568 | n24903;
  assign n68422 = (n52910 & n53122) | (n52910 & n53123) | (n53122 & n53123);
  assign n68423 = (n53122 & n53123) | (n53122 & n68282) | (n53123 & n68282);
  assign n68424 = (n52615 & n68422) | (n52615 & n68423) | (n68422 & n68423);
  assign n24906 = ~n68421 & n68424;
  assign n24907 = x147 & x184;
  assign n24908 = n24906 & n24907;
  assign n24909 = n24906 | n24907;
  assign n24910 = ~n24908 & n24909;
  assign n53072 = n24575 | n52958;
  assign n68425 = n24910 & n53072;
  assign n68376 = n24250 | n24575;
  assign n68377 = (n24575 & n24577) | (n24575 & n68376) | (n24577 & n68376);
  assign n68426 = n24910 & n68377;
  assign n68427 = (n52762 & n68425) | (n52762 & n68426) | (n68425 & n68426);
  assign n68428 = n24910 | n53072;
  assign n68429 = n24910 | n68377;
  assign n68430 = (n52762 & n68428) | (n52762 & n68429) | (n68428 & n68429);
  assign n24913 = ~n68427 & n68430;
  assign n24914 = x146 & x185;
  assign n24915 = n24913 & n24914;
  assign n24916 = n24913 | n24914;
  assign n24917 = ~n24915 & n24916;
  assign n53069 = n24582 | n24584;
  assign n68431 = n24917 & n53069;
  assign n68374 = n24257 | n24582;
  assign n68375 = (n24582 & n24584) | (n24582 & n68374) | (n24584 & n68374);
  assign n68432 = n24917 & n68375;
  assign n68433 = (n52804 & n68431) | (n52804 & n68432) | (n68431 & n68432);
  assign n68434 = n24917 | n53069;
  assign n68435 = n24917 | n68375;
  assign n68436 = (n52804 & n68434) | (n52804 & n68435) | (n68434 & n68435);
  assign n24920 = ~n68433 & n68436;
  assign n24921 = x145 & x186;
  assign n24922 = n24920 & n24921;
  assign n24923 = n24920 | n24921;
  assign n24924 = ~n24922 & n24923;
  assign n53066 = n24589 | n24591;
  assign n53125 = n24924 & n53066;
  assign n53126 = n24589 & n24924;
  assign n53127 = (n68280 & n53125) | (n68280 & n53126) | (n53125 & n53126);
  assign n53128 = n24924 | n53066;
  assign n53129 = n24589 | n24924;
  assign n53130 = (n68280 & n53128) | (n68280 & n53129) | (n53128 & n53129);
  assign n24927 = ~n53127 & n53130;
  assign n24928 = x144 & x187;
  assign n24929 = n24927 & n24928;
  assign n24930 = n24927 | n24928;
  assign n24931 = ~n24929 & n24930;
  assign n53131 = n24596 & n24931;
  assign n68437 = (n24931 & n52969) | (n24931 & n53131) | (n52969 & n53131);
  assign n68438 = (n24931 & n52968) | (n24931 & n53131) | (n52968 & n53131);
  assign n68439 = (n68169 & n68437) | (n68169 & n68438) | (n68437 & n68438);
  assign n53133 = n24596 | n24931;
  assign n68440 = n52969 | n53133;
  assign n68441 = n52968 | n53133;
  assign n68442 = (n68169 & n68440) | (n68169 & n68441) | (n68440 & n68441);
  assign n24934 = ~n68439 & n68442;
  assign n24935 = x143 & x188;
  assign n24936 = n24934 & n24935;
  assign n24937 = n24934 | n24935;
  assign n24938 = ~n24936 & n24937;
  assign n24939 = n68373 & n24938;
  assign n24940 = n68373 | n24938;
  assign n24941 = ~n24939 & n24940;
  assign n24942 = x142 & x189;
  assign n24943 = n24941 & n24942;
  assign n24944 = n24941 | n24942;
  assign n24945 = ~n24943 & n24944;
  assign n53061 = n24610 | n24612;
  assign n53135 = n24945 & n53061;
  assign n53136 = n24610 & n24945;
  assign n53137 = (n68275 & n53135) | (n68275 & n53136) | (n53135 & n53136);
  assign n53138 = n24945 | n53061;
  assign n53139 = n24610 | n24945;
  assign n53140 = (n68275 & n53138) | (n68275 & n53139) | (n53138 & n53139);
  assign n24948 = ~n53137 & n53140;
  assign n24949 = x141 & x190;
  assign n24950 = n24948 & n24949;
  assign n24951 = n24948 | n24949;
  assign n24952 = ~n24950 & n24951;
  assign n53141 = n24617 & n24952;
  assign n68443 = (n24952 & n52979) | (n24952 & n53141) | (n52979 & n53141);
  assign n68444 = (n24952 & n52978) | (n24952 & n53141) | (n52978 & n53141);
  assign n68445 = (n68164 & n68443) | (n68164 & n68444) | (n68443 & n68444);
  assign n53143 = n24617 | n24952;
  assign n68446 = n52979 | n53143;
  assign n68447 = n52978 | n53143;
  assign n68448 = (n68164 & n68446) | (n68164 & n68447) | (n68446 & n68447);
  assign n24955 = ~n68445 & n68448;
  assign n24956 = x140 & x191;
  assign n24957 = n24955 & n24956;
  assign n24958 = n24955 | n24956;
  assign n24959 = ~n24957 & n24958;
  assign n24960 = n68368 & n24959;
  assign n24961 = n68368 | n24959;
  assign n24962 = ~n24960 & n24961;
  assign n24963 = x139 & x192;
  assign n24964 = n24962 & n24963;
  assign n24965 = n24962 | n24963;
  assign n24966 = ~n24964 & n24965;
  assign n53056 = n24631 | n24633;
  assign n53145 = n24966 & n53056;
  assign n53146 = n24631 & n24966;
  assign n53147 = (n52896 & n53145) | (n52896 & n53146) | (n53145 & n53146);
  assign n53148 = n24966 | n53056;
  assign n53149 = n24631 | n24966;
  assign n53150 = (n52896 & n53148) | (n52896 & n53149) | (n53148 & n53149);
  assign n24969 = ~n53147 & n53150;
  assign n24970 = x138 & x193;
  assign n24971 = n24969 & n24970;
  assign n24972 = n24969 | n24970;
  assign n24973 = ~n24971 & n24972;
  assign n53151 = n24638 & n24973;
  assign n53152 = (n24973 & n68344) | (n24973 & n53151) | (n68344 & n53151);
  assign n53153 = n24638 | n24973;
  assign n53154 = n68344 | n53153;
  assign n24976 = ~n53152 & n53154;
  assign n24977 = x137 & x194;
  assign n24978 = n24976 & n24977;
  assign n24979 = n24976 | n24977;
  assign n24980 = ~n24978 & n24979;
  assign n53155 = n24645 & n24980;
  assign n53156 = (n24980 & n52993) | (n24980 & n53155) | (n52993 & n53155);
  assign n53157 = n24645 | n24980;
  assign n53158 = n52993 | n53157;
  assign n24983 = ~n53156 & n53158;
  assign n24984 = x136 & x195;
  assign n24985 = n24983 & n24984;
  assign n24986 = n24983 | n24984;
  assign n24987 = ~n24985 & n24986;
  assign n53159 = n24652 & n24987;
  assign n53160 = (n24987 & n52997) | (n24987 & n53159) | (n52997 & n53159);
  assign n53161 = n24652 | n24987;
  assign n53162 = n52997 | n53161;
  assign n24990 = ~n53160 & n53162;
  assign n24991 = x135 & x196;
  assign n24992 = n24990 & n24991;
  assign n24993 = n24990 | n24991;
  assign n24994 = ~n24992 & n24993;
  assign n53163 = n24659 & n24994;
  assign n53164 = (n24994 & n53001) | (n24994 & n53163) | (n53001 & n53163);
  assign n53165 = n24659 | n24994;
  assign n53166 = n53001 | n53165;
  assign n24997 = ~n53164 & n53166;
  assign n24998 = x134 & x197;
  assign n24999 = n24997 & n24998;
  assign n25000 = n24997 | n24998;
  assign n25001 = ~n24999 & n25000;
  assign n53167 = n24666 & n25001;
  assign n53168 = (n25001 & n53005) | (n25001 & n53167) | (n53005 & n53167);
  assign n53169 = n24666 | n25001;
  assign n53170 = n53005 | n53169;
  assign n25004 = ~n53168 & n53170;
  assign n25005 = x133 & x198;
  assign n25006 = n25004 & n25005;
  assign n25007 = n25004 | n25005;
  assign n25008 = ~n25006 & n25007;
  assign n53171 = n24673 & n25008;
  assign n53172 = (n25008 & n53009) | (n25008 & n53171) | (n53009 & n53171);
  assign n53173 = n24673 | n25008;
  assign n53174 = n53009 | n53173;
  assign n25011 = ~n53172 & n53174;
  assign n25012 = x132 & x199;
  assign n25013 = n25011 & n25012;
  assign n25014 = n25011 | n25012;
  assign n25015 = ~n25013 & n25014;
  assign n53175 = n24680 & n25015;
  assign n53176 = (n25015 & n53013) | (n25015 & n53175) | (n53013 & n53175);
  assign n53177 = n24680 | n25015;
  assign n53178 = n53013 | n53177;
  assign n25018 = ~n53176 & n53178;
  assign n25019 = x131 & x200;
  assign n25020 = n25018 & n25019;
  assign n25021 = n25018 | n25019;
  assign n25022 = ~n25020 & n25021;
  assign n53179 = n24687 & n25022;
  assign n53180 = (n25022 & n53017) | (n25022 & n53179) | (n53017 & n53179);
  assign n53181 = n24687 | n25022;
  assign n53182 = n53017 | n53181;
  assign n25025 = ~n53180 & n53182;
  assign n25026 = x130 & x201;
  assign n25027 = n25025 & n25026;
  assign n25028 = n25025 | n25026;
  assign n25029 = ~n25027 & n25028;
  assign n53183 = n24694 & n25029;
  assign n53184 = (n25029 & n53022) | (n25029 & n53183) | (n53022 & n53183);
  assign n53185 = n24694 | n25029;
  assign n53186 = n53022 | n53185;
  assign n25032 = ~n53184 & n53186;
  assign n25033 = x129 & x202;
  assign n25034 = n25032 & n25033;
  assign n25035 = n25032 | n25033;
  assign n25036 = ~n25034 & n25035;
  assign n53054 = n24701 | n24703;
  assign n53187 = n25036 & n53054;
  assign n53188 = n24701 & n25036;
  assign n53189 = (n52891 & n53187) | (n52891 & n53188) | (n53187 & n53188);
  assign n53190 = n25036 | n53054;
  assign n53191 = n24701 | n25036;
  assign n53192 = (n52891 & n53190) | (n52891 & n53191) | (n53190 & n53191);
  assign n25039 = ~n53189 & n53192;
  assign n25040 = x128 & x203;
  assign n25041 = n25039 & n25040;
  assign n25042 = n25039 | n25040;
  assign n25043 = ~n25041 & n25042;
  assign n53052 = n24708 | n24710;
  assign n68449 = n25043 & n53052;
  assign n68450 = n24708 & n25043;
  assign n68451 = (n52889 & n68449) | (n52889 & n68450) | (n68449 & n68450);
  assign n68452 = n25043 | n53052;
  assign n68453 = n24708 | n25043;
  assign n68454 = (n52889 & n68452) | (n52889 & n68453) | (n68452 & n68453);
  assign n25046 = ~n68451 & n68454;
  assign n25047 = x127 & x204;
  assign n25048 = n25046 & n25047;
  assign n25049 = n25046 | n25047;
  assign n25050 = ~n25048 & n25049;
  assign n53050 = n24715 | n24717;
  assign n68455 = n25050 & n53050;
  assign n68456 = n24715 & n25050;
  assign n68457 = (n52887 & n68455) | (n52887 & n68456) | (n68455 & n68456);
  assign n68458 = n25050 | n53050;
  assign n68459 = n24715 | n25050;
  assign n68460 = (n52887 & n68458) | (n52887 & n68459) | (n68458 & n68459);
  assign n25053 = ~n68457 & n68460;
  assign n25054 = x126 & x205;
  assign n25055 = n25053 & n25054;
  assign n25056 = n25053 | n25054;
  assign n25057 = ~n25055 & n25056;
  assign n25058 = n53049 & n25057;
  assign n25059 = n53049 | n25057;
  assign n25060 = ~n25058 & n25059;
  assign n25061 = x125 & x206;
  assign n25062 = n25060 & n25061;
  assign n25063 = n25060 | n25061;
  assign n25064 = ~n25062 & n25063;
  assign n25065 = n53047 & n25064;
  assign n25066 = n53047 | n25064;
  assign n25067 = ~n25065 & n25066;
  assign n25068 = x124 & x207;
  assign n25069 = n25067 & n25068;
  assign n25070 = n25067 | n25068;
  assign n25071 = ~n25069 & n25070;
  assign n25072 = n53045 & n25071;
  assign n25073 = n53045 | n25071;
  assign n25074 = ~n25072 & n25073;
  assign n25075 = x123 & x208;
  assign n25076 = n25074 & n25075;
  assign n25077 = n25074 | n25075;
  assign n25078 = ~n25076 & n25077;
  assign n25079 = n53043 & n25078;
  assign n25080 = n53043 | n25078;
  assign n25081 = ~n25079 & n25080;
  assign n25082 = x122 & x209;
  assign n25083 = n25081 & n25082;
  assign n25084 = n25081 | n25082;
  assign n25085 = ~n25083 & n25084;
  assign n25086 = n53041 & n25085;
  assign n25087 = n53041 | n25085;
  assign n25088 = ~n25086 & n25087;
  assign n25089 = x121 & x210;
  assign n25090 = n25088 & n25089;
  assign n25091 = n25088 | n25089;
  assign n25092 = ~n25090 & n25091;
  assign n25093 = n68363 & n25092;
  assign n25094 = n68363 | n25092;
  assign n25095 = ~n25093 & n25094;
  assign n25096 = x120 & x211;
  assign n25097 = n25095 & n25096;
  assign n25098 = n25095 | n25096;
  assign n25099 = ~n25097 & n25098;
  assign n25100 = n53039 & n25099;
  assign n25101 = n53039 | n25099;
  assign n25102 = ~n25100 & n25101;
  assign n25103 = x119 & x212;
  assign n25104 = n25102 & n25103;
  assign n25105 = n25102 | n25103;
  assign n25106 = ~n25104 & n25105;
  assign n25107 = n53037 & n25106;
  assign n25108 = n53037 | n25106;
  assign n25109 = ~n25107 & n25108;
  assign n25110 = x118 & x213;
  assign n25111 = n25109 & n25110;
  assign n25112 = n25109 | n25110;
  assign n25113 = ~n25111 & n25112;
  assign n25114 = n53035 & n25113;
  assign n25115 = n53035 | n25113;
  assign n25116 = ~n25114 & n25115;
  assign n25117 = x117 & x214;
  assign n25118 = n25116 & n25117;
  assign n25119 = n25116 | n25117;
  assign n25120 = ~n25118 & n25119;
  assign n25121 = n53033 & n25120;
  assign n25122 = n53033 | n25120;
  assign n25123 = ~n25121 & n25122;
  assign n25124 = x116 & x215;
  assign n25125 = n25123 & n25124;
  assign n25126 = n25123 | n25124;
  assign n25127 = ~n25125 & n25126;
  assign n25128 = n53031 & n25127;
  assign n25129 = n53031 | n25127;
  assign n25130 = ~n25128 & n25129;
  assign n25131 = x115 & x216;
  assign n25132 = n25130 & n25131;
  assign n25133 = n25130 | n25131;
  assign n25134 = ~n25132 & n25133;
  assign n25135 = n53029 & n25134;
  assign n25136 = n53029 | n25134;
  assign n25137 = ~n25135 & n25136;
  assign n25138 = x114 & x217;
  assign n25139 = n25137 & n25138;
  assign n25140 = n25137 | n25138;
  assign n25141 = ~n25139 & n25140;
  assign n25142 = n53027 & n25141;
  assign n25143 = n53027 | n25141;
  assign n25144 = ~n25142 & n25143;
  assign n25145 = x113 & x218;
  assign n25146 = n25144 & n25145;
  assign n25147 = n25144 | n25145;
  assign n25148 = ~n25146 & n25147;
  assign n25149 = n24813 & n25148;
  assign n25150 = n24813 | n25148;
  assign n25151 = ~n25149 & n25150;
  assign n25152 = x112 & x219;
  assign n25153 = n25151 & n25152;
  assign n25154 = n25151 | n25152;
  assign n25155 = ~n25153 & n25154;
  assign n53193 = n24813 | n25146;
  assign n53194 = (n25146 & n25148) | (n25146 & n53193) | (n25148 & n53193);
  assign n53195 = n25139 | n53027;
  assign n53196 = (n25139 & n25141) | (n25139 & n53195) | (n25141 & n53195);
  assign n53197 = n25132 | n53029;
  assign n53198 = (n25132 & n25134) | (n25132 & n53197) | (n25134 & n53197);
  assign n53199 = n25125 | n53031;
  assign n53200 = (n25125 & n25127) | (n25125 & n53199) | (n25127 & n53199);
  assign n53201 = n25118 | n53033;
  assign n53202 = (n25118 & n25120) | (n25118 & n53201) | (n25120 & n53201);
  assign n53203 = n25111 | n53035;
  assign n53204 = (n25111 & n25113) | (n25111 & n53203) | (n25113 & n53203);
  assign n53205 = n25104 | n53037;
  assign n53206 = (n25104 & n25106) | (n25104 & n53205) | (n25106 & n53205);
  assign n53207 = n25097 | n53039;
  assign n53208 = (n25097 & n25099) | (n25097 & n53207) | (n25099 & n53207);
  assign n53209 = n25090 | n25092;
  assign n53210 = (n68363 & n25090) | (n68363 & n53209) | (n25090 & n53209);
  assign n53211 = n25083 | n25085;
  assign n53212 = (n25083 & n53041) | (n25083 & n53211) | (n53041 & n53211);
  assign n53213 = n25076 | n25078;
  assign n53214 = (n25076 & n53043) | (n25076 & n53213) | (n53043 & n53213);
  assign n53215 = n25069 | n25071;
  assign n53216 = (n25069 & n53045) | (n25069 & n53215) | (n53045 & n53215);
  assign n53217 = n25062 | n25064;
  assign n53218 = (n25062 & n53047) | (n25062 & n53217) | (n53047 & n53217);
  assign n53051 = (n24715 & n52887) | (n24715 & n53050) | (n52887 & n53050);
  assign n53053 = (n24708 & n52889) | (n24708 & n53052) | (n52889 & n53052);
  assign n53231 = n24950 | n24952;
  assign n68463 = n24617 | n24950;
  assign n68464 = (n24950 & n24952) | (n24950 & n68463) | (n24952 & n68463);
  assign n68465 = (n52979 & n53231) | (n52979 & n68464) | (n53231 & n68464);
  assign n68466 = (n52978 & n53231) | (n52978 & n68464) | (n53231 & n68464);
  assign n68467 = (n68164 & n68465) | (n68164 & n68466) | (n68465 & n68466);
  assign n53236 = n24929 | n24931;
  assign n68468 = n24596 | n24929;
  assign n68469 = (n24929 & n24931) | (n24929 & n68468) | (n24931 & n68468);
  assign n68470 = (n52969 & n53236) | (n52969 & n68469) | (n53236 & n68469);
  assign n68471 = (n52968 & n53236) | (n52968 & n68469) | (n53236 & n68469);
  assign n68472 = (n68169 & n68470) | (n68169 & n68471) | (n68470 & n68471);
  assign n53070 = (n52804 & n68375) | (n52804 & n53069) | (n68375 & n53069);
  assign n68473 = n24568 | n24901;
  assign n68474 = (n24901 & n24903) | (n24901 & n68473) | (n24903 & n68473);
  assign n68475 = n24901 | n24903;
  assign n68476 = (n24901 & n53074) | (n24901 & n68475) | (n53074 & n68475);
  assign n68477 = (n52910 & n68474) | (n52910 & n68476) | (n68474 & n68476);
  assign n68478 = (n68282 & n68474) | (n68282 & n68476) | (n68474 & n68476);
  assign n68479 = (n52615 & n68477) | (n52615 & n68478) | (n68477 & n68478);
  assign n25198 = x156 & x176;
  assign n25199 = x155 & x177;
  assign n25200 = n25198 & n25199;
  assign n25201 = n25198 | n25199;
  assign n25202 = ~n25200 & n25201;
  assign n68486 = n24859 | n24861;
  assign n68487 = (n24859 & n68383) | (n24859 & n68486) | (n68383 & n68486);
  assign n53256 = n25202 & n68487;
  assign n68488 = (n24859 & n53089) | (n24859 & n68486) | (n53089 & n68486);
  assign n53257 = n25202 & n68488;
  assign n53258 = (n68195 & n53256) | (n68195 & n53257) | (n53256 & n53257);
  assign n53259 = n25202 | n68487;
  assign n53260 = n25202 | n68488;
  assign n53261 = (n68195 & n53259) | (n68195 & n53260) | (n53259 & n53260);
  assign n25205 = ~n53258 & n53261;
  assign n25206 = x154 & x178;
  assign n25207 = n25205 & n25206;
  assign n25208 = n25205 | n25206;
  assign n25209 = ~n25207 & n25208;
  assign n53262 = n24866 & n25209;
  assign n53263 = (n25209 & n68389) | (n25209 & n53262) | (n68389 & n53262);
  assign n53264 = n24866 | n25209;
  assign n53265 = n68389 | n53264;
  assign n25212 = ~n53263 & n53265;
  assign n25213 = x153 & x179;
  assign n25214 = n25212 & n25213;
  assign n25215 = n25212 | n25213;
  assign n25216 = ~n25214 & n25215;
  assign n68480 = n24873 | n24875;
  assign n68481 = (n24873 & n68394) | (n24873 & n68480) | (n68394 & n68480);
  assign n68482 = (n24873 & n68396) | (n24873 & n68480) | (n68396 & n68480);
  assign n68484 = (n68184 & n68481) | (n68184 & n68482) | (n68481 & n68482);
  assign n68489 = n25216 & n68484;
  assign n68483 = (n68183 & n68481) | (n68183 & n68482) | (n68481 & n68482);
  assign n68490 = n25216 & n68483;
  assign n68491 = (n67914 & n68489) | (n67914 & n68490) | (n68489 & n68490);
  assign n68492 = n25216 | n68484;
  assign n68493 = n25216 | n68483;
  assign n68494 = (n67914 & n68492) | (n67914 & n68493) | (n68492 & n68493);
  assign n25219 = ~n68491 & n68494;
  assign n25220 = x152 & x180;
  assign n25221 = n25219 & n25220;
  assign n25222 = n25219 | n25220;
  assign n25223 = ~n25221 & n25222;
  assign n53266 = n24880 & n25223;
  assign n53267 = (n25223 & n68409) | (n25223 & n53266) | (n68409 & n53266);
  assign n53268 = n24880 | n25223;
  assign n53269 = n68409 | n53268;
  assign n25226 = ~n53267 & n53269;
  assign n25227 = x151 & x181;
  assign n25228 = n25226 & n25227;
  assign n25229 = n25226 | n25227;
  assign n25230 = ~n25228 & n25229;
  assign n68495 = n24554 | n24887;
  assign n68496 = (n24887 & n24889) | (n24887 & n68495) | (n24889 & n68495);
  assign n53270 = n25230 & n68496;
  assign n53248 = n24887 | n24889;
  assign n53271 = n25230 & n53248;
  assign n53272 = (n68308 & n53270) | (n68308 & n53271) | (n53270 & n53271);
  assign n53273 = n25230 | n68496;
  assign n53274 = n25230 | n53248;
  assign n53275 = (n68308 & n53273) | (n68308 & n53274) | (n53273 & n53274);
  assign n25233 = ~n53272 & n53275;
  assign n25234 = x150 & x182;
  assign n25235 = n25233 & n25234;
  assign n25236 = n25233 | n25234;
  assign n25237 = ~n25235 & n25236;
  assign n53245 = n24894 | n24896;
  assign n53276 = n25237 & n53245;
  assign n53277 = n24894 & n25237;
  assign n68497 = (n53276 & n53277) | (n53276 & n68379) | (n53277 & n68379);
  assign n68498 = (n53276 & n53277) | (n53276 & n68381) | (n53277 & n68381);
  assign n68499 = (n68178 & n68497) | (n68178 & n68498) | (n68497 & n68498);
  assign n53279 = n25237 | n53245;
  assign n53280 = n24894 | n25237;
  assign n68500 = (n53279 & n53280) | (n53279 & n68379) | (n53280 & n68379);
  assign n68501 = (n53279 & n53280) | (n53279 & n68381) | (n53280 & n68381);
  assign n68502 = (n68178 & n68500) | (n68178 & n68501) | (n68500 & n68501);
  assign n25240 = ~n68499 & n68502;
  assign n25241 = x149 & x183;
  assign n25242 = n25240 & n25241;
  assign n25243 = n25240 | n25241;
  assign n25244 = ~n25242 & n25243;
  assign n25245 = n68479 & n25244;
  assign n25246 = n68479 | n25244;
  assign n25247 = ~n25245 & n25246;
  assign n25248 = x148 & x184;
  assign n25249 = n25247 & n25248;
  assign n25250 = n25247 | n25248;
  assign n25251 = ~n25249 & n25250;
  assign n53240 = n24908 | n24910;
  assign n53282 = n25251 & n53240;
  assign n53283 = n24908 & n25251;
  assign n68503 = (n53072 & n53282) | (n53072 & n53283) | (n53282 & n53283);
  assign n68504 = (n53282 & n53283) | (n53282 & n68377) | (n53283 & n68377);
  assign n68505 = (n52762 & n68503) | (n52762 & n68504) | (n68503 & n68504);
  assign n53285 = n25251 | n53240;
  assign n53286 = n24908 | n25251;
  assign n68506 = (n53072 & n53285) | (n53072 & n53286) | (n53285 & n53286);
  assign n68507 = (n53285 & n53286) | (n53285 & n68377) | (n53286 & n68377);
  assign n68508 = (n52762 & n68506) | (n52762 & n68507) | (n68506 & n68507);
  assign n25254 = ~n68505 & n68508;
  assign n25255 = x147 & x185;
  assign n25256 = n25254 & n25255;
  assign n25257 = n25254 | n25255;
  assign n25258 = ~n25256 & n25257;
  assign n53238 = n24915 | n24917;
  assign n53288 = n25258 & n53238;
  assign n53289 = n24915 & n25258;
  assign n53290 = (n53070 & n53288) | (n53070 & n53289) | (n53288 & n53289);
  assign n53291 = n25258 | n53238;
  assign n53292 = n24915 | n25258;
  assign n53293 = (n53070 & n53291) | (n53070 & n53292) | (n53291 & n53292);
  assign n25261 = ~n53290 & n53293;
  assign n25262 = x146 & x186;
  assign n25263 = n25261 & n25262;
  assign n25264 = n25261 | n25262;
  assign n25265 = ~n25263 & n25264;
  assign n53294 = n24922 & n25265;
  assign n53295 = (n25265 & n53127) | (n25265 & n53294) | (n53127 & n53294);
  assign n53296 = n24922 | n25265;
  assign n53297 = n53127 | n53296;
  assign n25268 = ~n53295 & n53297;
  assign n25269 = x145 & x187;
  assign n25270 = n25268 & n25269;
  assign n25271 = n25268 | n25269;
  assign n25272 = ~n25270 & n25271;
  assign n25273 = n68472 & n25272;
  assign n25274 = n68472 | n25272;
  assign n25275 = ~n25273 & n25274;
  assign n25276 = x144 & x188;
  assign n25277 = n25275 & n25276;
  assign n25278 = n25275 | n25276;
  assign n25279 = ~n25277 & n25278;
  assign n53233 = n24936 | n24938;
  assign n53298 = n25279 & n53233;
  assign n53299 = n24936 & n25279;
  assign n53300 = (n68373 & n53298) | (n68373 & n53299) | (n53298 & n53299);
  assign n53301 = n25279 | n53233;
  assign n53302 = n24936 | n25279;
  assign n53303 = (n68373 & n53301) | (n68373 & n53302) | (n53301 & n53302);
  assign n25282 = ~n53300 & n53303;
  assign n25283 = x143 & x189;
  assign n25284 = n25282 & n25283;
  assign n25285 = n25282 | n25283;
  assign n25286 = ~n25284 & n25285;
  assign n53304 = n24943 & n25286;
  assign n68509 = (n25286 & n53136) | (n25286 & n53304) | (n53136 & n53304);
  assign n68510 = (n25286 & n53135) | (n25286 & n53304) | (n53135 & n53304);
  assign n68511 = (n68275 & n68509) | (n68275 & n68510) | (n68509 & n68510);
  assign n53306 = n24943 | n25286;
  assign n68512 = n53136 | n53306;
  assign n68513 = n53135 | n53306;
  assign n68514 = (n68275 & n68512) | (n68275 & n68513) | (n68512 & n68513);
  assign n25289 = ~n68511 & n68514;
  assign n25290 = x142 & x190;
  assign n25291 = n25289 & n25290;
  assign n25292 = n25289 | n25290;
  assign n25293 = ~n25291 & n25292;
  assign n25294 = n68467 & n25293;
  assign n25295 = n68467 | n25293;
  assign n25296 = ~n25294 & n25295;
  assign n25297 = x141 & x191;
  assign n25298 = n25296 & n25297;
  assign n25299 = n25296 | n25297;
  assign n25300 = ~n25298 & n25299;
  assign n53228 = n24957 | n24959;
  assign n53308 = n25300 & n53228;
  assign n53309 = n24957 & n25300;
  assign n53310 = (n68368 & n53308) | (n68368 & n53309) | (n53308 & n53309);
  assign n53311 = n25300 | n53228;
  assign n53312 = n24957 | n25300;
  assign n53313 = (n68368 & n53311) | (n68368 & n53312) | (n53311 & n53312);
  assign n25303 = ~n53310 & n53313;
  assign n25304 = x140 & x192;
  assign n25305 = n25303 & n25304;
  assign n25306 = n25303 | n25304;
  assign n25307 = ~n25305 & n25306;
  assign n53314 = n24964 & n25307;
  assign n68515 = (n25307 & n53146) | (n25307 & n53314) | (n53146 & n53314);
  assign n68516 = (n25307 & n53145) | (n25307 & n53314) | (n53145 & n53314);
  assign n68517 = (n52896 & n68515) | (n52896 & n68516) | (n68515 & n68516);
  assign n53316 = n24964 | n25307;
  assign n68518 = n53146 | n53316;
  assign n68519 = n53145 | n53316;
  assign n68520 = (n52896 & n68518) | (n52896 & n68519) | (n68518 & n68519);
  assign n25310 = ~n68517 & n68520;
  assign n25311 = x139 & x193;
  assign n25312 = n25310 & n25311;
  assign n25313 = n25310 | n25311;
  assign n25314 = ~n25312 & n25313;
  assign n53226 = n24971 | n24973;
  assign n68521 = n25314 & n53226;
  assign n68461 = n24638 | n24971;
  assign n68462 = (n24971 & n24973) | (n24971 & n68461) | (n24973 & n68461);
  assign n68522 = n25314 & n68462;
  assign n68523 = (n68344 & n68521) | (n68344 & n68522) | (n68521 & n68522);
  assign n68524 = n25314 | n53226;
  assign n68525 = n25314 | n68462;
  assign n68526 = (n68344 & n68524) | (n68344 & n68525) | (n68524 & n68525);
  assign n25317 = ~n68523 & n68526;
  assign n25318 = x138 & x194;
  assign n25319 = n25317 & n25318;
  assign n25320 = n25317 | n25318;
  assign n25321 = ~n25319 & n25320;
  assign n53318 = n24978 & n25321;
  assign n68527 = (n25321 & n53155) | (n25321 & n53318) | (n53155 & n53318);
  assign n68528 = (n24980 & n25321) | (n24980 & n53318) | (n25321 & n53318);
  assign n68529 = (n52993 & n68527) | (n52993 & n68528) | (n68527 & n68528);
  assign n53320 = n24978 | n25321;
  assign n68530 = n53155 | n53320;
  assign n68531 = n24980 | n53320;
  assign n68532 = (n52993 & n68530) | (n52993 & n68531) | (n68530 & n68531);
  assign n25324 = ~n68529 & n68532;
  assign n25325 = x137 & x195;
  assign n25326 = n25324 & n25325;
  assign n25327 = n25324 | n25325;
  assign n25328 = ~n25326 & n25327;
  assign n53322 = n24985 & n25328;
  assign n53323 = (n25328 & n53160) | (n25328 & n53322) | (n53160 & n53322);
  assign n53324 = n24985 | n25328;
  assign n53325 = n53160 | n53324;
  assign n25331 = ~n53323 & n53325;
  assign n25332 = x136 & x196;
  assign n25333 = n25331 & n25332;
  assign n25334 = n25331 | n25332;
  assign n25335 = ~n25333 & n25334;
  assign n53326 = n24992 & n25335;
  assign n53327 = (n25335 & n53164) | (n25335 & n53326) | (n53164 & n53326);
  assign n53328 = n24992 | n25335;
  assign n53329 = n53164 | n53328;
  assign n25338 = ~n53327 & n53329;
  assign n25339 = x135 & x197;
  assign n25340 = n25338 & n25339;
  assign n25341 = n25338 | n25339;
  assign n25342 = ~n25340 & n25341;
  assign n53330 = n24999 & n25342;
  assign n53331 = (n25342 & n53168) | (n25342 & n53330) | (n53168 & n53330);
  assign n53332 = n24999 | n25342;
  assign n53333 = n53168 | n53332;
  assign n25345 = ~n53331 & n53333;
  assign n25346 = x134 & x198;
  assign n25347 = n25345 & n25346;
  assign n25348 = n25345 | n25346;
  assign n25349 = ~n25347 & n25348;
  assign n53334 = n25006 & n25349;
  assign n53335 = (n25349 & n53172) | (n25349 & n53334) | (n53172 & n53334);
  assign n53336 = n25006 | n25349;
  assign n53337 = n53172 | n53336;
  assign n25352 = ~n53335 & n53337;
  assign n25353 = x133 & x199;
  assign n25354 = n25352 & n25353;
  assign n25355 = n25352 | n25353;
  assign n25356 = ~n25354 & n25355;
  assign n53338 = n25013 & n25356;
  assign n53339 = (n25356 & n53176) | (n25356 & n53338) | (n53176 & n53338);
  assign n53340 = n25013 | n25356;
  assign n53341 = n53176 | n53340;
  assign n25359 = ~n53339 & n53341;
  assign n25360 = x132 & x200;
  assign n25361 = n25359 & n25360;
  assign n25362 = n25359 | n25360;
  assign n25363 = ~n25361 & n25362;
  assign n53342 = n25020 & n25363;
  assign n53343 = (n25363 & n53180) | (n25363 & n53342) | (n53180 & n53342);
  assign n53344 = n25020 | n25363;
  assign n53345 = n53180 | n53344;
  assign n25366 = ~n53343 & n53345;
  assign n25367 = x131 & x201;
  assign n25368 = n25366 & n25367;
  assign n25369 = n25366 | n25367;
  assign n25370 = ~n25368 & n25369;
  assign n53346 = n25027 & n25370;
  assign n53347 = (n25370 & n53184) | (n25370 & n53346) | (n53184 & n53346);
  assign n53348 = n25027 | n25370;
  assign n53349 = n53184 | n53348;
  assign n25373 = ~n53347 & n53349;
  assign n25374 = x130 & x202;
  assign n25375 = n25373 & n25374;
  assign n25376 = n25373 | n25374;
  assign n25377 = ~n25375 & n25376;
  assign n53350 = n25034 & n25377;
  assign n53351 = (n25377 & n53189) | (n25377 & n53350) | (n53189 & n53350);
  assign n53352 = n25034 | n25377;
  assign n53353 = n53189 | n53352;
  assign n25380 = ~n53351 & n53353;
  assign n25381 = x129 & x203;
  assign n25382 = n25380 & n25381;
  assign n25383 = n25380 | n25381;
  assign n25384 = ~n25382 & n25383;
  assign n53223 = n25041 | n25043;
  assign n53354 = n25384 & n53223;
  assign n53355 = n25041 & n25384;
  assign n53356 = (n53053 & n53354) | (n53053 & n53355) | (n53354 & n53355);
  assign n53357 = n25384 | n53223;
  assign n53358 = n25041 | n25384;
  assign n53359 = (n53053 & n53357) | (n53053 & n53358) | (n53357 & n53358);
  assign n25387 = ~n53356 & n53359;
  assign n25388 = x128 & x204;
  assign n25389 = n25387 & n25388;
  assign n25390 = n25387 | n25388;
  assign n25391 = ~n25389 & n25390;
  assign n53221 = n25048 | n25050;
  assign n68533 = n25391 & n53221;
  assign n68534 = n25048 & n25391;
  assign n68535 = (n53051 & n68533) | (n53051 & n68534) | (n68533 & n68534);
  assign n68536 = n25391 | n53221;
  assign n68537 = n25048 | n25391;
  assign n68538 = (n53051 & n68536) | (n53051 & n68537) | (n68536 & n68537);
  assign n25394 = ~n68535 & n68538;
  assign n25395 = x127 & x205;
  assign n25396 = n25394 & n25395;
  assign n25397 = n25394 | n25395;
  assign n25398 = ~n25396 & n25397;
  assign n53219 = n25055 | n25057;
  assign n68539 = n25398 & n53219;
  assign n68540 = n25055 & n25398;
  assign n68541 = (n53049 & n68539) | (n53049 & n68540) | (n68539 & n68540);
  assign n68542 = n25398 | n53219;
  assign n68543 = n25055 | n25398;
  assign n68544 = (n53049 & n68542) | (n53049 & n68543) | (n68542 & n68543);
  assign n25401 = ~n68541 & n68544;
  assign n25402 = x126 & x206;
  assign n25403 = n25401 & n25402;
  assign n25404 = n25401 | n25402;
  assign n25405 = ~n25403 & n25404;
  assign n25406 = n53218 & n25405;
  assign n25407 = n53218 | n25405;
  assign n25408 = ~n25406 & n25407;
  assign n25409 = x125 & x207;
  assign n25410 = n25408 & n25409;
  assign n25411 = n25408 | n25409;
  assign n25412 = ~n25410 & n25411;
  assign n25413 = n53216 & n25412;
  assign n25414 = n53216 | n25412;
  assign n25415 = ~n25413 & n25414;
  assign n25416 = x124 & x208;
  assign n25417 = n25415 & n25416;
  assign n25418 = n25415 | n25416;
  assign n25419 = ~n25417 & n25418;
  assign n25420 = n53214 & n25419;
  assign n25421 = n53214 | n25419;
  assign n25422 = ~n25420 & n25421;
  assign n25423 = x123 & x209;
  assign n25424 = n25422 & n25423;
  assign n25425 = n25422 | n25423;
  assign n25426 = ~n25424 & n25425;
  assign n25427 = n53212 & n25426;
  assign n25428 = n53212 | n25426;
  assign n25429 = ~n25427 & n25428;
  assign n25430 = x122 & x210;
  assign n25431 = n25429 & n25430;
  assign n25432 = n25429 | n25430;
  assign n25433 = ~n25431 & n25432;
  assign n25434 = n53210 & n25433;
  assign n25435 = n53210 | n25433;
  assign n25436 = ~n25434 & n25435;
  assign n25437 = x121 & x211;
  assign n25438 = n25436 & n25437;
  assign n25439 = n25436 | n25437;
  assign n25440 = ~n25438 & n25439;
  assign n25441 = n53208 & n25440;
  assign n25442 = n53208 | n25440;
  assign n25443 = ~n25441 & n25442;
  assign n25444 = x120 & x212;
  assign n25445 = n25443 & n25444;
  assign n25446 = n25443 | n25444;
  assign n25447 = ~n25445 & n25446;
  assign n25448 = n53206 & n25447;
  assign n25449 = n53206 | n25447;
  assign n25450 = ~n25448 & n25449;
  assign n25451 = x119 & x213;
  assign n25452 = n25450 & n25451;
  assign n25453 = n25450 | n25451;
  assign n25454 = ~n25452 & n25453;
  assign n25455 = n53204 & n25454;
  assign n25456 = n53204 | n25454;
  assign n25457 = ~n25455 & n25456;
  assign n25458 = x118 & x214;
  assign n25459 = n25457 & n25458;
  assign n25460 = n25457 | n25458;
  assign n25461 = ~n25459 & n25460;
  assign n25462 = n53202 & n25461;
  assign n25463 = n53202 | n25461;
  assign n25464 = ~n25462 & n25463;
  assign n25465 = x117 & x215;
  assign n25466 = n25464 & n25465;
  assign n25467 = n25464 | n25465;
  assign n25468 = ~n25466 & n25467;
  assign n25469 = n53200 & n25468;
  assign n25470 = n53200 | n25468;
  assign n25471 = ~n25469 & n25470;
  assign n25472 = x116 & x216;
  assign n25473 = n25471 & n25472;
  assign n25474 = n25471 | n25472;
  assign n25475 = ~n25473 & n25474;
  assign n25476 = n53198 & n25475;
  assign n25477 = n53198 | n25475;
  assign n25478 = ~n25476 & n25477;
  assign n25479 = x115 & x217;
  assign n25480 = n25478 & n25479;
  assign n25481 = n25478 | n25479;
  assign n25482 = ~n25480 & n25481;
  assign n25483 = n53196 & n25482;
  assign n25484 = n53196 | n25482;
  assign n25485 = ~n25483 & n25484;
  assign n25486 = x114 & x218;
  assign n25487 = n25485 & n25486;
  assign n25488 = n25485 | n25486;
  assign n25489 = ~n25487 & n25488;
  assign n25490 = n53194 & n25489;
  assign n25491 = n53194 | n25489;
  assign n25492 = ~n25490 & n25491;
  assign n25493 = x113 & x219;
  assign n25494 = n25492 & n25493;
  assign n25495 = n25492 | n25493;
  assign n25496 = ~n25494 & n25495;
  assign n25497 = n25153 & n25496;
  assign n25498 = n25153 | n25496;
  assign n25499 = ~n25497 & n25498;
  assign n25500 = x112 & x220;
  assign n25501 = n25499 & n25500;
  assign n25502 = n25499 | n25500;
  assign n25503 = ~n25501 & n25502;
  assign n68545 = n25153 | n25493;
  assign n68546 = (n25153 & n25492) | (n25153 & n68545) | (n25492 & n68545);
  assign n53361 = (n25494 & n25496) | (n25494 & n68546) | (n25496 & n68546);
  assign n68547 = n25487 | n53194;
  assign n68548 = (n25487 & n25489) | (n25487 & n68547) | (n25489 & n68547);
  assign n25506 = n25480 | n25483;
  assign n25507 = n25473 | n25476;
  assign n25508 = n25466 | n25469;
  assign n25509 = n25459 | n25462;
  assign n25510 = n25452 | n25455;
  assign n25511 = n25445 | n25448;
  assign n25512 = n25438 | n25441;
  assign n53362 = n25431 | n25433;
  assign n53363 = (n25431 & n53210) | (n25431 & n53362) | (n53210 & n53362);
  assign n53364 = n25424 | n25426;
  assign n53365 = (n25424 & n53212) | (n25424 & n53364) | (n53212 & n53364);
  assign n53366 = n25417 | n25419;
  assign n53367 = (n25417 & n53214) | (n25417 & n53366) | (n53214 & n53366);
  assign n53368 = n25410 | n25412;
  assign n53369 = (n25410 & n53216) | (n25410 & n53368) | (n53216 & n53368);
  assign n53220 = (n25055 & n53049) | (n25055 & n53219) | (n53049 & n53219);
  assign n53222 = (n25048 & n53051) | (n25048 & n53221) | (n53051 & n53221);
  assign n53227 = (n68344 & n68462) | (n68344 & n53226) | (n68462 & n53226);
  assign n53379 = n25305 | n25307;
  assign n68549 = n24964 | n25305;
  assign n68550 = (n25305 & n25307) | (n25305 & n68549) | (n25307 & n68549);
  assign n68551 = (n53146 & n53379) | (n53146 & n68550) | (n53379 & n68550);
  assign n68552 = (n53145 & n53379) | (n53145 & n68550) | (n53379 & n68550);
  assign n68553 = (n52896 & n68551) | (n52896 & n68552) | (n68551 & n68552);
  assign n53384 = n25284 | n25286;
  assign n68554 = n24943 | n25284;
  assign n68555 = (n25284 & n25286) | (n25284 & n68554) | (n25286 & n68554);
  assign n68556 = (n53136 & n53384) | (n53136 & n68555) | (n53384 & n68555);
  assign n68557 = (n53135 & n53384) | (n53135 & n68555) | (n53384 & n68555);
  assign n68558 = (n68275 & n68556) | (n68275 & n68557) | (n68556 & n68557);
  assign n53073 = (n52762 & n68377) | (n52762 & n53072) | (n68377 & n53072);
  assign n68563 = n25235 | n25237;
  assign n68564 = (n25235 & n53245) | (n25235 & n68563) | (n53245 & n68563);
  assign n68565 = n24894 | n25235;
  assign n68566 = (n25235 & n25237) | (n25235 & n68565) | (n25237 & n68565);
  assign n68567 = (n68379 & n68564) | (n68379 & n68566) | (n68564 & n68566);
  assign n68568 = (n68381 & n68564) | (n68381 & n68566) | (n68564 & n68566);
  assign n68569 = (n68178 & n68567) | (n68178 & n68568) | (n68567 & n68568);
  assign n25547 = x157 & x176;
  assign n25548 = x156 & x177;
  assign n25549 = n25547 & n25548;
  assign n25550 = n25547 | n25548;
  assign n25551 = ~n25549 & n25550;
  assign n68570 = n25200 | n25202;
  assign n68572 = n25551 & n68570;
  assign n68573 = n25200 & n25551;
  assign n68574 = (n68487 & n68572) | (n68487 & n68573) | (n68572 & n68573);
  assign n68576 = (n68488 & n68572) | (n68488 & n68573) | (n68572 & n68573);
  assign n53415 = (n68195 & n68574) | (n68195 & n68576) | (n68574 & n68576);
  assign n68577 = n25551 | n68570;
  assign n68578 = n25200 | n25551;
  assign n68579 = (n68487 & n68577) | (n68487 & n68578) | (n68577 & n68578);
  assign n68580 = (n68488 & n68577) | (n68488 & n68578) | (n68577 & n68578);
  assign n53418 = (n68195 & n68579) | (n68195 & n68580) | (n68579 & n68580);
  assign n25554 = ~n53415 & n53418;
  assign n25555 = x155 & x178;
  assign n25556 = n25554 & n25555;
  assign n25557 = n25554 | n25555;
  assign n25558 = ~n25556 & n25557;
  assign n68581 = n24866 | n25207;
  assign n68582 = (n25207 & n25209) | (n25207 & n68581) | (n25209 & n68581);
  assign n53419 = n25558 & n68582;
  assign n53408 = n25207 | n25209;
  assign n53420 = n25558 & n53408;
  assign n53421 = (n68389 & n53419) | (n68389 & n53420) | (n53419 & n53420);
  assign n53422 = n25558 | n68582;
  assign n53423 = n25558 | n53408;
  assign n53424 = (n68389 & n53422) | (n68389 & n53423) | (n53422 & n53423);
  assign n25561 = ~n53421 & n53424;
  assign n25562 = x154 & x179;
  assign n25563 = n25561 & n25562;
  assign n25564 = n25561 | n25562;
  assign n25565 = ~n25563 & n25564;
  assign n53405 = n25214 | n25216;
  assign n53425 = n25565 & n53405;
  assign n53426 = n25214 & n25565;
  assign n68583 = (n53425 & n53426) | (n53425 & n68484) | (n53426 & n68484);
  assign n68584 = (n53425 & n53426) | (n53425 & n68483) | (n53426 & n68483);
  assign n68585 = (n67914 & n68583) | (n67914 & n68584) | (n68583 & n68584);
  assign n53428 = n25565 | n53405;
  assign n53429 = n25214 | n25565;
  assign n68586 = (n53428 & n53429) | (n53428 & n68484) | (n53429 & n68484);
  assign n68587 = (n53428 & n53429) | (n53428 & n68483) | (n53429 & n68483);
  assign n68588 = (n67914 & n68586) | (n67914 & n68587) | (n68586 & n68587);
  assign n25568 = ~n68585 & n68588;
  assign n25569 = x153 & x180;
  assign n25570 = n25568 & n25569;
  assign n25571 = n25568 | n25569;
  assign n25572 = ~n25570 & n25571;
  assign n68589 = n24880 | n25221;
  assign n68590 = (n25221 & n25223) | (n25221 & n68589) | (n25223 & n68589);
  assign n53431 = n25572 & n68590;
  assign n53403 = n25221 | n25223;
  assign n53432 = n25572 & n53403;
  assign n53433 = (n68409 & n53431) | (n68409 & n53432) | (n53431 & n53432);
  assign n53434 = n25572 | n68590;
  assign n53435 = n25572 | n53403;
  assign n53436 = (n68409 & n53434) | (n68409 & n53435) | (n53434 & n53435);
  assign n25575 = ~n53433 & n53436;
  assign n25576 = x152 & x181;
  assign n25577 = n25575 & n25576;
  assign n25578 = n25575 | n25576;
  assign n25579 = ~n25577 & n25578;
  assign n53400 = n25228 | n53271;
  assign n68591 = n25579 & n53400;
  assign n53399 = n25228 | n53270;
  assign n68592 = n25579 & n53399;
  assign n68593 = (n68308 & n68591) | (n68308 & n68592) | (n68591 & n68592);
  assign n68594 = n25579 | n53400;
  assign n68595 = n25579 | n53399;
  assign n68596 = (n68308 & n68594) | (n68308 & n68595) | (n68594 & n68595);
  assign n25582 = ~n68593 & n68596;
  assign n25583 = x151 & x182;
  assign n25584 = n25582 & n25583;
  assign n25585 = n25582 | n25583;
  assign n25586 = ~n25584 & n25585;
  assign n25587 = n68569 & n25586;
  assign n25588 = n68569 | n25586;
  assign n25589 = ~n25587 & n25588;
  assign n25590 = x150 & x183;
  assign n25591 = n25589 & n25590;
  assign n25592 = n25589 | n25590;
  assign n25593 = ~n25591 & n25592;
  assign n53394 = n25242 | n25244;
  assign n53437 = n25593 & n53394;
  assign n53438 = n25242 & n25593;
  assign n53439 = (n68479 & n53437) | (n68479 & n53438) | (n53437 & n53438);
  assign n53440 = n25593 | n53394;
  assign n53441 = n25242 | n25593;
  assign n53442 = (n68479 & n53440) | (n68479 & n53441) | (n53440 & n53441);
  assign n25596 = ~n53439 & n53442;
  assign n25597 = x149 & x184;
  assign n25598 = n25596 & n25597;
  assign n25599 = n25596 | n25597;
  assign n25600 = ~n25598 & n25599;
  assign n53392 = n25249 | n53282;
  assign n68597 = n25600 & n53392;
  assign n68561 = n24908 | n25249;
  assign n68562 = (n25249 & n25251) | (n25249 & n68561) | (n25251 & n68561);
  assign n68598 = n25600 & n68562;
  assign n68599 = (n53073 & n68597) | (n53073 & n68598) | (n68597 & n68598);
  assign n68600 = n25600 | n53392;
  assign n68601 = n25600 | n68562;
  assign n68602 = (n53073 & n68600) | (n53073 & n68601) | (n68600 & n68601);
  assign n25603 = ~n68599 & n68602;
  assign n25604 = x148 & x185;
  assign n25605 = n25603 & n25604;
  assign n25606 = n25603 | n25604;
  assign n25607 = ~n25605 & n25606;
  assign n53443 = n25256 & n25607;
  assign n68603 = (n25607 & n53288) | (n25607 & n53443) | (n53288 & n53443);
  assign n68604 = (n25607 & n53289) | (n25607 & n53443) | (n53289 & n53443);
  assign n68605 = (n53070 & n68603) | (n53070 & n68604) | (n68603 & n68604);
  assign n53445 = n25256 | n25607;
  assign n68606 = n53288 | n53445;
  assign n68607 = n53289 | n53445;
  assign n68608 = (n53070 & n68606) | (n53070 & n68607) | (n68606 & n68607);
  assign n25610 = ~n68605 & n68608;
  assign n25611 = x147 & x186;
  assign n25612 = n25610 & n25611;
  assign n25613 = n25610 | n25611;
  assign n25614 = ~n25612 & n25613;
  assign n53389 = n25263 | n25265;
  assign n68609 = n25614 & n53389;
  assign n68559 = n24922 | n25263;
  assign n68560 = (n25263 & n25265) | (n25263 & n68559) | (n25265 & n68559);
  assign n68610 = n25614 & n68560;
  assign n68611 = (n53127 & n68609) | (n53127 & n68610) | (n68609 & n68610);
  assign n68612 = n25614 | n53389;
  assign n68613 = n25614 | n68560;
  assign n68614 = (n53127 & n68612) | (n53127 & n68613) | (n68612 & n68613);
  assign n25617 = ~n68611 & n68614;
  assign n25618 = x146 & x187;
  assign n25619 = n25617 & n25618;
  assign n25620 = n25617 | n25618;
  assign n25621 = ~n25619 & n25620;
  assign n53386 = n25270 | n25272;
  assign n53447 = n25621 & n53386;
  assign n53448 = n25270 & n25621;
  assign n53449 = (n68472 & n53447) | (n68472 & n53448) | (n53447 & n53448);
  assign n53450 = n25621 | n53386;
  assign n53451 = n25270 | n25621;
  assign n53452 = (n68472 & n53450) | (n68472 & n53451) | (n53450 & n53451);
  assign n25624 = ~n53449 & n53452;
  assign n25625 = x145 & x188;
  assign n25626 = n25624 & n25625;
  assign n25627 = n25624 | n25625;
  assign n25628 = ~n25626 & n25627;
  assign n53453 = n25277 & n25628;
  assign n68615 = (n25628 & n53299) | (n25628 & n53453) | (n53299 & n53453);
  assign n68616 = (n25628 & n53298) | (n25628 & n53453) | (n53298 & n53453);
  assign n68617 = (n68373 & n68615) | (n68373 & n68616) | (n68615 & n68616);
  assign n53455 = n25277 | n25628;
  assign n68618 = n53299 | n53455;
  assign n68619 = n53298 | n53455;
  assign n68620 = (n68373 & n68618) | (n68373 & n68619) | (n68618 & n68619);
  assign n25631 = ~n68617 & n68620;
  assign n25632 = x144 & x189;
  assign n25633 = n25631 & n25632;
  assign n25634 = n25631 | n25632;
  assign n25635 = ~n25633 & n25634;
  assign n25636 = n68558 & n25635;
  assign n25637 = n68558 | n25635;
  assign n25638 = ~n25636 & n25637;
  assign n25639 = x143 & x190;
  assign n25640 = n25638 & n25639;
  assign n25641 = n25638 | n25639;
  assign n25642 = ~n25640 & n25641;
  assign n53381 = n25291 | n25293;
  assign n53457 = n25642 & n53381;
  assign n53458 = n25291 & n25642;
  assign n53459 = (n68467 & n53457) | (n68467 & n53458) | (n53457 & n53458);
  assign n53460 = n25642 | n53381;
  assign n53461 = n25291 | n25642;
  assign n53462 = (n68467 & n53460) | (n68467 & n53461) | (n53460 & n53461);
  assign n25645 = ~n53459 & n53462;
  assign n25646 = x142 & x191;
  assign n25647 = n25645 & n25646;
  assign n25648 = n25645 | n25646;
  assign n25649 = ~n25647 & n25648;
  assign n53463 = n25298 & n25649;
  assign n68621 = (n25649 & n53309) | (n25649 & n53463) | (n53309 & n53463);
  assign n68622 = (n25649 & n53308) | (n25649 & n53463) | (n53308 & n53463);
  assign n68623 = (n68368 & n68621) | (n68368 & n68622) | (n68621 & n68622);
  assign n53465 = n25298 | n25649;
  assign n68624 = n53309 | n53465;
  assign n68625 = n53308 | n53465;
  assign n68626 = (n68368 & n68624) | (n68368 & n68625) | (n68624 & n68625);
  assign n25652 = ~n68623 & n68626;
  assign n25653 = x141 & x192;
  assign n25654 = n25652 & n25653;
  assign n25655 = n25652 | n25653;
  assign n25656 = ~n25654 & n25655;
  assign n25657 = n68553 & n25656;
  assign n25658 = n68553 | n25656;
  assign n25659 = ~n25657 & n25658;
  assign n25660 = x140 & x193;
  assign n25661 = n25659 & n25660;
  assign n25662 = n25659 | n25660;
  assign n25663 = ~n25661 & n25662;
  assign n53376 = n25312 | n25314;
  assign n53467 = n25663 & n53376;
  assign n53468 = n25312 & n25663;
  assign n53469 = (n53227 & n53467) | (n53227 & n53468) | (n53467 & n53468);
  assign n53470 = n25663 | n53376;
  assign n53471 = n25312 | n25663;
  assign n53472 = (n53227 & n53470) | (n53227 & n53471) | (n53470 & n53471);
  assign n25666 = ~n53469 & n53472;
  assign n25667 = x139 & x194;
  assign n25668 = n25666 & n25667;
  assign n25669 = n25666 | n25667;
  assign n25670 = ~n25668 & n25669;
  assign n53473 = n25319 & n25670;
  assign n53474 = (n25670 & n68529) | (n25670 & n53473) | (n68529 & n53473);
  assign n53475 = n25319 | n25670;
  assign n53476 = n68529 | n53475;
  assign n25673 = ~n53474 & n53476;
  assign n25674 = x138 & x195;
  assign n25675 = n25673 & n25674;
  assign n25676 = n25673 | n25674;
  assign n25677 = ~n25675 & n25676;
  assign n53477 = n25326 & n25677;
  assign n53478 = (n25677 & n53323) | (n25677 & n53477) | (n53323 & n53477);
  assign n53479 = n25326 | n25677;
  assign n53480 = n53323 | n53479;
  assign n25680 = ~n53478 & n53480;
  assign n25681 = x137 & x196;
  assign n25682 = n25680 & n25681;
  assign n25683 = n25680 | n25681;
  assign n25684 = ~n25682 & n25683;
  assign n53481 = n25333 & n25684;
  assign n53482 = (n25684 & n53327) | (n25684 & n53481) | (n53327 & n53481);
  assign n53483 = n25333 | n25684;
  assign n53484 = n53327 | n53483;
  assign n25687 = ~n53482 & n53484;
  assign n25688 = x136 & x197;
  assign n25689 = n25687 & n25688;
  assign n25690 = n25687 | n25688;
  assign n25691 = ~n25689 & n25690;
  assign n53485 = n25340 & n25691;
  assign n53486 = (n25691 & n53331) | (n25691 & n53485) | (n53331 & n53485);
  assign n53487 = n25340 | n25691;
  assign n53488 = n53331 | n53487;
  assign n25694 = ~n53486 & n53488;
  assign n25695 = x135 & x198;
  assign n25696 = n25694 & n25695;
  assign n25697 = n25694 | n25695;
  assign n25698 = ~n25696 & n25697;
  assign n53489 = n25347 & n25698;
  assign n53490 = (n25698 & n53335) | (n25698 & n53489) | (n53335 & n53489);
  assign n53491 = n25347 | n25698;
  assign n53492 = n53335 | n53491;
  assign n25701 = ~n53490 & n53492;
  assign n25702 = x134 & x199;
  assign n25703 = n25701 & n25702;
  assign n25704 = n25701 | n25702;
  assign n25705 = ~n25703 & n25704;
  assign n53493 = n25354 & n25705;
  assign n53494 = (n25705 & n53339) | (n25705 & n53493) | (n53339 & n53493);
  assign n53495 = n25354 | n25705;
  assign n53496 = n53339 | n53495;
  assign n25708 = ~n53494 & n53496;
  assign n25709 = x133 & x200;
  assign n25710 = n25708 & n25709;
  assign n25711 = n25708 | n25709;
  assign n25712 = ~n25710 & n25711;
  assign n53497 = n25361 & n25712;
  assign n53498 = (n25712 & n53343) | (n25712 & n53497) | (n53343 & n53497);
  assign n53499 = n25361 | n25712;
  assign n53500 = n53343 | n53499;
  assign n25715 = ~n53498 & n53500;
  assign n25716 = x132 & x201;
  assign n25717 = n25715 & n25716;
  assign n25718 = n25715 | n25716;
  assign n25719 = ~n25717 & n25718;
  assign n53501 = n25368 & n25719;
  assign n53502 = (n25719 & n53347) | (n25719 & n53501) | (n53347 & n53501);
  assign n53503 = n25368 | n25719;
  assign n53504 = n53347 | n53503;
  assign n25722 = ~n53502 & n53504;
  assign n25723 = x131 & x202;
  assign n25724 = n25722 & n25723;
  assign n25725 = n25722 | n25723;
  assign n25726 = ~n25724 & n25725;
  assign n53505 = n25375 & n25726;
  assign n53506 = (n25726 & n53351) | (n25726 & n53505) | (n53351 & n53505);
  assign n53507 = n25375 | n25726;
  assign n53508 = n53351 | n53507;
  assign n25729 = ~n53506 & n53508;
  assign n25730 = x130 & x203;
  assign n25731 = n25729 & n25730;
  assign n25732 = n25729 | n25730;
  assign n25733 = ~n25731 & n25732;
  assign n53509 = n25382 & n25733;
  assign n53510 = (n25733 & n53356) | (n25733 & n53509) | (n53356 & n53509);
  assign n53511 = n25382 | n25733;
  assign n53512 = n53356 | n53511;
  assign n25736 = ~n53510 & n53512;
  assign n25737 = x129 & x204;
  assign n25738 = n25736 & n25737;
  assign n25739 = n25736 | n25737;
  assign n25740 = ~n25738 & n25739;
  assign n53374 = n25389 | n25391;
  assign n53513 = n25740 & n53374;
  assign n53514 = n25389 & n25740;
  assign n53515 = (n53222 & n53513) | (n53222 & n53514) | (n53513 & n53514);
  assign n53516 = n25740 | n53374;
  assign n53517 = n25389 | n25740;
  assign n53518 = (n53222 & n53516) | (n53222 & n53517) | (n53516 & n53517);
  assign n25743 = ~n53515 & n53518;
  assign n25744 = x128 & x205;
  assign n25745 = n25743 & n25744;
  assign n25746 = n25743 | n25744;
  assign n25747 = ~n25745 & n25746;
  assign n53372 = n25396 | n25398;
  assign n68627 = n25747 & n53372;
  assign n68628 = n25396 & n25747;
  assign n68629 = (n53220 & n68627) | (n53220 & n68628) | (n68627 & n68628);
  assign n68630 = n25747 | n53372;
  assign n68631 = n25396 | n25747;
  assign n68632 = (n53220 & n68630) | (n53220 & n68631) | (n68630 & n68631);
  assign n25750 = ~n68629 & n68632;
  assign n25751 = x127 & x206;
  assign n25752 = n25750 & n25751;
  assign n25753 = n25750 | n25751;
  assign n25754 = ~n25752 & n25753;
  assign n53370 = n25403 | n25405;
  assign n68633 = n25754 & n53370;
  assign n68634 = n25403 & n25754;
  assign n68635 = (n53218 & n68633) | (n53218 & n68634) | (n68633 & n68634);
  assign n68636 = n25754 | n53370;
  assign n68637 = n25403 | n25754;
  assign n68638 = (n53218 & n68636) | (n53218 & n68637) | (n68636 & n68637);
  assign n25757 = ~n68635 & n68638;
  assign n25758 = x126 & x207;
  assign n25759 = n25757 & n25758;
  assign n25760 = n25757 | n25758;
  assign n25761 = ~n25759 & n25760;
  assign n25762 = n53369 & n25761;
  assign n25763 = n53369 | n25761;
  assign n25764 = ~n25762 & n25763;
  assign n25765 = x125 & x208;
  assign n25766 = n25764 & n25765;
  assign n25767 = n25764 | n25765;
  assign n25768 = ~n25766 & n25767;
  assign n25769 = n53367 & n25768;
  assign n25770 = n53367 | n25768;
  assign n25771 = ~n25769 & n25770;
  assign n25772 = x124 & x209;
  assign n25773 = n25771 & n25772;
  assign n25774 = n25771 | n25772;
  assign n25775 = ~n25773 & n25774;
  assign n25776 = n53365 & n25775;
  assign n25777 = n53365 | n25775;
  assign n25778 = ~n25776 & n25777;
  assign n25779 = x123 & x210;
  assign n25780 = n25778 & n25779;
  assign n25781 = n25778 | n25779;
  assign n25782 = ~n25780 & n25781;
  assign n25783 = n53363 & n25782;
  assign n25784 = n53363 | n25782;
  assign n25785 = ~n25783 & n25784;
  assign n25786 = x122 & x211;
  assign n25787 = n25785 & n25786;
  assign n25788 = n25785 | n25786;
  assign n25789 = ~n25787 & n25788;
  assign n25790 = n25512 & n25789;
  assign n25791 = n25512 | n25789;
  assign n25792 = ~n25790 & n25791;
  assign n25793 = x121 & x212;
  assign n25794 = n25792 & n25793;
  assign n25795 = n25792 | n25793;
  assign n25796 = ~n25794 & n25795;
  assign n25797 = n25511 & n25796;
  assign n25798 = n25511 | n25796;
  assign n25799 = ~n25797 & n25798;
  assign n25800 = x120 & x213;
  assign n25801 = n25799 & n25800;
  assign n25802 = n25799 | n25800;
  assign n25803 = ~n25801 & n25802;
  assign n25804 = n25510 & n25803;
  assign n25805 = n25510 | n25803;
  assign n25806 = ~n25804 & n25805;
  assign n25807 = x119 & x214;
  assign n25808 = n25806 & n25807;
  assign n25809 = n25806 | n25807;
  assign n25810 = ~n25808 & n25809;
  assign n25811 = n25509 & n25810;
  assign n25812 = n25509 | n25810;
  assign n25813 = ~n25811 & n25812;
  assign n25814 = x118 & x215;
  assign n25815 = n25813 & n25814;
  assign n25816 = n25813 | n25814;
  assign n25817 = ~n25815 & n25816;
  assign n25818 = n25508 & n25817;
  assign n25819 = n25508 | n25817;
  assign n25820 = ~n25818 & n25819;
  assign n25821 = x117 & x216;
  assign n25822 = n25820 & n25821;
  assign n25823 = n25820 | n25821;
  assign n25824 = ~n25822 & n25823;
  assign n25825 = n25507 & n25824;
  assign n25826 = n25507 | n25824;
  assign n25827 = ~n25825 & n25826;
  assign n25828 = x116 & x217;
  assign n25829 = n25827 & n25828;
  assign n25830 = n25827 | n25828;
  assign n25831 = ~n25829 & n25830;
  assign n25832 = n25506 & n25831;
  assign n25833 = n25506 | n25831;
  assign n25834 = ~n25832 & n25833;
  assign n25835 = x115 & x218;
  assign n25836 = n25834 & n25835;
  assign n25837 = n25834 | n25835;
  assign n25838 = ~n25836 & n25837;
  assign n25839 = n68548 & n25838;
  assign n25840 = n68548 | n25838;
  assign n25841 = ~n25839 & n25840;
  assign n25842 = x114 & x219;
  assign n25843 = n25841 & n25842;
  assign n25844 = n25841 | n25842;
  assign n25845 = ~n25843 & n25844;
  assign n25846 = n53361 & n25845;
  assign n25847 = n53361 | n25845;
  assign n25848 = ~n25846 & n25847;
  assign n25849 = x113 & x220;
  assign n25850 = n25848 & n25849;
  assign n25851 = n25848 | n25849;
  assign n25852 = ~n25850 & n25851;
  assign n25853 = n25501 & n25852;
  assign n25854 = n25501 | n25852;
  assign n25855 = ~n25853 & n25854;
  assign n25856 = x112 & x221;
  assign n25857 = n25855 & n25856;
  assign n25858 = n25855 | n25856;
  assign n25859 = ~n25857 & n25858;
  assign n68639 = n25501 | n25849;
  assign n68640 = (n25501 & n25848) | (n25501 & n68639) | (n25848 & n68639);
  assign n53520 = (n25850 & n25852) | (n25850 & n68640) | (n25852 & n68640);
  assign n53521 = n25843 | n53361;
  assign n53522 = (n25843 & n25845) | (n25843 & n53521) | (n25845 & n53521);
  assign n68641 = n25836 | n68548;
  assign n68642 = (n25836 & n25838) | (n25836 & n68641) | (n25838 & n68641);
  assign n25863 = n25829 | n25832;
  assign n25864 = n25822 | n25825;
  assign n25865 = n25815 | n25818;
  assign n25866 = n25808 | n25811;
  assign n25867 = n25801 | n25804;
  assign n25868 = n25794 | n25797;
  assign n53523 = n25787 | n25789;
  assign n53524 = (n25512 & n25787) | (n25512 & n53523) | (n25787 & n53523);
  assign n53525 = n25780 | n25782;
  assign n53526 = (n25780 & n53363) | (n25780 & n53525) | (n53363 & n53525);
  assign n53527 = n25773 | n25775;
  assign n53528 = (n25773 & n53365) | (n25773 & n53527) | (n53365 & n53527);
  assign n53529 = n25766 | n25768;
  assign n53530 = (n25766 & n53367) | (n25766 & n53529) | (n53367 & n53529);
  assign n53371 = (n25403 & n53218) | (n25403 & n53370) | (n53218 & n53370);
  assign n53373 = (n25396 & n53220) | (n25396 & n53372) | (n53220 & n53372);
  assign n53543 = n25647 | n25649;
  assign n68645 = n25298 | n25647;
  assign n68646 = (n25647 & n25649) | (n25647 & n68645) | (n25649 & n68645);
  assign n68647 = (n53309 & n53543) | (n53309 & n68646) | (n53543 & n68646);
  assign n68648 = (n53308 & n53543) | (n53308 & n68646) | (n53543 & n68646);
  assign n68649 = (n68368 & n68647) | (n68368 & n68648) | (n68647 & n68648);
  assign n53548 = n25626 | n25628;
  assign n68650 = n25277 | n25626;
  assign n68651 = (n25626 & n25628) | (n25626 & n68650) | (n25628 & n68650);
  assign n68652 = (n53299 & n53548) | (n53299 & n68651) | (n53548 & n68651);
  assign n68653 = (n53298 & n53548) | (n53298 & n68651) | (n53548 & n68651);
  assign n68654 = (n68373 & n68652) | (n68373 & n68653) | (n68652 & n68653);
  assign n53390 = (n53127 & n68560) | (n53127 & n53389) | (n68560 & n53389);
  assign n53553 = n25605 | n25607;
  assign n68655 = n25256 | n25605;
  assign n68656 = (n25605 & n25607) | (n25605 & n68655) | (n25607 & n68655);
  assign n68657 = (n53288 & n53553) | (n53288 & n68656) | (n53553 & n68656);
  assign n68658 = (n53289 & n53553) | (n53289 & n68656) | (n53553 & n68656);
  assign n68659 = (n53070 & n68657) | (n53070 & n68658) | (n68657 & n68658);
  assign n25904 = x158 & x176;
  assign n25905 = x157 & x177;
  assign n25906 = n25904 & n25905;
  assign n25907 = n25904 | n25905;
  assign n25908 = ~n25906 & n25907;
  assign n68665 = n25549 & n25908;
  assign n68666 = (n25908 & n68574) | (n25908 & n68665) | (n68574 & n68665);
  assign n68667 = (n25908 & n68576) | (n25908 & n68665) | (n68576 & n68665);
  assign n53578 = (n68195 & n68666) | (n68195 & n68667) | (n68666 & n68667);
  assign n68668 = n25549 | n25908;
  assign n68669 = n68574 | n68668;
  assign n68670 = n68576 | n68668;
  assign n53581 = (n68195 & n68669) | (n68195 & n68670) | (n68669 & n68670);
  assign n25911 = ~n53578 & n53581;
  assign n25912 = x156 & x178;
  assign n25913 = n25911 & n25912;
  assign n25914 = n25911 | n25912;
  assign n25915 = ~n25913 & n25914;
  assign n68671 = n25556 | n25558;
  assign n68672 = (n25556 & n68582) | (n25556 & n68671) | (n68582 & n68671);
  assign n53582 = n25915 & n68672;
  assign n68673 = (n25556 & n53408) | (n25556 & n68671) | (n53408 & n68671);
  assign n53583 = n25915 & n68673;
  assign n53584 = (n68389 & n53582) | (n68389 & n53583) | (n53582 & n53583);
  assign n53585 = n25915 | n68672;
  assign n53586 = n25915 | n68673;
  assign n53587 = (n68389 & n53585) | (n68389 & n53586) | (n53585 & n53586);
  assign n25918 = ~n53584 & n53587;
  assign n25919 = x155 & x179;
  assign n25920 = n25918 & n25919;
  assign n25921 = n25918 | n25919;
  assign n25922 = ~n25920 & n25921;
  assign n68674 = n25563 | n25565;
  assign n68675 = (n25563 & n53405) | (n25563 & n68674) | (n53405 & n68674);
  assign n53588 = n25922 & n68675;
  assign n68676 = n25214 | n25563;
  assign n68677 = (n25563 & n25565) | (n25563 & n68676) | (n25565 & n68676);
  assign n53589 = n25922 & n68677;
  assign n68678 = (n53588 & n53589) | (n53588 & n68484) | (n53589 & n68484);
  assign n68679 = (n53588 & n53589) | (n53588 & n68483) | (n53589 & n68483);
  assign n68680 = (n67914 & n68678) | (n67914 & n68679) | (n68678 & n68679);
  assign n53591 = n25922 | n68675;
  assign n53592 = n25922 | n68677;
  assign n68681 = (n53591 & n53592) | (n53591 & n68484) | (n53592 & n68484);
  assign n68682 = (n53591 & n53592) | (n53591 & n68483) | (n53592 & n68483);
  assign n68683 = (n67914 & n68681) | (n67914 & n68682) | (n68681 & n68682);
  assign n25925 = ~n68680 & n68683;
  assign n25926 = x154 & x180;
  assign n25927 = n25925 & n25926;
  assign n25928 = n25925 | n25926;
  assign n25929 = ~n25927 & n25928;
  assign n68662 = n25570 | n25572;
  assign n68664 = (n25570 & n53403) | (n25570 & n68662) | (n53403 & n68662);
  assign n68684 = n25929 & n68664;
  assign n68663 = (n25570 & n68590) | (n25570 & n68662) | (n68590 & n68662);
  assign n68685 = n25929 & n68663;
  assign n68686 = (n68409 & n68684) | (n68409 & n68685) | (n68684 & n68685);
  assign n68687 = n25929 | n68664;
  assign n68688 = n25929 | n68663;
  assign n68689 = (n68409 & n68687) | (n68409 & n68688) | (n68687 & n68688);
  assign n25932 = ~n68686 & n68689;
  assign n25933 = x153 & x181;
  assign n25934 = n25932 & n25933;
  assign n25935 = n25932 | n25933;
  assign n25936 = ~n25934 & n25935;
  assign n53562 = n25577 | n25579;
  assign n53594 = n25936 & n53562;
  assign n53595 = n25577 & n25936;
  assign n68690 = (n53400 & n53594) | (n53400 & n53595) | (n53594 & n53595);
  assign n68691 = (n53399 & n53594) | (n53399 & n53595) | (n53594 & n53595);
  assign n68692 = (n68308 & n68690) | (n68308 & n68691) | (n68690 & n68691);
  assign n53597 = n25936 | n53562;
  assign n53598 = n25577 | n25936;
  assign n68693 = (n53400 & n53597) | (n53400 & n53598) | (n53597 & n53598);
  assign n68694 = (n53399 & n53597) | (n53399 & n53598) | (n53597 & n53598);
  assign n68695 = (n68308 & n68693) | (n68308 & n68694) | (n68693 & n68694);
  assign n25939 = ~n68692 & n68695;
  assign n25940 = x152 & x182;
  assign n25941 = n25939 & n25940;
  assign n25942 = n25939 | n25940;
  assign n25943 = ~n25941 & n25942;
  assign n53560 = n25584 | n25586;
  assign n53600 = n25943 & n53560;
  assign n53601 = n25584 & n25943;
  assign n53602 = (n68569 & n53600) | (n68569 & n53601) | (n53600 & n53601);
  assign n53603 = n25943 | n53560;
  assign n53604 = n25584 | n25943;
  assign n53605 = (n68569 & n53603) | (n68569 & n53604) | (n53603 & n53604);
  assign n25946 = ~n53602 & n53605;
  assign n25947 = x151 & x183;
  assign n25948 = n25946 & n25947;
  assign n25949 = n25946 | n25947;
  assign n25950 = ~n25948 & n25949;
  assign n53558 = n25591 | n53437;
  assign n68696 = n25950 & n53558;
  assign n68660 = n25242 | n25591;
  assign n68661 = (n25591 & n25593) | (n25591 & n68660) | (n25593 & n68660);
  assign n68697 = n25950 & n68661;
  assign n68698 = (n68479 & n68696) | (n68479 & n68697) | (n68696 & n68697);
  assign n68699 = n25950 | n53558;
  assign n68700 = n25950 | n68661;
  assign n68701 = (n68479 & n68699) | (n68479 & n68700) | (n68699 & n68700);
  assign n25953 = ~n68698 & n68701;
  assign n25954 = x150 & x184;
  assign n25955 = n25953 & n25954;
  assign n25956 = n25953 | n25954;
  assign n25957 = ~n25955 & n25956;
  assign n53555 = n25598 | n25600;
  assign n53606 = n25957 & n53555;
  assign n53607 = n25598 & n25957;
  assign n68702 = (n53392 & n53606) | (n53392 & n53607) | (n53606 & n53607);
  assign n68703 = (n53606 & n53607) | (n53606 & n68562) | (n53607 & n68562);
  assign n68704 = (n53073 & n68702) | (n53073 & n68703) | (n68702 & n68703);
  assign n53609 = n25957 | n53555;
  assign n53610 = n25598 | n25957;
  assign n68705 = (n53392 & n53609) | (n53392 & n53610) | (n53609 & n53610);
  assign n68706 = (n53609 & n53610) | (n53609 & n68562) | (n53610 & n68562);
  assign n68707 = (n53073 & n68705) | (n53073 & n68706) | (n68705 & n68706);
  assign n25960 = ~n68704 & n68707;
  assign n25961 = x149 & x185;
  assign n25962 = n25960 & n25961;
  assign n25963 = n25960 | n25961;
  assign n25964 = ~n25962 & n25963;
  assign n25965 = n68659 & n25964;
  assign n25966 = n68659 | n25964;
  assign n25967 = ~n25965 & n25966;
  assign n25968 = x148 & x186;
  assign n25969 = n25967 & n25968;
  assign n25970 = n25967 | n25968;
  assign n25971 = ~n25969 & n25970;
  assign n53550 = n25612 | n25614;
  assign n53612 = n25971 & n53550;
  assign n53613 = n25612 & n25971;
  assign n53614 = (n53390 & n53612) | (n53390 & n53613) | (n53612 & n53613);
  assign n53615 = n25971 | n53550;
  assign n53616 = n25612 | n25971;
  assign n53617 = (n53390 & n53615) | (n53390 & n53616) | (n53615 & n53616);
  assign n25974 = ~n53614 & n53617;
  assign n25975 = x147 & x187;
  assign n25976 = n25974 & n25975;
  assign n25977 = n25974 | n25975;
  assign n25978 = ~n25976 & n25977;
  assign n53618 = n25619 & n25978;
  assign n53619 = (n25978 & n53449) | (n25978 & n53618) | (n53449 & n53618);
  assign n53620 = n25619 | n25978;
  assign n53621 = n53449 | n53620;
  assign n25981 = ~n53619 & n53621;
  assign n25982 = x146 & x188;
  assign n25983 = n25981 & n25982;
  assign n25984 = n25981 | n25982;
  assign n25985 = ~n25983 & n25984;
  assign n25986 = n68654 & n25985;
  assign n25987 = n68654 | n25985;
  assign n25988 = ~n25986 & n25987;
  assign n25989 = x145 & x189;
  assign n25990 = n25988 & n25989;
  assign n25991 = n25988 | n25989;
  assign n25992 = ~n25990 & n25991;
  assign n53545 = n25633 | n25635;
  assign n53622 = n25992 & n53545;
  assign n53623 = n25633 & n25992;
  assign n53624 = (n68558 & n53622) | (n68558 & n53623) | (n53622 & n53623);
  assign n53625 = n25992 | n53545;
  assign n53626 = n25633 | n25992;
  assign n53627 = (n68558 & n53625) | (n68558 & n53626) | (n53625 & n53626);
  assign n25995 = ~n53624 & n53627;
  assign n25996 = x144 & x190;
  assign n25997 = n25995 & n25996;
  assign n25998 = n25995 | n25996;
  assign n25999 = ~n25997 & n25998;
  assign n53628 = n25640 & n25999;
  assign n68708 = (n25999 & n53458) | (n25999 & n53628) | (n53458 & n53628);
  assign n68709 = (n25999 & n53457) | (n25999 & n53628) | (n53457 & n53628);
  assign n68710 = (n68467 & n68708) | (n68467 & n68709) | (n68708 & n68709);
  assign n53630 = n25640 | n25999;
  assign n68711 = n53458 | n53630;
  assign n68712 = n53457 | n53630;
  assign n68713 = (n68467 & n68711) | (n68467 & n68712) | (n68711 & n68712);
  assign n26002 = ~n68710 & n68713;
  assign n26003 = x143 & x191;
  assign n26004 = n26002 & n26003;
  assign n26005 = n26002 | n26003;
  assign n26006 = ~n26004 & n26005;
  assign n26007 = n68649 & n26006;
  assign n26008 = n68649 | n26006;
  assign n26009 = ~n26007 & n26008;
  assign n26010 = x142 & x192;
  assign n26011 = n26009 & n26010;
  assign n26012 = n26009 | n26010;
  assign n26013 = ~n26011 & n26012;
  assign n53540 = n25654 | n25656;
  assign n53632 = n26013 & n53540;
  assign n53633 = n25654 & n26013;
  assign n53634 = (n68553 & n53632) | (n68553 & n53633) | (n53632 & n53633);
  assign n53635 = n26013 | n53540;
  assign n53636 = n25654 | n26013;
  assign n53637 = (n68553 & n53635) | (n68553 & n53636) | (n53635 & n53636);
  assign n26016 = ~n53634 & n53637;
  assign n26017 = x141 & x193;
  assign n26018 = n26016 & n26017;
  assign n26019 = n26016 | n26017;
  assign n26020 = ~n26018 & n26019;
  assign n53638 = n25661 & n26020;
  assign n68714 = (n26020 & n53468) | (n26020 & n53638) | (n53468 & n53638);
  assign n68715 = (n26020 & n53467) | (n26020 & n53638) | (n53467 & n53638);
  assign n68716 = (n53227 & n68714) | (n53227 & n68715) | (n68714 & n68715);
  assign n53640 = n25661 | n26020;
  assign n68717 = n53468 | n53640;
  assign n68718 = n53467 | n53640;
  assign n68719 = (n53227 & n68717) | (n53227 & n68718) | (n68717 & n68718);
  assign n26023 = ~n68716 & n68719;
  assign n26024 = x140 & x194;
  assign n26025 = n26023 & n26024;
  assign n26026 = n26023 | n26024;
  assign n26027 = ~n26025 & n26026;
  assign n53538 = n25668 | n25670;
  assign n68720 = n26027 & n53538;
  assign n68643 = n25319 | n25668;
  assign n68644 = (n25668 & n25670) | (n25668 & n68643) | (n25670 & n68643);
  assign n68721 = n26027 & n68644;
  assign n68722 = (n68529 & n68720) | (n68529 & n68721) | (n68720 & n68721);
  assign n68723 = n26027 | n53538;
  assign n68724 = n26027 | n68644;
  assign n68725 = (n68529 & n68723) | (n68529 & n68724) | (n68723 & n68724);
  assign n26030 = ~n68722 & n68725;
  assign n26031 = x139 & x195;
  assign n26032 = n26030 & n26031;
  assign n26033 = n26030 | n26031;
  assign n26034 = ~n26032 & n26033;
  assign n53642 = n25675 & n26034;
  assign n68726 = (n26034 & n53477) | (n26034 & n53642) | (n53477 & n53642);
  assign n68727 = (n25677 & n26034) | (n25677 & n53642) | (n26034 & n53642);
  assign n68728 = (n53323 & n68726) | (n53323 & n68727) | (n68726 & n68727);
  assign n53644 = n25675 | n26034;
  assign n68729 = n53477 | n53644;
  assign n68730 = n25677 | n53644;
  assign n68731 = (n53323 & n68729) | (n53323 & n68730) | (n68729 & n68730);
  assign n26037 = ~n68728 & n68731;
  assign n26038 = x138 & x196;
  assign n26039 = n26037 & n26038;
  assign n26040 = n26037 | n26038;
  assign n26041 = ~n26039 & n26040;
  assign n53646 = n25682 & n26041;
  assign n53647 = (n26041 & n53482) | (n26041 & n53646) | (n53482 & n53646);
  assign n53648 = n25682 | n26041;
  assign n53649 = n53482 | n53648;
  assign n26044 = ~n53647 & n53649;
  assign n26045 = x137 & x197;
  assign n26046 = n26044 & n26045;
  assign n26047 = n26044 | n26045;
  assign n26048 = ~n26046 & n26047;
  assign n53650 = n25689 & n26048;
  assign n53651 = (n26048 & n53486) | (n26048 & n53650) | (n53486 & n53650);
  assign n53652 = n25689 | n26048;
  assign n53653 = n53486 | n53652;
  assign n26051 = ~n53651 & n53653;
  assign n26052 = x136 & x198;
  assign n26053 = n26051 & n26052;
  assign n26054 = n26051 | n26052;
  assign n26055 = ~n26053 & n26054;
  assign n53654 = n25696 & n26055;
  assign n53655 = (n26055 & n53490) | (n26055 & n53654) | (n53490 & n53654);
  assign n53656 = n25696 | n26055;
  assign n53657 = n53490 | n53656;
  assign n26058 = ~n53655 & n53657;
  assign n26059 = x135 & x199;
  assign n26060 = n26058 & n26059;
  assign n26061 = n26058 | n26059;
  assign n26062 = ~n26060 & n26061;
  assign n53658 = n25703 & n26062;
  assign n53659 = (n26062 & n53494) | (n26062 & n53658) | (n53494 & n53658);
  assign n53660 = n25703 | n26062;
  assign n53661 = n53494 | n53660;
  assign n26065 = ~n53659 & n53661;
  assign n26066 = x134 & x200;
  assign n26067 = n26065 & n26066;
  assign n26068 = n26065 | n26066;
  assign n26069 = ~n26067 & n26068;
  assign n53662 = n25710 & n26069;
  assign n53663 = (n26069 & n53498) | (n26069 & n53662) | (n53498 & n53662);
  assign n53664 = n25710 | n26069;
  assign n53665 = n53498 | n53664;
  assign n26072 = ~n53663 & n53665;
  assign n26073 = x133 & x201;
  assign n26074 = n26072 & n26073;
  assign n26075 = n26072 | n26073;
  assign n26076 = ~n26074 & n26075;
  assign n53666 = n25717 & n26076;
  assign n53667 = (n26076 & n53502) | (n26076 & n53666) | (n53502 & n53666);
  assign n53668 = n25717 | n26076;
  assign n53669 = n53502 | n53668;
  assign n26079 = ~n53667 & n53669;
  assign n26080 = x132 & x202;
  assign n26081 = n26079 & n26080;
  assign n26082 = n26079 | n26080;
  assign n26083 = ~n26081 & n26082;
  assign n53670 = n25724 & n26083;
  assign n53671 = (n26083 & n53506) | (n26083 & n53670) | (n53506 & n53670);
  assign n53672 = n25724 | n26083;
  assign n53673 = n53506 | n53672;
  assign n26086 = ~n53671 & n53673;
  assign n26087 = x131 & x203;
  assign n26088 = n26086 & n26087;
  assign n26089 = n26086 | n26087;
  assign n26090 = ~n26088 & n26089;
  assign n53674 = n25731 & n26090;
  assign n53675 = (n26090 & n53510) | (n26090 & n53674) | (n53510 & n53674);
  assign n53676 = n25731 | n26090;
  assign n53677 = n53510 | n53676;
  assign n26093 = ~n53675 & n53677;
  assign n26094 = x130 & x204;
  assign n26095 = n26093 & n26094;
  assign n26096 = n26093 | n26094;
  assign n26097 = ~n26095 & n26096;
  assign n53678 = n25738 & n26097;
  assign n53679 = (n26097 & n53515) | (n26097 & n53678) | (n53515 & n53678);
  assign n53680 = n25738 | n26097;
  assign n53681 = n53515 | n53680;
  assign n26100 = ~n53679 & n53681;
  assign n26101 = x129 & x205;
  assign n26102 = n26100 & n26101;
  assign n26103 = n26100 | n26101;
  assign n26104 = ~n26102 & n26103;
  assign n53535 = n25745 | n25747;
  assign n53682 = n26104 & n53535;
  assign n53683 = n25745 & n26104;
  assign n53684 = (n53373 & n53682) | (n53373 & n53683) | (n53682 & n53683);
  assign n53685 = n26104 | n53535;
  assign n53686 = n25745 | n26104;
  assign n53687 = (n53373 & n53685) | (n53373 & n53686) | (n53685 & n53686);
  assign n26107 = ~n53684 & n53687;
  assign n26108 = x128 & x206;
  assign n26109 = n26107 & n26108;
  assign n26110 = n26107 | n26108;
  assign n26111 = ~n26109 & n26110;
  assign n53533 = n25752 | n25754;
  assign n68732 = n26111 & n53533;
  assign n68733 = n25752 & n26111;
  assign n68734 = (n53371 & n68732) | (n53371 & n68733) | (n68732 & n68733);
  assign n68735 = n26111 | n53533;
  assign n68736 = n25752 | n26111;
  assign n68737 = (n53371 & n68735) | (n53371 & n68736) | (n68735 & n68736);
  assign n26114 = ~n68734 & n68737;
  assign n26115 = x127 & x207;
  assign n26116 = n26114 & n26115;
  assign n26117 = n26114 | n26115;
  assign n26118 = ~n26116 & n26117;
  assign n53531 = n25759 | n25761;
  assign n68738 = n26118 & n53531;
  assign n68739 = n25759 & n26118;
  assign n68740 = (n53369 & n68738) | (n53369 & n68739) | (n68738 & n68739);
  assign n68741 = n26118 | n53531;
  assign n68742 = n25759 | n26118;
  assign n68743 = (n53369 & n68741) | (n53369 & n68742) | (n68741 & n68742);
  assign n26121 = ~n68740 & n68743;
  assign n26122 = x126 & x208;
  assign n26123 = n26121 & n26122;
  assign n26124 = n26121 | n26122;
  assign n26125 = ~n26123 & n26124;
  assign n26126 = n53530 & n26125;
  assign n26127 = n53530 | n26125;
  assign n26128 = ~n26126 & n26127;
  assign n26129 = x125 & x209;
  assign n26130 = n26128 & n26129;
  assign n26131 = n26128 | n26129;
  assign n26132 = ~n26130 & n26131;
  assign n26133 = n53528 & n26132;
  assign n26134 = n53528 | n26132;
  assign n26135 = ~n26133 & n26134;
  assign n26136 = x124 & x210;
  assign n26137 = n26135 & n26136;
  assign n26138 = n26135 | n26136;
  assign n26139 = ~n26137 & n26138;
  assign n26140 = n53526 & n26139;
  assign n26141 = n53526 | n26139;
  assign n26142 = ~n26140 & n26141;
  assign n26143 = x123 & x211;
  assign n26144 = n26142 & n26143;
  assign n26145 = n26142 | n26143;
  assign n26146 = ~n26144 & n26145;
  assign n26147 = n53524 & n26146;
  assign n26148 = n53524 | n26146;
  assign n26149 = ~n26147 & n26148;
  assign n26150 = x122 & x212;
  assign n26151 = n26149 & n26150;
  assign n26152 = n26149 | n26150;
  assign n26153 = ~n26151 & n26152;
  assign n26154 = n25868 & n26153;
  assign n26155 = n25868 | n26153;
  assign n26156 = ~n26154 & n26155;
  assign n26157 = x121 & x213;
  assign n26158 = n26156 & n26157;
  assign n26159 = n26156 | n26157;
  assign n26160 = ~n26158 & n26159;
  assign n26161 = n25867 & n26160;
  assign n26162 = n25867 | n26160;
  assign n26163 = ~n26161 & n26162;
  assign n26164 = x120 & x214;
  assign n26165 = n26163 & n26164;
  assign n26166 = n26163 | n26164;
  assign n26167 = ~n26165 & n26166;
  assign n26168 = n25866 & n26167;
  assign n26169 = n25866 | n26167;
  assign n26170 = ~n26168 & n26169;
  assign n26171 = x119 & x215;
  assign n26172 = n26170 & n26171;
  assign n26173 = n26170 | n26171;
  assign n26174 = ~n26172 & n26173;
  assign n26175 = n25865 & n26174;
  assign n26176 = n25865 | n26174;
  assign n26177 = ~n26175 & n26176;
  assign n26178 = x118 & x216;
  assign n26179 = n26177 & n26178;
  assign n26180 = n26177 | n26178;
  assign n26181 = ~n26179 & n26180;
  assign n26182 = n25864 & n26181;
  assign n26183 = n25864 | n26181;
  assign n26184 = ~n26182 & n26183;
  assign n26185 = x117 & x217;
  assign n26186 = n26184 & n26185;
  assign n26187 = n26184 | n26185;
  assign n26188 = ~n26186 & n26187;
  assign n26189 = n25863 & n26188;
  assign n26190 = n25863 | n26188;
  assign n26191 = ~n26189 & n26190;
  assign n26192 = x116 & x218;
  assign n26193 = n26191 & n26192;
  assign n26194 = n26191 | n26192;
  assign n26195 = ~n26193 & n26194;
  assign n26196 = n68642 & n26195;
  assign n26197 = n68642 | n26195;
  assign n26198 = ~n26196 & n26197;
  assign n26199 = x115 & x219;
  assign n26200 = n26198 & n26199;
  assign n26201 = n26198 | n26199;
  assign n26202 = ~n26200 & n26201;
  assign n26203 = n53522 & n26202;
  assign n26204 = n53522 | n26202;
  assign n26205 = ~n26203 & n26204;
  assign n26206 = x114 & x220;
  assign n26207 = n26205 & n26206;
  assign n26208 = n26205 | n26206;
  assign n26209 = ~n26207 & n26208;
  assign n26210 = n53520 & n26209;
  assign n26211 = n53520 | n26209;
  assign n26212 = ~n26210 & n26211;
  assign n26213 = x113 & x221;
  assign n26214 = n26212 & n26213;
  assign n26215 = n26212 | n26213;
  assign n26216 = ~n26214 & n26215;
  assign n26217 = n25857 & n26216;
  assign n26218 = n25857 | n26216;
  assign n26219 = ~n26217 & n26218;
  assign n26220 = x112 & x222;
  assign n26221 = n26219 & n26220;
  assign n26222 = n26219 | n26220;
  assign n26223 = ~n26221 & n26222;
  assign n68744 = n25857 | n26213;
  assign n68745 = (n25857 & n26212) | (n25857 & n68744) | (n26212 & n68744);
  assign n53689 = (n26214 & n26216) | (n26214 & n68745) | (n26216 & n68745);
  assign n53690 = n26207 | n53520;
  assign n53691 = (n26207 & n26209) | (n26207 & n53690) | (n26209 & n53690);
  assign n53692 = n26200 | n53522;
  assign n53693 = (n26200 & n26202) | (n26200 & n53692) | (n26202 & n53692);
  assign n68746 = n26193 | n68642;
  assign n68747 = (n26193 & n26195) | (n26193 & n68746) | (n26195 & n68746);
  assign n26228 = n26186 | n26189;
  assign n26229 = n26179 | n26182;
  assign n26230 = n26172 | n26175;
  assign n26231 = n26165 | n26168;
  assign n26232 = n26158 | n26161;
  assign n53694 = n26151 | n26153;
  assign n53695 = (n25868 & n26151) | (n25868 & n53694) | (n26151 & n53694);
  assign n53696 = n26144 | n26146;
  assign n53697 = (n26144 & n53524) | (n26144 & n53696) | (n53524 & n53696);
  assign n53698 = n26137 | n26139;
  assign n53699 = (n26137 & n53526) | (n26137 & n53698) | (n53526 & n53698);
  assign n53700 = n26130 | n26132;
  assign n53701 = (n26130 & n53528) | (n26130 & n53700) | (n53528 & n53700);
  assign n53532 = (n25759 & n53369) | (n25759 & n53531) | (n53369 & n53531);
  assign n53534 = (n25752 & n53371) | (n25752 & n53533) | (n53371 & n53533);
  assign n53539 = (n68529 & n68644) | (n68529 & n53538) | (n68644 & n53538);
  assign n53711 = n26018 | n26020;
  assign n68748 = n25661 | n26018;
  assign n68749 = (n26018 & n26020) | (n26018 & n68748) | (n26020 & n68748);
  assign n68750 = (n53468 & n53711) | (n53468 & n68749) | (n53711 & n68749);
  assign n68751 = (n53467 & n53711) | (n53467 & n68749) | (n53711 & n68749);
  assign n68752 = (n53227 & n68750) | (n53227 & n68751) | (n68750 & n68751);
  assign n53716 = n25997 | n25999;
  assign n68753 = n25640 | n25997;
  assign n68754 = (n25997 & n25999) | (n25997 & n68753) | (n25999 & n68753);
  assign n68755 = (n53458 & n53716) | (n53458 & n68754) | (n53716 & n68754);
  assign n68756 = (n53457 & n53716) | (n53457 & n68754) | (n53716 & n68754);
  assign n68757 = (n68467 & n68755) | (n68467 & n68756) | (n68755 & n68756);
  assign n68760 = n25598 | n25955;
  assign n68761 = (n25955 & n25957) | (n25955 & n68760) | (n25957 & n68760);
  assign n68762 = n25955 | n25957;
  assign n68763 = (n25955 & n53555) | (n25955 & n68762) | (n53555 & n68762);
  assign n68764 = (n53392 & n68761) | (n53392 & n68763) | (n68761 & n68763);
  assign n68765 = (n68562 & n68761) | (n68562 & n68763) | (n68761 & n68763);
  assign n68766 = (n53073 & n68764) | (n53073 & n68765) | (n68764 & n68765);
  assign n53401 = (n68308 & n53399) | (n68308 & n53400) | (n53399 & n53400);
  assign n68771 = n25920 | n25922;
  assign n68772 = (n25920 & n68675) | (n25920 & n68771) | (n68675 & n68771);
  assign n68773 = (n25920 & n68677) | (n25920 & n68771) | (n68677 & n68771);
  assign n68774 = (n68484 & n68772) | (n68484 & n68773) | (n68772 & n68773);
  assign n68775 = (n68483 & n68772) | (n68483 & n68773) | (n68772 & n68773);
  assign n68776 = (n67914 & n68774) | (n67914 & n68775) | (n68774 & n68775);
  assign n26269 = x159 & x176;
  assign n26270 = x158 & x177;
  assign n26271 = n26269 & n26270;
  assign n26272 = n26269 | n26270;
  assign n26273 = ~n26271 & n26272;
  assign n68777 = n25906 | n68665;
  assign n68780 = n26273 & n68777;
  assign n68778 = n25906 | n25908;
  assign n68781 = n26273 & n68778;
  assign n68782 = (n68574 & n68780) | (n68574 & n68781) | (n68780 & n68781);
  assign n68784 = (n68576 & n68780) | (n68576 & n68781) | (n68780 & n68781);
  assign n53749 = (n68195 & n68782) | (n68195 & n68784) | (n68782 & n68784);
  assign n68785 = n26273 | n68777;
  assign n68786 = n26273 | n68778;
  assign n68787 = (n68574 & n68785) | (n68574 & n68786) | (n68785 & n68786);
  assign n68788 = (n68576 & n68785) | (n68576 & n68786) | (n68785 & n68786);
  assign n53752 = (n68195 & n68787) | (n68195 & n68788) | (n68787 & n68788);
  assign n26276 = ~n53749 & n53752;
  assign n26277 = x157 & x178;
  assign n26278 = n26276 & n26277;
  assign n26279 = n26276 | n26277;
  assign n26280 = ~n26278 & n26279;
  assign n68789 = n25913 | n25915;
  assign n68791 = n26280 & n68789;
  assign n68792 = n25913 & n26280;
  assign n68793 = (n68672 & n68791) | (n68672 & n68792) | (n68791 & n68792);
  assign n68795 = (n68673 & n68791) | (n68673 & n68792) | (n68791 & n68792);
  assign n53755 = (n68389 & n68793) | (n68389 & n68795) | (n68793 & n68795);
  assign n68796 = n26280 | n68789;
  assign n68797 = n25913 | n26280;
  assign n68798 = (n68672 & n68796) | (n68672 & n68797) | (n68796 & n68797);
  assign n68799 = (n68673 & n68796) | (n68673 & n68797) | (n68796 & n68797);
  assign n53758 = (n68389 & n68798) | (n68389 & n68799) | (n68798 & n68799);
  assign n26283 = ~n53755 & n53758;
  assign n26284 = x156 & x179;
  assign n26285 = n26283 & n26284;
  assign n26286 = n26283 | n26284;
  assign n26287 = ~n26285 & n26286;
  assign n26288 = n68776 & n26287;
  assign n26289 = n68776 | n26287;
  assign n26290 = ~n26288 & n26289;
  assign n26291 = x155 & x180;
  assign n26292 = n26290 & n26291;
  assign n26293 = n26290 | n26291;
  assign n26294 = ~n26292 & n26293;
  assign n53736 = n25927 | n25929;
  assign n53759 = n26294 & n53736;
  assign n53760 = n25927 & n26294;
  assign n68800 = (n53759 & n53760) | (n53759 & n68664) | (n53760 & n68664);
  assign n68801 = (n53759 & n53760) | (n53759 & n68663) | (n53760 & n68663);
  assign n68802 = (n68409 & n68800) | (n68409 & n68801) | (n68800 & n68801);
  assign n53762 = n26294 | n53736;
  assign n53763 = n25927 | n26294;
  assign n68803 = (n53762 & n53763) | (n53762 & n68664) | (n53763 & n68664);
  assign n68804 = (n53762 & n53763) | (n53762 & n68663) | (n53763 & n68663);
  assign n68805 = (n68409 & n68803) | (n68409 & n68804) | (n68803 & n68804);
  assign n26297 = ~n68802 & n68805;
  assign n26298 = x154 & x181;
  assign n26299 = n26297 & n26298;
  assign n26300 = n26297 | n26298;
  assign n26301 = ~n26299 & n26300;
  assign n68806 = n25934 | n25936;
  assign n68807 = (n25934 & n53562) | (n25934 & n68806) | (n53562 & n68806);
  assign n53765 = n26301 & n68807;
  assign n68808 = n25577 | n25934;
  assign n68809 = (n25934 & n25936) | (n25934 & n68808) | (n25936 & n68808);
  assign n53766 = n26301 & n68809;
  assign n53767 = (n53401 & n53765) | (n53401 & n53766) | (n53765 & n53766);
  assign n53768 = n26301 | n68807;
  assign n53769 = n26301 | n68809;
  assign n53770 = (n53401 & n53768) | (n53401 & n53769) | (n53768 & n53769);
  assign n26304 = ~n53767 & n53770;
  assign n26305 = x153 & x182;
  assign n26306 = n26304 & n26305;
  assign n26307 = n26304 | n26305;
  assign n26308 = ~n26306 & n26307;
  assign n68767 = n25941 | n25943;
  assign n68768 = (n25941 & n53560) | (n25941 & n68767) | (n53560 & n68767);
  assign n68810 = n26308 & n68768;
  assign n68769 = n25584 | n25941;
  assign n68770 = (n25941 & n25943) | (n25941 & n68769) | (n25943 & n68769);
  assign n68811 = n26308 & n68770;
  assign n68812 = (n68569 & n68810) | (n68569 & n68811) | (n68810 & n68811);
  assign n68813 = n26308 | n68768;
  assign n68814 = n26308 | n68770;
  assign n68815 = (n68569 & n68813) | (n68569 & n68814) | (n68813 & n68814);
  assign n26311 = ~n68812 & n68815;
  assign n26312 = x152 & x183;
  assign n26313 = n26311 & n26312;
  assign n26314 = n26311 | n26312;
  assign n26315 = ~n26313 & n26314;
  assign n53728 = n25948 | n25950;
  assign n53771 = n26315 & n53728;
  assign n53772 = n25948 & n26315;
  assign n68816 = (n53558 & n53771) | (n53558 & n53772) | (n53771 & n53772);
  assign n68817 = (n53771 & n53772) | (n53771 & n68661) | (n53772 & n68661);
  assign n68818 = (n68479 & n68816) | (n68479 & n68817) | (n68816 & n68817);
  assign n53774 = n26315 | n53728;
  assign n53775 = n25948 | n26315;
  assign n68819 = (n53558 & n53774) | (n53558 & n53775) | (n53774 & n53775);
  assign n68820 = (n53774 & n53775) | (n53774 & n68661) | (n53775 & n68661);
  assign n68821 = (n68479 & n68819) | (n68479 & n68820) | (n68819 & n68820);
  assign n26318 = ~n68818 & n68821;
  assign n26319 = x151 & x184;
  assign n26320 = n26318 & n26319;
  assign n26321 = n26318 | n26319;
  assign n26322 = ~n26320 & n26321;
  assign n26323 = n68766 & n26322;
  assign n26324 = n68766 | n26322;
  assign n26325 = ~n26323 & n26324;
  assign n26326 = x150 & x185;
  assign n26327 = n26325 & n26326;
  assign n26328 = n26325 | n26326;
  assign n26329 = ~n26327 & n26328;
  assign n53723 = n25962 | n25964;
  assign n53777 = n26329 & n53723;
  assign n53778 = n25962 & n26329;
  assign n53779 = (n68659 & n53777) | (n68659 & n53778) | (n53777 & n53778);
  assign n53780 = n26329 | n53723;
  assign n53781 = n25962 | n26329;
  assign n53782 = (n68659 & n53780) | (n68659 & n53781) | (n53780 & n53781);
  assign n26332 = ~n53779 & n53782;
  assign n26333 = x149 & x186;
  assign n26334 = n26332 & n26333;
  assign n26335 = n26332 | n26333;
  assign n26336 = ~n26334 & n26335;
  assign n53783 = n25969 & n26336;
  assign n68822 = (n26336 & n53613) | (n26336 & n53783) | (n53613 & n53783);
  assign n68823 = (n26336 & n53612) | (n26336 & n53783) | (n53612 & n53783);
  assign n68824 = (n53390 & n68822) | (n53390 & n68823) | (n68822 & n68823);
  assign n53785 = n25969 | n26336;
  assign n68825 = n53613 | n53785;
  assign n68826 = n53612 | n53785;
  assign n68827 = (n53390 & n68825) | (n53390 & n68826) | (n68825 & n68826);
  assign n26339 = ~n68824 & n68827;
  assign n26340 = x148 & x187;
  assign n26341 = n26339 & n26340;
  assign n26342 = n26339 | n26340;
  assign n26343 = ~n26341 & n26342;
  assign n53721 = n25976 | n25978;
  assign n68828 = n26343 & n53721;
  assign n68758 = n25619 | n25976;
  assign n68759 = (n25976 & n25978) | (n25976 & n68758) | (n25978 & n68758);
  assign n68829 = n26343 & n68759;
  assign n68830 = (n53449 & n68828) | (n53449 & n68829) | (n68828 & n68829);
  assign n68831 = n26343 | n53721;
  assign n68832 = n26343 | n68759;
  assign n68833 = (n53449 & n68831) | (n53449 & n68832) | (n68831 & n68832);
  assign n26346 = ~n68830 & n68833;
  assign n26347 = x147 & x188;
  assign n26348 = n26346 & n26347;
  assign n26349 = n26346 | n26347;
  assign n26350 = ~n26348 & n26349;
  assign n53718 = n25983 | n25985;
  assign n53787 = n26350 & n53718;
  assign n53788 = n25983 & n26350;
  assign n53789 = (n68654 & n53787) | (n68654 & n53788) | (n53787 & n53788);
  assign n53790 = n26350 | n53718;
  assign n53791 = n25983 | n26350;
  assign n53792 = (n68654 & n53790) | (n68654 & n53791) | (n53790 & n53791);
  assign n26353 = ~n53789 & n53792;
  assign n26354 = x146 & x189;
  assign n26355 = n26353 & n26354;
  assign n26356 = n26353 | n26354;
  assign n26357 = ~n26355 & n26356;
  assign n53793 = n25990 & n26357;
  assign n68834 = (n26357 & n53623) | (n26357 & n53793) | (n53623 & n53793);
  assign n68835 = (n26357 & n53622) | (n26357 & n53793) | (n53622 & n53793);
  assign n68836 = (n68558 & n68834) | (n68558 & n68835) | (n68834 & n68835);
  assign n53795 = n25990 | n26357;
  assign n68837 = n53623 | n53795;
  assign n68838 = n53622 | n53795;
  assign n68839 = (n68558 & n68837) | (n68558 & n68838) | (n68837 & n68838);
  assign n26360 = ~n68836 & n68839;
  assign n26361 = x145 & x190;
  assign n26362 = n26360 & n26361;
  assign n26363 = n26360 | n26361;
  assign n26364 = ~n26362 & n26363;
  assign n26365 = n68757 & n26364;
  assign n26366 = n68757 | n26364;
  assign n26367 = ~n26365 & n26366;
  assign n26368 = x144 & x191;
  assign n26369 = n26367 & n26368;
  assign n26370 = n26367 | n26368;
  assign n26371 = ~n26369 & n26370;
  assign n53713 = n26004 | n26006;
  assign n53797 = n26371 & n53713;
  assign n53798 = n26004 & n26371;
  assign n53799 = (n68649 & n53797) | (n68649 & n53798) | (n53797 & n53798);
  assign n53800 = n26371 | n53713;
  assign n53801 = n26004 | n26371;
  assign n53802 = (n68649 & n53800) | (n68649 & n53801) | (n53800 & n53801);
  assign n26374 = ~n53799 & n53802;
  assign n26375 = x143 & x192;
  assign n26376 = n26374 & n26375;
  assign n26377 = n26374 | n26375;
  assign n26378 = ~n26376 & n26377;
  assign n53803 = n26011 & n26378;
  assign n68840 = (n26378 & n53633) | (n26378 & n53803) | (n53633 & n53803);
  assign n68841 = (n26378 & n53632) | (n26378 & n53803) | (n53632 & n53803);
  assign n68842 = (n68553 & n68840) | (n68553 & n68841) | (n68840 & n68841);
  assign n53805 = n26011 | n26378;
  assign n68843 = n53633 | n53805;
  assign n68844 = n53632 | n53805;
  assign n68845 = (n68553 & n68843) | (n68553 & n68844) | (n68843 & n68844);
  assign n26381 = ~n68842 & n68845;
  assign n26382 = x142 & x193;
  assign n26383 = n26381 & n26382;
  assign n26384 = n26381 | n26382;
  assign n26385 = ~n26383 & n26384;
  assign n26386 = n68752 & n26385;
  assign n26387 = n68752 | n26385;
  assign n26388 = ~n26386 & n26387;
  assign n26389 = x141 & x194;
  assign n26390 = n26388 & n26389;
  assign n26391 = n26388 | n26389;
  assign n26392 = ~n26390 & n26391;
  assign n53708 = n26025 | n26027;
  assign n53807 = n26392 & n53708;
  assign n53808 = n26025 & n26392;
  assign n53809 = (n53539 & n53807) | (n53539 & n53808) | (n53807 & n53808);
  assign n53810 = n26392 | n53708;
  assign n53811 = n26025 | n26392;
  assign n53812 = (n53539 & n53810) | (n53539 & n53811) | (n53810 & n53811);
  assign n26395 = ~n53809 & n53812;
  assign n26396 = x140 & x195;
  assign n26397 = n26395 & n26396;
  assign n26398 = n26395 | n26396;
  assign n26399 = ~n26397 & n26398;
  assign n53813 = n26032 & n26399;
  assign n53814 = (n26399 & n68728) | (n26399 & n53813) | (n68728 & n53813);
  assign n53815 = n26032 | n26399;
  assign n53816 = n68728 | n53815;
  assign n26402 = ~n53814 & n53816;
  assign n26403 = x139 & x196;
  assign n26404 = n26402 & n26403;
  assign n26405 = n26402 | n26403;
  assign n26406 = ~n26404 & n26405;
  assign n53817 = n26039 & n26406;
  assign n53818 = (n26406 & n53647) | (n26406 & n53817) | (n53647 & n53817);
  assign n53819 = n26039 | n26406;
  assign n53820 = n53647 | n53819;
  assign n26409 = ~n53818 & n53820;
  assign n26410 = x138 & x197;
  assign n26411 = n26409 & n26410;
  assign n26412 = n26409 | n26410;
  assign n26413 = ~n26411 & n26412;
  assign n53821 = n26046 & n26413;
  assign n53822 = (n26413 & n53651) | (n26413 & n53821) | (n53651 & n53821);
  assign n53823 = n26046 | n26413;
  assign n53824 = n53651 | n53823;
  assign n26416 = ~n53822 & n53824;
  assign n26417 = x137 & x198;
  assign n26418 = n26416 & n26417;
  assign n26419 = n26416 | n26417;
  assign n26420 = ~n26418 & n26419;
  assign n53825 = n26053 & n26420;
  assign n53826 = (n26420 & n53655) | (n26420 & n53825) | (n53655 & n53825);
  assign n53827 = n26053 | n26420;
  assign n53828 = n53655 | n53827;
  assign n26423 = ~n53826 & n53828;
  assign n26424 = x136 & x199;
  assign n26425 = n26423 & n26424;
  assign n26426 = n26423 | n26424;
  assign n26427 = ~n26425 & n26426;
  assign n53829 = n26060 & n26427;
  assign n53830 = (n26427 & n53659) | (n26427 & n53829) | (n53659 & n53829);
  assign n53831 = n26060 | n26427;
  assign n53832 = n53659 | n53831;
  assign n26430 = ~n53830 & n53832;
  assign n26431 = x135 & x200;
  assign n26432 = n26430 & n26431;
  assign n26433 = n26430 | n26431;
  assign n26434 = ~n26432 & n26433;
  assign n53833 = n26067 & n26434;
  assign n53834 = (n26434 & n53663) | (n26434 & n53833) | (n53663 & n53833);
  assign n53835 = n26067 | n26434;
  assign n53836 = n53663 | n53835;
  assign n26437 = ~n53834 & n53836;
  assign n26438 = x134 & x201;
  assign n26439 = n26437 & n26438;
  assign n26440 = n26437 | n26438;
  assign n26441 = ~n26439 & n26440;
  assign n53837 = n26074 & n26441;
  assign n53838 = (n26441 & n53667) | (n26441 & n53837) | (n53667 & n53837);
  assign n53839 = n26074 | n26441;
  assign n53840 = n53667 | n53839;
  assign n26444 = ~n53838 & n53840;
  assign n26445 = x133 & x202;
  assign n26446 = n26444 & n26445;
  assign n26447 = n26444 | n26445;
  assign n26448 = ~n26446 & n26447;
  assign n53841 = n26081 & n26448;
  assign n53842 = (n26448 & n53671) | (n26448 & n53841) | (n53671 & n53841);
  assign n53843 = n26081 | n26448;
  assign n53844 = n53671 | n53843;
  assign n26451 = ~n53842 & n53844;
  assign n26452 = x132 & x203;
  assign n26453 = n26451 & n26452;
  assign n26454 = n26451 | n26452;
  assign n26455 = ~n26453 & n26454;
  assign n53845 = n26088 & n26455;
  assign n53846 = (n26455 & n53675) | (n26455 & n53845) | (n53675 & n53845);
  assign n53847 = n26088 | n26455;
  assign n53848 = n53675 | n53847;
  assign n26458 = ~n53846 & n53848;
  assign n26459 = x131 & x204;
  assign n26460 = n26458 & n26459;
  assign n26461 = n26458 | n26459;
  assign n26462 = ~n26460 & n26461;
  assign n53849 = n26095 & n26462;
  assign n53850 = (n26462 & n53679) | (n26462 & n53849) | (n53679 & n53849);
  assign n53851 = n26095 | n26462;
  assign n53852 = n53679 | n53851;
  assign n26465 = ~n53850 & n53852;
  assign n26466 = x130 & x205;
  assign n26467 = n26465 & n26466;
  assign n26468 = n26465 | n26466;
  assign n26469 = ~n26467 & n26468;
  assign n53853 = n26102 & n26469;
  assign n53854 = (n26469 & n53684) | (n26469 & n53853) | (n53684 & n53853);
  assign n53855 = n26102 | n26469;
  assign n53856 = n53684 | n53855;
  assign n26472 = ~n53854 & n53856;
  assign n26473 = x129 & x206;
  assign n26474 = n26472 & n26473;
  assign n26475 = n26472 | n26473;
  assign n26476 = ~n26474 & n26475;
  assign n53706 = n26109 | n26111;
  assign n53857 = n26476 & n53706;
  assign n53858 = n26109 & n26476;
  assign n53859 = (n53534 & n53857) | (n53534 & n53858) | (n53857 & n53858);
  assign n53860 = n26476 | n53706;
  assign n53861 = n26109 | n26476;
  assign n53862 = (n53534 & n53860) | (n53534 & n53861) | (n53860 & n53861);
  assign n26479 = ~n53859 & n53862;
  assign n26480 = x128 & x207;
  assign n26481 = n26479 & n26480;
  assign n26482 = n26479 | n26480;
  assign n26483 = ~n26481 & n26482;
  assign n53704 = n26116 | n26118;
  assign n68846 = n26483 & n53704;
  assign n68847 = n26116 & n26483;
  assign n68848 = (n53532 & n68846) | (n53532 & n68847) | (n68846 & n68847);
  assign n68849 = n26483 | n53704;
  assign n68850 = n26116 | n26483;
  assign n68851 = (n53532 & n68849) | (n53532 & n68850) | (n68849 & n68850);
  assign n26486 = ~n68848 & n68851;
  assign n26487 = x127 & x208;
  assign n26488 = n26486 & n26487;
  assign n26489 = n26486 | n26487;
  assign n26490 = ~n26488 & n26489;
  assign n53702 = n26123 | n26125;
  assign n68852 = n26490 & n53702;
  assign n68853 = n26123 & n26490;
  assign n68854 = (n53530 & n68852) | (n53530 & n68853) | (n68852 & n68853);
  assign n68855 = n26490 | n53702;
  assign n68856 = n26123 | n26490;
  assign n68857 = (n53530 & n68855) | (n53530 & n68856) | (n68855 & n68856);
  assign n26493 = ~n68854 & n68857;
  assign n26494 = x126 & x209;
  assign n26495 = n26493 & n26494;
  assign n26496 = n26493 | n26494;
  assign n26497 = ~n26495 & n26496;
  assign n26498 = n53701 & n26497;
  assign n26499 = n53701 | n26497;
  assign n26500 = ~n26498 & n26499;
  assign n26501 = x125 & x210;
  assign n26502 = n26500 & n26501;
  assign n26503 = n26500 | n26501;
  assign n26504 = ~n26502 & n26503;
  assign n26505 = n53699 & n26504;
  assign n26506 = n53699 | n26504;
  assign n26507 = ~n26505 & n26506;
  assign n26508 = x124 & x211;
  assign n26509 = n26507 & n26508;
  assign n26510 = n26507 | n26508;
  assign n26511 = ~n26509 & n26510;
  assign n26512 = n53697 & n26511;
  assign n26513 = n53697 | n26511;
  assign n26514 = ~n26512 & n26513;
  assign n26515 = x123 & x212;
  assign n26516 = n26514 & n26515;
  assign n26517 = n26514 | n26515;
  assign n26518 = ~n26516 & n26517;
  assign n26519 = n53695 & n26518;
  assign n26520 = n53695 | n26518;
  assign n26521 = ~n26519 & n26520;
  assign n26522 = x122 & x213;
  assign n26523 = n26521 & n26522;
  assign n26524 = n26521 | n26522;
  assign n26525 = ~n26523 & n26524;
  assign n26526 = n26232 & n26525;
  assign n26527 = n26232 | n26525;
  assign n26528 = ~n26526 & n26527;
  assign n26529 = x121 & x214;
  assign n26530 = n26528 & n26529;
  assign n26531 = n26528 | n26529;
  assign n26532 = ~n26530 & n26531;
  assign n26533 = n26231 & n26532;
  assign n26534 = n26231 | n26532;
  assign n26535 = ~n26533 & n26534;
  assign n26536 = x120 & x215;
  assign n26537 = n26535 & n26536;
  assign n26538 = n26535 | n26536;
  assign n26539 = ~n26537 & n26538;
  assign n26540 = n26230 & n26539;
  assign n26541 = n26230 | n26539;
  assign n26542 = ~n26540 & n26541;
  assign n26543 = x119 & x216;
  assign n26544 = n26542 & n26543;
  assign n26545 = n26542 | n26543;
  assign n26546 = ~n26544 & n26545;
  assign n26547 = n26229 & n26546;
  assign n26548 = n26229 | n26546;
  assign n26549 = ~n26547 & n26548;
  assign n26550 = x118 & x217;
  assign n26551 = n26549 & n26550;
  assign n26552 = n26549 | n26550;
  assign n26553 = ~n26551 & n26552;
  assign n26554 = n26228 & n26553;
  assign n26555 = n26228 | n26553;
  assign n26556 = ~n26554 & n26555;
  assign n26557 = x117 & x218;
  assign n26558 = n26556 & n26557;
  assign n26559 = n26556 | n26557;
  assign n26560 = ~n26558 & n26559;
  assign n26561 = n68747 & n26560;
  assign n26562 = n68747 | n26560;
  assign n26563 = ~n26561 & n26562;
  assign n26564 = x116 & x219;
  assign n26565 = n26563 & n26564;
  assign n26566 = n26563 | n26564;
  assign n26567 = ~n26565 & n26566;
  assign n26568 = n53693 & n26567;
  assign n26569 = n53693 | n26567;
  assign n26570 = ~n26568 & n26569;
  assign n26571 = x115 & x220;
  assign n26572 = n26570 & n26571;
  assign n26573 = n26570 | n26571;
  assign n26574 = ~n26572 & n26573;
  assign n26575 = n53691 & n26574;
  assign n26576 = n53691 | n26574;
  assign n26577 = ~n26575 & n26576;
  assign n26578 = x114 & x221;
  assign n26579 = n26577 & n26578;
  assign n26580 = n26577 | n26578;
  assign n26581 = ~n26579 & n26580;
  assign n26582 = n53689 & n26581;
  assign n26583 = n53689 | n26581;
  assign n26584 = ~n26582 & n26583;
  assign n26585 = x113 & x222;
  assign n26586 = n26584 & n26585;
  assign n26587 = n26584 | n26585;
  assign n26588 = ~n26586 & n26587;
  assign n26589 = n26221 & n26588;
  assign n26590 = n26221 | n26588;
  assign n26591 = ~n26589 & n26590;
  assign n26592 = x112 & x223;
  assign n26593 = n26591 & n26592;
  assign n26594 = n26591 | n26592;
  assign n26595 = ~n26593 & n26594;
  assign n68858 = n26221 | n26585;
  assign n68859 = (n26221 & n26584) | (n26221 & n68858) | (n26584 & n68858);
  assign n53864 = (n26586 & n26588) | (n26586 & n68859) | (n26588 & n68859);
  assign n53865 = n26579 | n53689;
  assign n53866 = (n26579 & n26581) | (n26579 & n53865) | (n26581 & n53865);
  assign n53867 = n26572 | n53691;
  assign n53868 = (n26572 & n26574) | (n26572 & n53867) | (n26574 & n53867);
  assign n53869 = n26565 | n53693;
  assign n53870 = (n26565 & n26567) | (n26565 & n53869) | (n26567 & n53869);
  assign n68860 = n26558 | n68747;
  assign n68861 = (n26558 & n26560) | (n26558 & n68860) | (n26560 & n68860);
  assign n26601 = n26551 | n26554;
  assign n26602 = n26544 | n26547;
  assign n26603 = n26537 | n26540;
  assign n26604 = n26530 | n26533;
  assign n53871 = n26523 | n26525;
  assign n53872 = (n26232 & n26523) | (n26232 & n53871) | (n26523 & n53871);
  assign n53873 = n26516 | n26518;
  assign n53874 = (n26516 & n53695) | (n26516 & n53873) | (n53695 & n53873);
  assign n53875 = n26509 | n26511;
  assign n53876 = (n26509 & n53697) | (n26509 & n53875) | (n53697 & n53875);
  assign n53877 = n26502 | n26504;
  assign n53878 = (n26502 & n53699) | (n26502 & n53877) | (n53699 & n53877);
  assign n53703 = (n26123 & n53530) | (n26123 & n53702) | (n53530 & n53702);
  assign n53705 = (n26116 & n53532) | (n26116 & n53704) | (n53532 & n53704);
  assign n53891 = n26376 | n26378;
  assign n68864 = n26011 | n26376;
  assign n68865 = (n26376 & n26378) | (n26376 & n68864) | (n26378 & n68864);
  assign n68866 = (n53633 & n53891) | (n53633 & n68865) | (n53891 & n68865);
  assign n68867 = (n53632 & n53891) | (n53632 & n68865) | (n53891 & n68865);
  assign n68868 = (n68553 & n68866) | (n68553 & n68867) | (n68866 & n68867);
  assign n53896 = n26355 | n26357;
  assign n68869 = n25990 | n26355;
  assign n68870 = (n26355 & n26357) | (n26355 & n68869) | (n26357 & n68869);
  assign n68871 = (n53623 & n53896) | (n53623 & n68870) | (n53896 & n68870);
  assign n68872 = (n53622 & n53896) | (n53622 & n68870) | (n53896 & n68870);
  assign n68873 = (n68558 & n68871) | (n68558 & n68872) | (n68871 & n68872);
  assign n53722 = (n53449 & n68759) | (n53449 & n53721) | (n68759 & n53721);
  assign n53901 = n26334 | n26336;
  assign n68874 = n25969 | n26334;
  assign n68875 = (n26334 & n26336) | (n26334 & n68874) | (n26336 & n68874);
  assign n68876 = (n53613 & n53901) | (n53613 & n68875) | (n53901 & n68875);
  assign n68877 = (n53612 & n53901) | (n53612 & n68875) | (n53901 & n68875);
  assign n68878 = (n53390 & n68876) | (n53390 & n68877) | (n68876 & n68877);
  assign n68879 = n25962 | n26327;
  assign n68880 = (n26327 & n26329) | (n26327 & n68879) | (n26329 & n68879);
  assign n53904 = n26327 | n53777;
  assign n53905 = (n68659 & n68880) | (n68659 & n53904) | (n68880 & n53904);
  assign n68881 = n25948 | n26313;
  assign n68882 = (n26313 & n26315) | (n26313 & n68881) | (n26315 & n68881);
  assign n68883 = n26313 | n26315;
  assign n68884 = (n26313 & n53728) | (n26313 & n68883) | (n53728 & n68883);
  assign n68885 = (n53558 & n68882) | (n53558 & n68884) | (n68882 & n68884);
  assign n68886 = (n68661 & n68882) | (n68661 & n68884) | (n68882 & n68884);
  assign n68887 = (n68479 & n68885) | (n68479 & n68886) | (n68885 & n68886);
  assign n26642 = x160 & x176;
  assign n26643 = x159 & x177;
  assign n26644 = n26642 & n26643;
  assign n26645 = n26642 | n26643;
  assign n26646 = ~n26644 & n26645;
  assign n53919 = n26271 | n68784;
  assign n68888 = n26646 & n53919;
  assign n53918 = n26271 | n68782;
  assign n68889 = n26646 & n53918;
  assign n68890 = (n68195 & n68888) | (n68195 & n68889) | (n68888 & n68889);
  assign n68891 = n26646 | n53919;
  assign n68892 = n26646 | n53918;
  assign n68893 = (n68195 & n68891) | (n68195 & n68892) | (n68891 & n68892);
  assign n26649 = ~n68890 & n68893;
  assign n26650 = x158 & x178;
  assign n26651 = n26649 & n26650;
  assign n26652 = n26649 | n26650;
  assign n26653 = ~n26651 & n26652;
  assign n53921 = n26278 & n26653;
  assign n68894 = (n26653 & n53921) | (n26653 & n68795) | (n53921 & n68795);
  assign n68895 = (n26653 & n53921) | (n26653 & n68793) | (n53921 & n68793);
  assign n68896 = (n68389 & n68894) | (n68389 & n68895) | (n68894 & n68895);
  assign n53923 = n26278 | n26653;
  assign n68897 = n53923 | n68795;
  assign n68898 = n53923 | n68793;
  assign n68899 = (n68389 & n68897) | (n68389 & n68898) | (n68897 & n68898);
  assign n26656 = ~n68896 & n68899;
  assign n26657 = x157 & x179;
  assign n26658 = n26656 & n26657;
  assign n26659 = n26656 | n26657;
  assign n26660 = ~n26658 & n26659;
  assign n53916 = n26285 | n26287;
  assign n53925 = n26660 & n53916;
  assign n53926 = n26285 & n26660;
  assign n53927 = (n68776 & n53925) | (n68776 & n53926) | (n53925 & n53926);
  assign n53928 = n26660 | n53916;
  assign n53929 = n26285 | n26660;
  assign n53930 = (n68776 & n53928) | (n68776 & n53929) | (n53928 & n53929);
  assign n26663 = ~n53927 & n53930;
  assign n26664 = x156 & x180;
  assign n26665 = n26663 & n26664;
  assign n26666 = n26663 | n26664;
  assign n26667 = ~n26665 & n26666;
  assign n68902 = n25927 | n26292;
  assign n68903 = (n26292 & n26294) | (n26292 & n68902) | (n26294 & n68902);
  assign n53932 = n26667 & n68903;
  assign n68900 = n26292 & n26667;
  assign n68901 = (n26667 & n53759) | (n26667 & n68900) | (n53759 & n68900);
  assign n68904 = (n53932 & n68664) | (n53932 & n68901) | (n68664 & n68901);
  assign n68905 = (n53932 & n68663) | (n53932 & n68901) | (n68663 & n68901);
  assign n68906 = (n68409 & n68904) | (n68409 & n68905) | (n68904 & n68905);
  assign n53935 = n26667 | n68903;
  assign n68907 = n26292 | n26667;
  assign n68908 = n53759 | n68907;
  assign n68909 = (n53935 & n68664) | (n53935 & n68908) | (n68664 & n68908);
  assign n68910 = (n53935 & n68663) | (n53935 & n68908) | (n68663 & n68908);
  assign n68911 = (n68409 & n68909) | (n68409 & n68910) | (n68909 & n68910);
  assign n26670 = ~n68906 & n68911;
  assign n26671 = x155 & x181;
  assign n26672 = n26670 & n26671;
  assign n26673 = n26670 | n26671;
  assign n26674 = ~n26672 & n26673;
  assign n53937 = n26299 & n26674;
  assign n68912 = (n26674 & n53765) | (n26674 & n53937) | (n53765 & n53937);
  assign n68913 = (n26674 & n53766) | (n26674 & n53937) | (n53766 & n53937);
  assign n68914 = (n53401 & n68912) | (n53401 & n68913) | (n68912 & n68913);
  assign n53939 = n26299 | n26674;
  assign n68915 = n53765 | n53939;
  assign n68916 = n53766 | n53939;
  assign n68917 = (n53401 & n68915) | (n53401 & n68916) | (n68915 & n68916);
  assign n26677 = ~n68914 & n68917;
  assign n26678 = x154 & x182;
  assign n26679 = n26677 & n26678;
  assign n26680 = n26677 | n26678;
  assign n26681 = ~n26679 & n26680;
  assign n53911 = n26306 | n26308;
  assign n53941 = n26681 & n53911;
  assign n53942 = n26306 & n26681;
  assign n68918 = (n53941 & n53942) | (n53941 & n68768) | (n53942 & n68768);
  assign n68919 = (n53941 & n53942) | (n53941 & n68770) | (n53942 & n68770);
  assign n68920 = (n68569 & n68918) | (n68569 & n68919) | (n68918 & n68919);
  assign n53944 = n26681 | n53911;
  assign n53945 = n26306 | n26681;
  assign n68921 = (n53944 & n53945) | (n53944 & n68768) | (n53945 & n68768);
  assign n68922 = (n53944 & n53945) | (n53944 & n68770) | (n53945 & n68770);
  assign n68923 = (n68569 & n68921) | (n68569 & n68922) | (n68921 & n68922);
  assign n26684 = ~n68920 & n68923;
  assign n26685 = x153 & x183;
  assign n26686 = n26684 & n26685;
  assign n26687 = n26684 | n26685;
  assign n26688 = ~n26686 & n26687;
  assign n26689 = n68887 & n26688;
  assign n26690 = n68887 | n26688;
  assign n26691 = ~n26689 & n26690;
  assign n26692 = x152 & x184;
  assign n26693 = n26691 & n26692;
  assign n26694 = n26691 | n26692;
  assign n26695 = ~n26693 & n26694;
  assign n53906 = n26320 | n26322;
  assign n53947 = n26695 & n53906;
  assign n53948 = n26320 & n26695;
  assign n53949 = (n68766 & n53947) | (n68766 & n53948) | (n53947 & n53948);
  assign n53950 = n26695 | n53906;
  assign n53951 = n26320 | n26695;
  assign n53952 = (n68766 & n53950) | (n68766 & n53951) | (n53950 & n53951);
  assign n26698 = ~n53949 & n53952;
  assign n26699 = x151 & x185;
  assign n26700 = n26698 & n26699;
  assign n26701 = n26698 | n26699;
  assign n26702 = ~n26700 & n26701;
  assign n26703 = n53905 & n26702;
  assign n26704 = n53905 | n26702;
  assign n26705 = ~n26703 & n26704;
  assign n26706 = x150 & x186;
  assign n26707 = n26705 & n26706;
  assign n26708 = n26705 | n26706;
  assign n26709 = ~n26707 & n26708;
  assign n26710 = n68878 & n26709;
  assign n26711 = n68878 | n26709;
  assign n26712 = ~n26710 & n26711;
  assign n26713 = x149 & x187;
  assign n26714 = n26712 & n26713;
  assign n26715 = n26712 | n26713;
  assign n26716 = ~n26714 & n26715;
  assign n53898 = n26341 | n26343;
  assign n53953 = n26716 & n53898;
  assign n53954 = n26341 & n26716;
  assign n53955 = (n53722 & n53953) | (n53722 & n53954) | (n53953 & n53954);
  assign n53956 = n26716 | n53898;
  assign n53957 = n26341 | n26716;
  assign n53958 = (n53722 & n53956) | (n53722 & n53957) | (n53956 & n53957);
  assign n26719 = ~n53955 & n53958;
  assign n26720 = x148 & x188;
  assign n26721 = n26719 & n26720;
  assign n26722 = n26719 | n26720;
  assign n26723 = ~n26721 & n26722;
  assign n53959 = n26348 & n26723;
  assign n53960 = (n26723 & n53789) | (n26723 & n53959) | (n53789 & n53959);
  assign n53961 = n26348 | n26723;
  assign n53962 = n53789 | n53961;
  assign n26726 = ~n53960 & n53962;
  assign n26727 = x147 & x189;
  assign n26728 = n26726 & n26727;
  assign n26729 = n26726 | n26727;
  assign n26730 = ~n26728 & n26729;
  assign n26731 = n68873 & n26730;
  assign n26732 = n68873 | n26730;
  assign n26733 = ~n26731 & n26732;
  assign n26734 = x146 & x190;
  assign n26735 = n26733 & n26734;
  assign n26736 = n26733 | n26734;
  assign n26737 = ~n26735 & n26736;
  assign n53893 = n26362 | n26364;
  assign n53963 = n26737 & n53893;
  assign n53964 = n26362 & n26737;
  assign n53965 = (n68757 & n53963) | (n68757 & n53964) | (n53963 & n53964);
  assign n53966 = n26737 | n53893;
  assign n53967 = n26362 | n26737;
  assign n53968 = (n68757 & n53966) | (n68757 & n53967) | (n53966 & n53967);
  assign n26740 = ~n53965 & n53968;
  assign n26741 = x145 & x191;
  assign n26742 = n26740 & n26741;
  assign n26743 = n26740 | n26741;
  assign n26744 = ~n26742 & n26743;
  assign n53969 = n26369 & n26744;
  assign n68924 = (n26744 & n53798) | (n26744 & n53969) | (n53798 & n53969);
  assign n68925 = (n26744 & n53797) | (n26744 & n53969) | (n53797 & n53969);
  assign n68926 = (n68649 & n68924) | (n68649 & n68925) | (n68924 & n68925);
  assign n53971 = n26369 | n26744;
  assign n68927 = n53798 | n53971;
  assign n68928 = n53797 | n53971;
  assign n68929 = (n68649 & n68927) | (n68649 & n68928) | (n68927 & n68928);
  assign n26747 = ~n68926 & n68929;
  assign n26748 = x144 & x192;
  assign n26749 = n26747 & n26748;
  assign n26750 = n26747 | n26748;
  assign n26751 = ~n26749 & n26750;
  assign n26752 = n68868 & n26751;
  assign n26753 = n68868 | n26751;
  assign n26754 = ~n26752 & n26753;
  assign n26755 = x143 & x193;
  assign n26756 = n26754 & n26755;
  assign n26757 = n26754 | n26755;
  assign n26758 = ~n26756 & n26757;
  assign n53888 = n26383 | n26385;
  assign n53973 = n26758 & n53888;
  assign n53974 = n26383 & n26758;
  assign n53975 = (n68752 & n53973) | (n68752 & n53974) | (n53973 & n53974);
  assign n53976 = n26758 | n53888;
  assign n53977 = n26383 | n26758;
  assign n53978 = (n68752 & n53976) | (n68752 & n53977) | (n53976 & n53977);
  assign n26761 = ~n53975 & n53978;
  assign n26762 = x142 & x194;
  assign n26763 = n26761 & n26762;
  assign n26764 = n26761 | n26762;
  assign n26765 = ~n26763 & n26764;
  assign n53979 = n26390 & n26765;
  assign n68930 = (n26765 & n53808) | (n26765 & n53979) | (n53808 & n53979);
  assign n68931 = (n26765 & n53807) | (n26765 & n53979) | (n53807 & n53979);
  assign n68932 = (n53539 & n68930) | (n53539 & n68931) | (n68930 & n68931);
  assign n53981 = n26390 | n26765;
  assign n68933 = n53808 | n53981;
  assign n68934 = n53807 | n53981;
  assign n68935 = (n53539 & n68933) | (n53539 & n68934) | (n68933 & n68934);
  assign n26768 = ~n68932 & n68935;
  assign n26769 = x141 & x195;
  assign n26770 = n26768 & n26769;
  assign n26771 = n26768 | n26769;
  assign n26772 = ~n26770 & n26771;
  assign n53886 = n26397 | n26399;
  assign n68936 = n26772 & n53886;
  assign n68862 = n26032 | n26397;
  assign n68863 = (n26397 & n26399) | (n26397 & n68862) | (n26399 & n68862);
  assign n68937 = n26772 & n68863;
  assign n68938 = (n68728 & n68936) | (n68728 & n68937) | (n68936 & n68937);
  assign n68939 = n26772 | n53886;
  assign n68940 = n26772 | n68863;
  assign n68941 = (n68728 & n68939) | (n68728 & n68940) | (n68939 & n68940);
  assign n26775 = ~n68938 & n68941;
  assign n26776 = x140 & x196;
  assign n26777 = n26775 & n26776;
  assign n26778 = n26775 | n26776;
  assign n26779 = ~n26777 & n26778;
  assign n53983 = n26404 & n26779;
  assign n68942 = (n26779 & n53817) | (n26779 & n53983) | (n53817 & n53983);
  assign n68943 = (n26406 & n26779) | (n26406 & n53983) | (n26779 & n53983);
  assign n68944 = (n53647 & n68942) | (n53647 & n68943) | (n68942 & n68943);
  assign n53985 = n26404 | n26779;
  assign n68945 = n53817 | n53985;
  assign n68946 = n26406 | n53985;
  assign n68947 = (n53647 & n68945) | (n53647 & n68946) | (n68945 & n68946);
  assign n26782 = ~n68944 & n68947;
  assign n26783 = x139 & x197;
  assign n26784 = n26782 & n26783;
  assign n26785 = n26782 | n26783;
  assign n26786 = ~n26784 & n26785;
  assign n53987 = n26411 & n26786;
  assign n53988 = (n26786 & n53822) | (n26786 & n53987) | (n53822 & n53987);
  assign n53989 = n26411 | n26786;
  assign n53990 = n53822 | n53989;
  assign n26789 = ~n53988 & n53990;
  assign n26790 = x138 & x198;
  assign n26791 = n26789 & n26790;
  assign n26792 = n26789 | n26790;
  assign n26793 = ~n26791 & n26792;
  assign n53991 = n26418 & n26793;
  assign n53992 = (n26793 & n53826) | (n26793 & n53991) | (n53826 & n53991);
  assign n53993 = n26418 | n26793;
  assign n53994 = n53826 | n53993;
  assign n26796 = ~n53992 & n53994;
  assign n26797 = x137 & x199;
  assign n26798 = n26796 & n26797;
  assign n26799 = n26796 | n26797;
  assign n26800 = ~n26798 & n26799;
  assign n53995 = n26425 & n26800;
  assign n53996 = (n26800 & n53830) | (n26800 & n53995) | (n53830 & n53995);
  assign n53997 = n26425 | n26800;
  assign n53998 = n53830 | n53997;
  assign n26803 = ~n53996 & n53998;
  assign n26804 = x136 & x200;
  assign n26805 = n26803 & n26804;
  assign n26806 = n26803 | n26804;
  assign n26807 = ~n26805 & n26806;
  assign n53999 = n26432 & n26807;
  assign n54000 = (n26807 & n53834) | (n26807 & n53999) | (n53834 & n53999);
  assign n54001 = n26432 | n26807;
  assign n54002 = n53834 | n54001;
  assign n26810 = ~n54000 & n54002;
  assign n26811 = x135 & x201;
  assign n26812 = n26810 & n26811;
  assign n26813 = n26810 | n26811;
  assign n26814 = ~n26812 & n26813;
  assign n54003 = n26439 & n26814;
  assign n54004 = (n26814 & n53838) | (n26814 & n54003) | (n53838 & n54003);
  assign n54005 = n26439 | n26814;
  assign n54006 = n53838 | n54005;
  assign n26817 = ~n54004 & n54006;
  assign n26818 = x134 & x202;
  assign n26819 = n26817 & n26818;
  assign n26820 = n26817 | n26818;
  assign n26821 = ~n26819 & n26820;
  assign n54007 = n26446 & n26821;
  assign n54008 = (n26821 & n53842) | (n26821 & n54007) | (n53842 & n54007);
  assign n54009 = n26446 | n26821;
  assign n54010 = n53842 | n54009;
  assign n26824 = ~n54008 & n54010;
  assign n26825 = x133 & x203;
  assign n26826 = n26824 & n26825;
  assign n26827 = n26824 | n26825;
  assign n26828 = ~n26826 & n26827;
  assign n54011 = n26453 & n26828;
  assign n54012 = (n26828 & n53846) | (n26828 & n54011) | (n53846 & n54011);
  assign n54013 = n26453 | n26828;
  assign n54014 = n53846 | n54013;
  assign n26831 = ~n54012 & n54014;
  assign n26832 = x132 & x204;
  assign n26833 = n26831 & n26832;
  assign n26834 = n26831 | n26832;
  assign n26835 = ~n26833 & n26834;
  assign n54015 = n26460 & n26835;
  assign n54016 = (n26835 & n53850) | (n26835 & n54015) | (n53850 & n54015);
  assign n54017 = n26460 | n26835;
  assign n54018 = n53850 | n54017;
  assign n26838 = ~n54016 & n54018;
  assign n26839 = x131 & x205;
  assign n26840 = n26838 & n26839;
  assign n26841 = n26838 | n26839;
  assign n26842 = ~n26840 & n26841;
  assign n54019 = n26467 & n26842;
  assign n54020 = (n26842 & n53854) | (n26842 & n54019) | (n53854 & n54019);
  assign n54021 = n26467 | n26842;
  assign n54022 = n53854 | n54021;
  assign n26845 = ~n54020 & n54022;
  assign n26846 = x130 & x206;
  assign n26847 = n26845 & n26846;
  assign n26848 = n26845 | n26846;
  assign n26849 = ~n26847 & n26848;
  assign n54023 = n26474 & n26849;
  assign n54024 = (n26849 & n53859) | (n26849 & n54023) | (n53859 & n54023);
  assign n54025 = n26474 | n26849;
  assign n54026 = n53859 | n54025;
  assign n26852 = ~n54024 & n54026;
  assign n26853 = x129 & x207;
  assign n26854 = n26852 & n26853;
  assign n26855 = n26852 | n26853;
  assign n26856 = ~n26854 & n26855;
  assign n53883 = n26481 | n26483;
  assign n54027 = n26856 & n53883;
  assign n54028 = n26481 & n26856;
  assign n54029 = (n53705 & n54027) | (n53705 & n54028) | (n54027 & n54028);
  assign n54030 = n26856 | n53883;
  assign n54031 = n26481 | n26856;
  assign n54032 = (n53705 & n54030) | (n53705 & n54031) | (n54030 & n54031);
  assign n26859 = ~n54029 & n54032;
  assign n26860 = x128 & x208;
  assign n26861 = n26859 & n26860;
  assign n26862 = n26859 | n26860;
  assign n26863 = ~n26861 & n26862;
  assign n53881 = n26488 | n26490;
  assign n68948 = n26863 & n53881;
  assign n68949 = n26488 & n26863;
  assign n68950 = (n53703 & n68948) | (n53703 & n68949) | (n68948 & n68949);
  assign n68951 = n26863 | n53881;
  assign n68952 = n26488 | n26863;
  assign n68953 = (n53703 & n68951) | (n53703 & n68952) | (n68951 & n68952);
  assign n26866 = ~n68950 & n68953;
  assign n26867 = x127 & x209;
  assign n26868 = n26866 & n26867;
  assign n26869 = n26866 | n26867;
  assign n26870 = ~n26868 & n26869;
  assign n53879 = n26495 | n26497;
  assign n68954 = n26870 & n53879;
  assign n68955 = n26495 & n26870;
  assign n68956 = (n53701 & n68954) | (n53701 & n68955) | (n68954 & n68955);
  assign n68957 = n26870 | n53879;
  assign n68958 = n26495 | n26870;
  assign n68959 = (n53701 & n68957) | (n53701 & n68958) | (n68957 & n68958);
  assign n26873 = ~n68956 & n68959;
  assign n26874 = x126 & x210;
  assign n26875 = n26873 & n26874;
  assign n26876 = n26873 | n26874;
  assign n26877 = ~n26875 & n26876;
  assign n26878 = n53878 & n26877;
  assign n26879 = n53878 | n26877;
  assign n26880 = ~n26878 & n26879;
  assign n26881 = x125 & x211;
  assign n26882 = n26880 & n26881;
  assign n26883 = n26880 | n26881;
  assign n26884 = ~n26882 & n26883;
  assign n26885 = n53876 & n26884;
  assign n26886 = n53876 | n26884;
  assign n26887 = ~n26885 & n26886;
  assign n26888 = x124 & x212;
  assign n26889 = n26887 & n26888;
  assign n26890 = n26887 | n26888;
  assign n26891 = ~n26889 & n26890;
  assign n26892 = n53874 & n26891;
  assign n26893 = n53874 | n26891;
  assign n26894 = ~n26892 & n26893;
  assign n26895 = x123 & x213;
  assign n26896 = n26894 & n26895;
  assign n26897 = n26894 | n26895;
  assign n26898 = ~n26896 & n26897;
  assign n26899 = n53872 & n26898;
  assign n26900 = n53872 | n26898;
  assign n26901 = ~n26899 & n26900;
  assign n26902 = x122 & x214;
  assign n26903 = n26901 & n26902;
  assign n26904 = n26901 | n26902;
  assign n26905 = ~n26903 & n26904;
  assign n26906 = n26604 & n26905;
  assign n26907 = n26604 | n26905;
  assign n26908 = ~n26906 & n26907;
  assign n26909 = x121 & x215;
  assign n26910 = n26908 & n26909;
  assign n26911 = n26908 | n26909;
  assign n26912 = ~n26910 & n26911;
  assign n26913 = n26603 & n26912;
  assign n26914 = n26603 | n26912;
  assign n26915 = ~n26913 & n26914;
  assign n26916 = x120 & x216;
  assign n26917 = n26915 & n26916;
  assign n26918 = n26915 | n26916;
  assign n26919 = ~n26917 & n26918;
  assign n26920 = n26602 & n26919;
  assign n26921 = n26602 | n26919;
  assign n26922 = ~n26920 & n26921;
  assign n26923 = x119 & x217;
  assign n26924 = n26922 & n26923;
  assign n26925 = n26922 | n26923;
  assign n26926 = ~n26924 & n26925;
  assign n26927 = n26601 & n26926;
  assign n26928 = n26601 | n26926;
  assign n26929 = ~n26927 & n26928;
  assign n26930 = x118 & x218;
  assign n26931 = n26929 & n26930;
  assign n26932 = n26929 | n26930;
  assign n26933 = ~n26931 & n26932;
  assign n26934 = n68861 & n26933;
  assign n26935 = n68861 | n26933;
  assign n26936 = ~n26934 & n26935;
  assign n26937 = x117 & x219;
  assign n26938 = n26936 & n26937;
  assign n26939 = n26936 | n26937;
  assign n26940 = ~n26938 & n26939;
  assign n26941 = n53870 & n26940;
  assign n26942 = n53870 | n26940;
  assign n26943 = ~n26941 & n26942;
  assign n26944 = x116 & x220;
  assign n26945 = n26943 & n26944;
  assign n26946 = n26943 | n26944;
  assign n26947 = ~n26945 & n26946;
  assign n26948 = n53868 & n26947;
  assign n26949 = n53868 | n26947;
  assign n26950 = ~n26948 & n26949;
  assign n26951 = x115 & x221;
  assign n26952 = n26950 & n26951;
  assign n26953 = n26950 | n26951;
  assign n26954 = ~n26952 & n26953;
  assign n26955 = n53866 & n26954;
  assign n26956 = n53866 | n26954;
  assign n26957 = ~n26955 & n26956;
  assign n26958 = x114 & x222;
  assign n26959 = n26957 & n26958;
  assign n26960 = n26957 | n26958;
  assign n26961 = ~n26959 & n26960;
  assign n26962 = n53864 & n26961;
  assign n26963 = n53864 | n26961;
  assign n26964 = ~n26962 & n26963;
  assign n26965 = x113 & x223;
  assign n26966 = n26964 & n26965;
  assign n26967 = n26964 | n26965;
  assign n26968 = ~n26966 & n26967;
  assign n26969 = n26593 & n26968;
  assign n26970 = n26593 | n26968;
  assign n26971 = ~n26969 & n26970;
  assign n26972 = x112 & x224;
  assign n26973 = n26971 & n26972;
  assign n26974 = n26971 | n26972;
  assign n26975 = ~n26973 & n26974;
  assign n68960 = n26593 | n26965;
  assign n68961 = (n26593 & n26964) | (n26593 & n68960) | (n26964 & n68960);
  assign n54034 = (n26966 & n26968) | (n26966 & n68961) | (n26968 & n68961);
  assign n54035 = n26959 | n53864;
  assign n54036 = (n26959 & n26961) | (n26959 & n54035) | (n26961 & n54035);
  assign n54037 = n26952 | n53866;
  assign n54038 = (n26952 & n26954) | (n26952 & n54037) | (n26954 & n54037);
  assign n54039 = n26945 | n53868;
  assign n54040 = (n26945 & n26947) | (n26945 & n54039) | (n26947 & n54039);
  assign n54041 = n26938 | n53870;
  assign n54042 = (n26938 & n26940) | (n26938 & n54041) | (n26940 & n54041);
  assign n68962 = n26931 | n68861;
  assign n68963 = (n26931 & n26933) | (n26931 & n68962) | (n26933 & n68962);
  assign n26982 = n26924 | n26927;
  assign n26983 = n26917 | n26920;
  assign n26984 = n26910 | n26913;
  assign n54043 = n26903 | n26905;
  assign n54044 = (n26604 & n26903) | (n26604 & n54043) | (n26903 & n54043);
  assign n54045 = n26896 | n26898;
  assign n54046 = (n26896 & n53872) | (n26896 & n54045) | (n53872 & n54045);
  assign n54047 = n26889 | n26891;
  assign n54048 = (n26889 & n53874) | (n26889 & n54047) | (n53874 & n54047);
  assign n54049 = n26882 | n26884;
  assign n54050 = (n26882 & n53876) | (n26882 & n54049) | (n53876 & n54049);
  assign n53880 = (n26495 & n53701) | (n26495 & n53879) | (n53701 & n53879);
  assign n53882 = (n26488 & n53703) | (n26488 & n53881) | (n53703 & n53881);
  assign n53887 = (n68728 & n68863) | (n68728 & n53886) | (n68863 & n53886);
  assign n54060 = n26763 | n26765;
  assign n68964 = n26390 | n26763;
  assign n68965 = (n26763 & n26765) | (n26763 & n68964) | (n26765 & n68964);
  assign n68966 = (n53808 & n54060) | (n53808 & n68965) | (n54060 & n68965);
  assign n68967 = (n53807 & n54060) | (n53807 & n68965) | (n54060 & n68965);
  assign n68968 = (n53539 & n68966) | (n53539 & n68967) | (n68966 & n68967);
  assign n54065 = n26742 | n26744;
  assign n68969 = n26369 | n26742;
  assign n68970 = (n26742 & n26744) | (n26742 & n68969) | (n26744 & n68969);
  assign n68971 = (n53798 & n54065) | (n53798 & n68970) | (n54065 & n68970);
  assign n68972 = (n53797 & n54065) | (n53797 & n68970) | (n54065 & n68970);
  assign n68973 = (n68649 & n68971) | (n68649 & n68972) | (n68971 & n68972);
  assign n53732 = (n68569 & n68768) | (n68569 & n68770) | (n68768 & n68770);
  assign n54088 = n26665 | n68901;
  assign n68978 = n26665 | n26667;
  assign n68979 = (n26665 & n68903) | (n26665 & n68978) | (n68903 & n68978);
  assign n68980 = (n54088 & n68664) | (n54088 & n68979) | (n68664 & n68979);
  assign n68981 = (n54088 & n68663) | (n54088 & n68979) | (n68663 & n68979);
  assign n68982 = (n68409 & n68980) | (n68409 & n68981) | (n68980 & n68981);
  assign n27023 = x161 & x176;
  assign n27024 = x160 & x177;
  assign n27025 = n27023 & n27024;
  assign n27026 = n27023 | n27024;
  assign n27027 = ~n27025 & n27026;
  assign n54096 = n26644 | n26646;
  assign n54098 = n27027 & n54096;
  assign n54099 = n26644 & n27027;
  assign n68983 = (n53919 & n54098) | (n53919 & n54099) | (n54098 & n54099);
  assign n68984 = (n53918 & n54098) | (n53918 & n54099) | (n54098 & n54099);
  assign n68985 = (n68195 & n68983) | (n68195 & n68984) | (n68983 & n68984);
  assign n54101 = n27027 | n54096;
  assign n54102 = n26644 | n27027;
  assign n68986 = (n53919 & n54101) | (n53919 & n54102) | (n54101 & n54102);
  assign n68987 = (n53918 & n54101) | (n53918 & n54102) | (n54101 & n54102);
  assign n68988 = (n68195 & n68986) | (n68195 & n68987) | (n68986 & n68987);
  assign n27030 = ~n68985 & n68988;
  assign n27031 = x159 & x178;
  assign n27032 = n27030 & n27031;
  assign n27033 = n27030 | n27031;
  assign n27034 = ~n27032 & n27033;
  assign n68989 = n26278 | n26651;
  assign n68990 = (n26651 & n26653) | (n26651 & n68989) | (n26653 & n68989);
  assign n54104 = n27034 & n68990;
  assign n54094 = n26651 | n26653;
  assign n54105 = n27034 & n54094;
  assign n68991 = (n54104 & n54105) | (n54104 & n68795) | (n54105 & n68795);
  assign n68992 = (n54104 & n54105) | (n54104 & n68793) | (n54105 & n68793);
  assign n68993 = (n68389 & n68991) | (n68389 & n68992) | (n68991 & n68992);
  assign n54107 = n27034 | n68990;
  assign n54108 = n27034 | n54094;
  assign n68994 = (n54107 & n54108) | (n54107 & n68795) | (n54108 & n68795);
  assign n68995 = (n54107 & n54108) | (n54107 & n68793) | (n54108 & n68793);
  assign n68996 = (n68389 & n68994) | (n68389 & n68995) | (n68994 & n68995);
  assign n27037 = ~n68993 & n68996;
  assign n27038 = x158 & x179;
  assign n27039 = n27037 & n27038;
  assign n27040 = n27037 | n27038;
  assign n27041 = ~n27039 & n27040;
  assign n68997 = n26658 | n26660;
  assign n68998 = (n26658 & n53916) | (n26658 & n68997) | (n53916 & n68997);
  assign n54110 = n27041 & n68998;
  assign n68999 = n26285 | n26658;
  assign n69000 = (n26658 & n26660) | (n26658 & n68999) | (n26660 & n68999);
  assign n54111 = n27041 & n69000;
  assign n54112 = (n68776 & n54110) | (n68776 & n54111) | (n54110 & n54111);
  assign n54113 = n27041 | n68998;
  assign n54114 = n27041 | n69000;
  assign n54115 = (n68776 & n54113) | (n68776 & n54114) | (n54113 & n54114);
  assign n27044 = ~n54112 & n54115;
  assign n27045 = x157 & x180;
  assign n27046 = n27044 & n27045;
  assign n27047 = n27044 | n27045;
  assign n27048 = ~n27046 & n27047;
  assign n27049 = n68982 & n27048;
  assign n27050 = n68982 | n27048;
  assign n27051 = ~n27049 & n27050;
  assign n27052 = x156 & x181;
  assign n27053 = n27051 & n27052;
  assign n27054 = n27051 | n27052;
  assign n27055 = ~n27053 & n27054;
  assign n69001 = n26299 | n26672;
  assign n69002 = (n26672 & n26674) | (n26672 & n69001) | (n26674 & n69001);
  assign n54116 = n27055 & n69002;
  assign n54085 = n26672 | n26674;
  assign n54117 = n27055 & n54085;
  assign n69003 = (n53765 & n54116) | (n53765 & n54117) | (n54116 & n54117);
  assign n69004 = (n53766 & n54116) | (n53766 & n54117) | (n54116 & n54117);
  assign n69005 = (n53401 & n69003) | (n53401 & n69004) | (n69003 & n69004);
  assign n54119 = n27055 | n69002;
  assign n54120 = n27055 | n54085;
  assign n69006 = (n53765 & n54119) | (n53765 & n54120) | (n54119 & n54120);
  assign n69007 = (n53766 & n54119) | (n53766 & n54120) | (n54119 & n54120);
  assign n69008 = (n53401 & n69006) | (n53401 & n69007) | (n69006 & n69007);
  assign n27058 = ~n69005 & n69008;
  assign n27059 = x155 & x182;
  assign n27060 = n27058 & n27059;
  assign n27061 = n27058 | n27059;
  assign n27062 = ~n27060 & n27061;
  assign n69009 = n26679 | n26681;
  assign n69010 = (n26679 & n53911) | (n26679 & n69009) | (n53911 & n69009);
  assign n54122 = n27062 & n69010;
  assign n69011 = n26306 | n26679;
  assign n69012 = (n26679 & n26681) | (n26679 & n69011) | (n26681 & n69011);
  assign n54123 = n27062 & n69012;
  assign n54124 = (n53732 & n54122) | (n53732 & n54123) | (n54122 & n54123);
  assign n54125 = n27062 | n69010;
  assign n54126 = n27062 | n69012;
  assign n54127 = (n53732 & n54125) | (n53732 & n54126) | (n54125 & n54126);
  assign n27065 = ~n54124 & n54127;
  assign n27066 = x154 & x183;
  assign n27067 = n27065 & n27066;
  assign n27068 = n27065 | n27066;
  assign n27069 = ~n27067 & n27068;
  assign n54079 = n26686 | n26688;
  assign n54128 = n27069 & n54079;
  assign n54129 = n26686 & n27069;
  assign n54130 = (n68887 & n54128) | (n68887 & n54129) | (n54128 & n54129);
  assign n54131 = n27069 | n54079;
  assign n54132 = n26686 | n27069;
  assign n54133 = (n68887 & n54131) | (n68887 & n54132) | (n54131 & n54132);
  assign n27072 = ~n54130 & n54133;
  assign n27073 = x153 & x184;
  assign n27074 = n27072 & n27073;
  assign n27075 = n27072 | n27073;
  assign n27076 = ~n27074 & n27075;
  assign n54077 = n26693 | n53947;
  assign n69013 = n27076 & n54077;
  assign n68976 = n26320 | n26693;
  assign n68977 = (n26693 & n26695) | (n26693 & n68976) | (n26695 & n68976);
  assign n69014 = n27076 & n68977;
  assign n69015 = (n68766 & n69013) | (n68766 & n69014) | (n69013 & n69014);
  assign n69016 = n27076 | n54077;
  assign n69017 = n27076 | n68977;
  assign n69018 = (n68766 & n69016) | (n68766 & n69017) | (n69016 & n69017);
  assign n27079 = ~n69015 & n69018;
  assign n27080 = x152 & x185;
  assign n27081 = n27079 & n27080;
  assign n27082 = n27079 | n27080;
  assign n27083 = ~n27081 & n27082;
  assign n54074 = n26700 | n26702;
  assign n54134 = n27083 & n54074;
  assign n54135 = n26700 & n27083;
  assign n54136 = (n53905 & n54134) | (n53905 & n54135) | (n54134 & n54135);
  assign n54137 = n27083 | n54074;
  assign n54138 = n26700 | n27083;
  assign n54139 = (n53905 & n54137) | (n53905 & n54138) | (n54137 & n54138);
  assign n27086 = ~n54136 & n54139;
  assign n27087 = x151 & x186;
  assign n27088 = n27086 & n27087;
  assign n27089 = n27086 | n27087;
  assign n27090 = ~n27088 & n27089;
  assign n54072 = n26707 | n26709;
  assign n54140 = n27090 & n54072;
  assign n54141 = n26707 & n27090;
  assign n54142 = (n68878 & n54140) | (n68878 & n54141) | (n54140 & n54141);
  assign n54143 = n27090 | n54072;
  assign n54144 = n26707 | n27090;
  assign n54145 = (n68878 & n54143) | (n68878 & n54144) | (n54143 & n54144);
  assign n27093 = ~n54142 & n54145;
  assign n27094 = x150 & x187;
  assign n27095 = n27093 & n27094;
  assign n27096 = n27093 | n27094;
  assign n27097 = ~n27095 & n27096;
  assign n54146 = n26714 & n27097;
  assign n69019 = (n27097 & n53954) | (n27097 & n54146) | (n53954 & n54146);
  assign n69020 = (n27097 & n53953) | (n27097 & n54146) | (n53953 & n54146);
  assign n69021 = (n53722 & n69019) | (n53722 & n69020) | (n69019 & n69020);
  assign n54148 = n26714 | n27097;
  assign n69022 = n53954 | n54148;
  assign n69023 = n53953 | n54148;
  assign n69024 = (n53722 & n69022) | (n53722 & n69023) | (n69022 & n69023);
  assign n27100 = ~n69021 & n69024;
  assign n27101 = x149 & x188;
  assign n27102 = n27100 & n27101;
  assign n27103 = n27100 | n27101;
  assign n27104 = ~n27102 & n27103;
  assign n54070 = n26721 | n26723;
  assign n69025 = n27104 & n54070;
  assign n68974 = n26348 | n26721;
  assign n68975 = (n26721 & n26723) | (n26721 & n68974) | (n26723 & n68974);
  assign n69026 = n27104 & n68975;
  assign n69027 = (n53789 & n69025) | (n53789 & n69026) | (n69025 & n69026);
  assign n69028 = n27104 | n54070;
  assign n69029 = n27104 | n68975;
  assign n69030 = (n53789 & n69028) | (n53789 & n69029) | (n69028 & n69029);
  assign n27107 = ~n69027 & n69030;
  assign n27108 = x148 & x189;
  assign n27109 = n27107 & n27108;
  assign n27110 = n27107 | n27108;
  assign n27111 = ~n27109 & n27110;
  assign n54067 = n26728 | n26730;
  assign n54150 = n27111 & n54067;
  assign n54151 = n26728 & n27111;
  assign n54152 = (n68873 & n54150) | (n68873 & n54151) | (n54150 & n54151);
  assign n54153 = n27111 | n54067;
  assign n54154 = n26728 | n27111;
  assign n54155 = (n68873 & n54153) | (n68873 & n54154) | (n54153 & n54154);
  assign n27114 = ~n54152 & n54155;
  assign n27115 = x147 & x190;
  assign n27116 = n27114 & n27115;
  assign n27117 = n27114 | n27115;
  assign n27118 = ~n27116 & n27117;
  assign n54156 = n26735 & n27118;
  assign n69031 = (n27118 & n53964) | (n27118 & n54156) | (n53964 & n54156);
  assign n69032 = (n27118 & n53963) | (n27118 & n54156) | (n53963 & n54156);
  assign n69033 = (n68757 & n69031) | (n68757 & n69032) | (n69031 & n69032);
  assign n54158 = n26735 | n27118;
  assign n69034 = n53964 | n54158;
  assign n69035 = n53963 | n54158;
  assign n69036 = (n68757 & n69034) | (n68757 & n69035) | (n69034 & n69035);
  assign n27121 = ~n69033 & n69036;
  assign n27122 = x146 & x191;
  assign n27123 = n27121 & n27122;
  assign n27124 = n27121 | n27122;
  assign n27125 = ~n27123 & n27124;
  assign n27126 = n68973 & n27125;
  assign n27127 = n68973 | n27125;
  assign n27128 = ~n27126 & n27127;
  assign n27129 = x145 & x192;
  assign n27130 = n27128 & n27129;
  assign n27131 = n27128 | n27129;
  assign n27132 = ~n27130 & n27131;
  assign n54062 = n26749 | n26751;
  assign n54160 = n27132 & n54062;
  assign n54161 = n26749 & n27132;
  assign n54162 = (n68868 & n54160) | (n68868 & n54161) | (n54160 & n54161);
  assign n54163 = n27132 | n54062;
  assign n54164 = n26749 | n27132;
  assign n54165 = (n68868 & n54163) | (n68868 & n54164) | (n54163 & n54164);
  assign n27135 = ~n54162 & n54165;
  assign n27136 = x144 & x193;
  assign n27137 = n27135 & n27136;
  assign n27138 = n27135 | n27136;
  assign n27139 = ~n27137 & n27138;
  assign n54166 = n26756 & n27139;
  assign n69037 = (n27139 & n53974) | (n27139 & n54166) | (n53974 & n54166);
  assign n69038 = (n27139 & n53973) | (n27139 & n54166) | (n53973 & n54166);
  assign n69039 = (n68752 & n69037) | (n68752 & n69038) | (n69037 & n69038);
  assign n54168 = n26756 | n27139;
  assign n69040 = n53974 | n54168;
  assign n69041 = n53973 | n54168;
  assign n69042 = (n68752 & n69040) | (n68752 & n69041) | (n69040 & n69041);
  assign n27142 = ~n69039 & n69042;
  assign n27143 = x143 & x194;
  assign n27144 = n27142 & n27143;
  assign n27145 = n27142 | n27143;
  assign n27146 = ~n27144 & n27145;
  assign n27147 = n68968 & n27146;
  assign n27148 = n68968 | n27146;
  assign n27149 = ~n27147 & n27148;
  assign n27150 = x142 & x195;
  assign n27151 = n27149 & n27150;
  assign n27152 = n27149 | n27150;
  assign n27153 = ~n27151 & n27152;
  assign n54057 = n26770 | n26772;
  assign n54170 = n27153 & n54057;
  assign n54171 = n26770 & n27153;
  assign n54172 = (n53887 & n54170) | (n53887 & n54171) | (n54170 & n54171);
  assign n54173 = n27153 | n54057;
  assign n54174 = n26770 | n27153;
  assign n54175 = (n53887 & n54173) | (n53887 & n54174) | (n54173 & n54174);
  assign n27156 = ~n54172 & n54175;
  assign n27157 = x141 & x196;
  assign n27158 = n27156 & n27157;
  assign n27159 = n27156 | n27157;
  assign n27160 = ~n27158 & n27159;
  assign n54176 = n26777 & n27160;
  assign n54177 = (n27160 & n68944) | (n27160 & n54176) | (n68944 & n54176);
  assign n54178 = n26777 | n27160;
  assign n54179 = n68944 | n54178;
  assign n27163 = ~n54177 & n54179;
  assign n27164 = x140 & x197;
  assign n27165 = n27163 & n27164;
  assign n27166 = n27163 | n27164;
  assign n27167 = ~n27165 & n27166;
  assign n54180 = n26784 & n27167;
  assign n54181 = (n27167 & n53988) | (n27167 & n54180) | (n53988 & n54180);
  assign n54182 = n26784 | n27167;
  assign n54183 = n53988 | n54182;
  assign n27170 = ~n54181 & n54183;
  assign n27171 = x139 & x198;
  assign n27172 = n27170 & n27171;
  assign n27173 = n27170 | n27171;
  assign n27174 = ~n27172 & n27173;
  assign n54184 = n26791 & n27174;
  assign n54185 = (n27174 & n53992) | (n27174 & n54184) | (n53992 & n54184);
  assign n54186 = n26791 | n27174;
  assign n54187 = n53992 | n54186;
  assign n27177 = ~n54185 & n54187;
  assign n27178 = x138 & x199;
  assign n27179 = n27177 & n27178;
  assign n27180 = n27177 | n27178;
  assign n27181 = ~n27179 & n27180;
  assign n54188 = n26798 & n27181;
  assign n54189 = (n27181 & n53996) | (n27181 & n54188) | (n53996 & n54188);
  assign n54190 = n26798 | n27181;
  assign n54191 = n53996 | n54190;
  assign n27184 = ~n54189 & n54191;
  assign n27185 = x137 & x200;
  assign n27186 = n27184 & n27185;
  assign n27187 = n27184 | n27185;
  assign n27188 = ~n27186 & n27187;
  assign n54192 = n26805 & n27188;
  assign n54193 = (n27188 & n54000) | (n27188 & n54192) | (n54000 & n54192);
  assign n54194 = n26805 | n27188;
  assign n54195 = n54000 | n54194;
  assign n27191 = ~n54193 & n54195;
  assign n27192 = x136 & x201;
  assign n27193 = n27191 & n27192;
  assign n27194 = n27191 | n27192;
  assign n27195 = ~n27193 & n27194;
  assign n54196 = n26812 & n27195;
  assign n54197 = (n27195 & n54004) | (n27195 & n54196) | (n54004 & n54196);
  assign n54198 = n26812 | n27195;
  assign n54199 = n54004 | n54198;
  assign n27198 = ~n54197 & n54199;
  assign n27199 = x135 & x202;
  assign n27200 = n27198 & n27199;
  assign n27201 = n27198 | n27199;
  assign n27202 = ~n27200 & n27201;
  assign n54200 = n26819 & n27202;
  assign n54201 = (n27202 & n54008) | (n27202 & n54200) | (n54008 & n54200);
  assign n54202 = n26819 | n27202;
  assign n54203 = n54008 | n54202;
  assign n27205 = ~n54201 & n54203;
  assign n27206 = x134 & x203;
  assign n27207 = n27205 & n27206;
  assign n27208 = n27205 | n27206;
  assign n27209 = ~n27207 & n27208;
  assign n54204 = n26826 & n27209;
  assign n54205 = (n27209 & n54012) | (n27209 & n54204) | (n54012 & n54204);
  assign n54206 = n26826 | n27209;
  assign n54207 = n54012 | n54206;
  assign n27212 = ~n54205 & n54207;
  assign n27213 = x133 & x204;
  assign n27214 = n27212 & n27213;
  assign n27215 = n27212 | n27213;
  assign n27216 = ~n27214 & n27215;
  assign n54208 = n26833 & n27216;
  assign n54209 = (n27216 & n54016) | (n27216 & n54208) | (n54016 & n54208);
  assign n54210 = n26833 | n27216;
  assign n54211 = n54016 | n54210;
  assign n27219 = ~n54209 & n54211;
  assign n27220 = x132 & x205;
  assign n27221 = n27219 & n27220;
  assign n27222 = n27219 | n27220;
  assign n27223 = ~n27221 & n27222;
  assign n54212 = n26840 & n27223;
  assign n54213 = (n27223 & n54020) | (n27223 & n54212) | (n54020 & n54212);
  assign n54214 = n26840 | n27223;
  assign n54215 = n54020 | n54214;
  assign n27226 = ~n54213 & n54215;
  assign n27227 = x131 & x206;
  assign n27228 = n27226 & n27227;
  assign n27229 = n27226 | n27227;
  assign n27230 = ~n27228 & n27229;
  assign n54216 = n26847 & n27230;
  assign n54217 = (n27230 & n54024) | (n27230 & n54216) | (n54024 & n54216);
  assign n54218 = n26847 | n27230;
  assign n54219 = n54024 | n54218;
  assign n27233 = ~n54217 & n54219;
  assign n27234 = x130 & x207;
  assign n27235 = n27233 & n27234;
  assign n27236 = n27233 | n27234;
  assign n27237 = ~n27235 & n27236;
  assign n54220 = n26854 & n27237;
  assign n54221 = (n27237 & n54029) | (n27237 & n54220) | (n54029 & n54220);
  assign n54222 = n26854 | n27237;
  assign n54223 = n54029 | n54222;
  assign n27240 = ~n54221 & n54223;
  assign n27241 = x129 & x208;
  assign n27242 = n27240 & n27241;
  assign n27243 = n27240 | n27241;
  assign n27244 = ~n27242 & n27243;
  assign n54055 = n26861 | n26863;
  assign n54224 = n27244 & n54055;
  assign n54225 = n26861 & n27244;
  assign n54226 = (n53882 & n54224) | (n53882 & n54225) | (n54224 & n54225);
  assign n54227 = n27244 | n54055;
  assign n54228 = n26861 | n27244;
  assign n54229 = (n53882 & n54227) | (n53882 & n54228) | (n54227 & n54228);
  assign n27247 = ~n54226 & n54229;
  assign n27248 = x128 & x209;
  assign n27249 = n27247 & n27248;
  assign n27250 = n27247 | n27248;
  assign n27251 = ~n27249 & n27250;
  assign n54053 = n26868 | n26870;
  assign n69043 = n27251 & n54053;
  assign n69044 = n26868 & n27251;
  assign n69045 = (n53880 & n69043) | (n53880 & n69044) | (n69043 & n69044);
  assign n69046 = n27251 | n54053;
  assign n69047 = n26868 | n27251;
  assign n69048 = (n53880 & n69046) | (n53880 & n69047) | (n69046 & n69047);
  assign n27254 = ~n69045 & n69048;
  assign n27255 = x127 & x210;
  assign n27256 = n27254 & n27255;
  assign n27257 = n27254 | n27255;
  assign n27258 = ~n27256 & n27257;
  assign n54051 = n26875 | n26877;
  assign n69049 = n27258 & n54051;
  assign n69050 = n26875 & n27258;
  assign n69051 = (n53878 & n69049) | (n53878 & n69050) | (n69049 & n69050);
  assign n69052 = n27258 | n54051;
  assign n69053 = n26875 | n27258;
  assign n69054 = (n53878 & n69052) | (n53878 & n69053) | (n69052 & n69053);
  assign n27261 = ~n69051 & n69054;
  assign n27262 = x126 & x211;
  assign n27263 = n27261 & n27262;
  assign n27264 = n27261 | n27262;
  assign n27265 = ~n27263 & n27264;
  assign n27266 = n54050 & n27265;
  assign n27267 = n54050 | n27265;
  assign n27268 = ~n27266 & n27267;
  assign n27269 = x125 & x212;
  assign n27270 = n27268 & n27269;
  assign n27271 = n27268 | n27269;
  assign n27272 = ~n27270 & n27271;
  assign n27273 = n54048 & n27272;
  assign n27274 = n54048 | n27272;
  assign n27275 = ~n27273 & n27274;
  assign n27276 = x124 & x213;
  assign n27277 = n27275 & n27276;
  assign n27278 = n27275 | n27276;
  assign n27279 = ~n27277 & n27278;
  assign n27280 = n54046 & n27279;
  assign n27281 = n54046 | n27279;
  assign n27282 = ~n27280 & n27281;
  assign n27283 = x123 & x214;
  assign n27284 = n27282 & n27283;
  assign n27285 = n27282 | n27283;
  assign n27286 = ~n27284 & n27285;
  assign n27287 = n54044 & n27286;
  assign n27288 = n54044 | n27286;
  assign n27289 = ~n27287 & n27288;
  assign n27290 = x122 & x215;
  assign n27291 = n27289 & n27290;
  assign n27292 = n27289 | n27290;
  assign n27293 = ~n27291 & n27292;
  assign n27294 = n26984 & n27293;
  assign n27295 = n26984 | n27293;
  assign n27296 = ~n27294 & n27295;
  assign n27297 = x121 & x216;
  assign n27298 = n27296 & n27297;
  assign n27299 = n27296 | n27297;
  assign n27300 = ~n27298 & n27299;
  assign n27301 = n26983 & n27300;
  assign n27302 = n26983 | n27300;
  assign n27303 = ~n27301 & n27302;
  assign n27304 = x120 & x217;
  assign n27305 = n27303 & n27304;
  assign n27306 = n27303 | n27304;
  assign n27307 = ~n27305 & n27306;
  assign n27308 = n26982 & n27307;
  assign n27309 = n26982 | n27307;
  assign n27310 = ~n27308 & n27309;
  assign n27311 = x119 & x218;
  assign n27312 = n27310 & n27311;
  assign n27313 = n27310 | n27311;
  assign n27314 = ~n27312 & n27313;
  assign n27315 = n68963 & n27314;
  assign n27316 = n68963 | n27314;
  assign n27317 = ~n27315 & n27316;
  assign n27318 = x118 & x219;
  assign n27319 = n27317 & n27318;
  assign n27320 = n27317 | n27318;
  assign n27321 = ~n27319 & n27320;
  assign n27322 = n54042 & n27321;
  assign n27323 = n54042 | n27321;
  assign n27324 = ~n27322 & n27323;
  assign n27325 = x117 & x220;
  assign n27326 = n27324 & n27325;
  assign n27327 = n27324 | n27325;
  assign n27328 = ~n27326 & n27327;
  assign n27329 = n54040 & n27328;
  assign n27330 = n54040 | n27328;
  assign n27331 = ~n27329 & n27330;
  assign n27332 = x116 & x221;
  assign n27333 = n27331 & n27332;
  assign n27334 = n27331 | n27332;
  assign n27335 = ~n27333 & n27334;
  assign n27336 = n54038 & n27335;
  assign n27337 = n54038 | n27335;
  assign n27338 = ~n27336 & n27337;
  assign n27339 = x115 & x222;
  assign n27340 = n27338 & n27339;
  assign n27341 = n27338 | n27339;
  assign n27342 = ~n27340 & n27341;
  assign n27343 = n54036 & n27342;
  assign n27344 = n54036 | n27342;
  assign n27345 = ~n27343 & n27344;
  assign n27346 = x114 & x223;
  assign n27347 = n27345 & n27346;
  assign n27348 = n27345 | n27346;
  assign n27349 = ~n27347 & n27348;
  assign n27350 = n54034 & n27349;
  assign n27351 = n54034 | n27349;
  assign n27352 = ~n27350 & n27351;
  assign n27353 = x113 & x224;
  assign n27354 = n27352 & n27353;
  assign n27355 = n27352 | n27353;
  assign n27356 = ~n27354 & n27355;
  assign n27357 = n26973 & n27356;
  assign n27358 = n26973 | n27356;
  assign n27359 = ~n27357 & n27358;
  assign n27360 = x112 & x225;
  assign n27361 = n27359 & n27360;
  assign n27362 = n27359 | n27360;
  assign n27363 = ~n27361 & n27362;
  assign n69055 = n26973 | n27353;
  assign n69056 = (n26973 & n27352) | (n26973 & n69055) | (n27352 & n69055);
  assign n54231 = (n27354 & n27356) | (n27354 & n69056) | (n27356 & n69056);
  assign n54232 = n27347 | n54034;
  assign n54233 = (n27347 & n27349) | (n27347 & n54232) | (n27349 & n54232);
  assign n54234 = n27340 | n54036;
  assign n54235 = (n27340 & n27342) | (n27340 & n54234) | (n27342 & n54234);
  assign n54236 = n27333 | n54038;
  assign n54237 = (n27333 & n27335) | (n27333 & n54236) | (n27335 & n54236);
  assign n54238 = n27326 | n54040;
  assign n54239 = (n27326 & n27328) | (n27326 & n54238) | (n27328 & n54238);
  assign n54240 = n27319 | n54042;
  assign n54241 = (n27319 & n27321) | (n27319 & n54240) | (n27321 & n54240);
  assign n69057 = n27312 | n68963;
  assign n69058 = (n27312 & n27314) | (n27312 & n69057) | (n27314 & n69057);
  assign n27371 = n27305 | n27308;
  assign n27372 = n27298 | n27301;
  assign n54242 = n27291 | n27293;
  assign n54243 = (n26984 & n27291) | (n26984 & n54242) | (n27291 & n54242);
  assign n54244 = n27284 | n27286;
  assign n54245 = (n27284 & n54044) | (n27284 & n54244) | (n54044 & n54244);
  assign n54246 = n27277 | n27279;
  assign n54247 = (n27277 & n54046) | (n27277 & n54246) | (n54046 & n54246);
  assign n54248 = n27270 | n27272;
  assign n54249 = (n27270 & n54048) | (n27270 & n54248) | (n54048 & n54248);
  assign n54052 = (n26875 & n53878) | (n26875 & n54051) | (n53878 & n54051);
  assign n54054 = (n26868 & n53880) | (n26868 & n54053) | (n53880 & n54053);
  assign n54262 = n27137 | n27139;
  assign n69061 = n26756 | n27137;
  assign n69062 = (n27137 & n27139) | (n27137 & n69061) | (n27139 & n69061);
  assign n69063 = (n53974 & n54262) | (n53974 & n69062) | (n54262 & n69062);
  assign n69064 = (n53973 & n54262) | (n53973 & n69062) | (n54262 & n69062);
  assign n69065 = (n68752 & n69063) | (n68752 & n69064) | (n69063 & n69064);
  assign n54267 = n27116 | n27118;
  assign n69066 = n26735 | n27116;
  assign n69067 = (n27116 & n27118) | (n27116 & n69066) | (n27118 & n69066);
  assign n69068 = (n53964 & n54267) | (n53964 & n69067) | (n54267 & n69067);
  assign n69069 = (n53963 & n54267) | (n53963 & n69067) | (n54267 & n69067);
  assign n69070 = (n68757 & n69068) | (n68757 & n69069) | (n69068 & n69069);
  assign n54071 = (n53789 & n68975) | (n53789 & n54070) | (n68975 & n54070);
  assign n54272 = n27095 | n27097;
  assign n69071 = n26714 | n27095;
  assign n69072 = (n27095 & n27097) | (n27095 & n69071) | (n27097 & n69071);
  assign n69073 = (n53954 & n54272) | (n53954 & n69072) | (n54272 & n69072);
  assign n69074 = (n53953 & n54272) | (n53953 & n69072) | (n54272 & n69072);
  assign n69075 = (n53722 & n69073) | (n53722 & n69074) | (n69073 & n69074);
  assign n54282 = n27053 | n54116;
  assign n54283 = n27053 | n54117;
  assign n69082 = (n53765 & n54282) | (n53765 & n54283) | (n54282 & n54283);
  assign n69083 = (n53766 & n54282) | (n53766 & n54283) | (n54282 & n54283);
  assign n69084 = (n53401 & n69082) | (n53401 & n69083) | (n69082 & n69083);
  assign n27412 = x162 & x176;
  assign n27413 = x161 & x177;
  assign n27414 = n27412 & n27413;
  assign n27415 = n27412 | n27413;
  assign n27416 = ~n27414 & n27415;
  assign n69085 = n27025 | n27027;
  assign n69086 = (n27025 & n54096) | (n27025 & n69085) | (n54096 & n69085);
  assign n54296 = n27416 & n69086;
  assign n69087 = n26644 | n27025;
  assign n69088 = (n27025 & n27027) | (n27025 & n69087) | (n27027 & n69087);
  assign n54297 = n27416 & n69088;
  assign n69089 = (n53919 & n54296) | (n53919 & n54297) | (n54296 & n54297);
  assign n69090 = (n53918 & n54296) | (n53918 & n54297) | (n54296 & n54297);
  assign n69091 = (n68195 & n69089) | (n68195 & n69090) | (n69089 & n69090);
  assign n54299 = n27416 | n69086;
  assign n54300 = n27416 | n69088;
  assign n69092 = (n53919 & n54299) | (n53919 & n54300) | (n54299 & n54300);
  assign n69093 = (n53918 & n54299) | (n53918 & n54300) | (n54299 & n54300);
  assign n69094 = (n68195 & n69092) | (n68195 & n69093) | (n69092 & n69093);
  assign n27419 = ~n69091 & n69094;
  assign n27420 = x160 & x178;
  assign n27421 = n27419 & n27420;
  assign n27422 = n27419 | n27420;
  assign n27423 = ~n27421 & n27422;
  assign n69095 = n27032 | n27034;
  assign n69096 = (n27032 & n68990) | (n27032 & n69095) | (n68990 & n69095);
  assign n54302 = n27423 & n69096;
  assign n69097 = (n27032 & n54094) | (n27032 & n69095) | (n54094 & n69095);
  assign n54303 = n27423 & n69097;
  assign n69098 = (n54302 & n54303) | (n54302 & n68795) | (n54303 & n68795);
  assign n69099 = (n54302 & n54303) | (n54302 & n68793) | (n54303 & n68793);
  assign n69100 = (n68389 & n69098) | (n68389 & n69099) | (n69098 & n69099);
  assign n54305 = n27423 | n69096;
  assign n54306 = n27423 | n69097;
  assign n69101 = (n54305 & n54306) | (n54305 & n68795) | (n54306 & n68795);
  assign n69102 = (n54305 & n54306) | (n54305 & n68793) | (n54306 & n68793);
  assign n69103 = (n68389 & n69101) | (n68389 & n69102) | (n69101 & n69102);
  assign n27426 = ~n69100 & n69103;
  assign n27427 = x159 & x179;
  assign n27428 = n27426 & n27427;
  assign n27429 = n27426 | n27427;
  assign n27430 = ~n27428 & n27429;
  assign n69104 = n27039 | n27041;
  assign n69106 = n27430 & n69104;
  assign n69107 = n27039 & n27430;
  assign n69108 = (n68998 & n69106) | (n68998 & n69107) | (n69106 & n69107);
  assign n69109 = (n27039 & n69000) | (n27039 & n69104) | (n69000 & n69104);
  assign n54309 = n27430 & n69109;
  assign n54310 = (n68776 & n69108) | (n68776 & n54309) | (n69108 & n54309);
  assign n69110 = n27430 | n69104;
  assign n69111 = n27039 | n27430;
  assign n69112 = (n68998 & n69110) | (n68998 & n69111) | (n69110 & n69111);
  assign n54312 = n27430 | n69109;
  assign n54313 = (n68776 & n69112) | (n68776 & n54312) | (n69112 & n54312);
  assign n27433 = ~n54310 & n54313;
  assign n27434 = x158 & x180;
  assign n27435 = n27433 & n27434;
  assign n27436 = n27433 | n27434;
  assign n27437 = ~n27435 & n27436;
  assign n54285 = n27046 | n27048;
  assign n54314 = n27437 & n54285;
  assign n54315 = n27046 & n27437;
  assign n54316 = (n68982 & n54314) | (n68982 & n54315) | (n54314 & n54315);
  assign n54317 = n27437 | n54285;
  assign n54318 = n27046 | n27437;
  assign n54319 = (n68982 & n54317) | (n68982 & n54318) | (n54317 & n54318);
  assign n27440 = ~n54316 & n54319;
  assign n27441 = x157 & x181;
  assign n27442 = n27440 & n27441;
  assign n27443 = n27440 | n27441;
  assign n27444 = ~n27442 & n27443;
  assign n27445 = n69084 & n27444;
  assign n27446 = n69084 | n27444;
  assign n27447 = ~n27445 & n27446;
  assign n27448 = x156 & x182;
  assign n27449 = n27447 & n27448;
  assign n27450 = n27447 | n27448;
  assign n27451 = ~n27449 & n27450;
  assign n54320 = n27060 & n27451;
  assign n69113 = (n27451 & n54122) | (n27451 & n54320) | (n54122 & n54320);
  assign n69114 = (n27451 & n54123) | (n27451 & n54320) | (n54123 & n54320);
  assign n69115 = (n53732 & n69113) | (n53732 & n69114) | (n69113 & n69114);
  assign n54322 = n27060 | n27451;
  assign n69116 = n54122 | n54322;
  assign n69117 = n54123 | n54322;
  assign n69118 = (n53732 & n69116) | (n53732 & n69117) | (n69116 & n69117);
  assign n27454 = ~n69115 & n69118;
  assign n27455 = x155 & x183;
  assign n27456 = n27454 & n27455;
  assign n27457 = n27454 | n27455;
  assign n27458 = ~n27456 & n27457;
  assign n54279 = n27067 | n54128;
  assign n69119 = n27458 & n54279;
  assign n69080 = n26686 | n27067;
  assign n69081 = (n27067 & n27069) | (n27067 & n69080) | (n27069 & n69080);
  assign n69120 = n27458 & n69081;
  assign n69121 = (n68887 & n69119) | (n68887 & n69120) | (n69119 & n69120);
  assign n69122 = n27458 | n54279;
  assign n69123 = n27458 | n69081;
  assign n69124 = (n68887 & n69122) | (n68887 & n69123) | (n69122 & n69123);
  assign n27461 = ~n69121 & n69124;
  assign n27462 = x154 & x184;
  assign n27463 = n27461 & n27462;
  assign n27464 = n27461 | n27462;
  assign n27465 = ~n27463 & n27464;
  assign n54277 = n27074 | n27076;
  assign n54324 = n27465 & n54277;
  assign n54325 = n27074 & n27465;
  assign n69125 = (n54077 & n54324) | (n54077 & n54325) | (n54324 & n54325);
  assign n69126 = (n54324 & n54325) | (n54324 & n68977) | (n54325 & n68977);
  assign n69127 = (n68766 & n69125) | (n68766 & n69126) | (n69125 & n69126);
  assign n54327 = n27465 | n54277;
  assign n54328 = n27074 | n27465;
  assign n69128 = (n54077 & n54327) | (n54077 & n54328) | (n54327 & n54328);
  assign n69129 = (n54327 & n54328) | (n54327 & n68977) | (n54328 & n68977);
  assign n69130 = (n68766 & n69128) | (n68766 & n69129) | (n69128 & n69129);
  assign n27468 = ~n69127 & n69130;
  assign n27469 = x153 & x185;
  assign n27470 = n27468 & n27469;
  assign n27471 = n27468 | n27469;
  assign n27472 = ~n27470 & n27471;
  assign n69078 = n27081 | n27083;
  assign n69079 = (n27081 & n54074) | (n27081 & n69078) | (n54074 & n69078);
  assign n69131 = n27472 & n69079;
  assign n69076 = n26700 | n27081;
  assign n69077 = (n27081 & n27083) | (n27081 & n69076) | (n27083 & n69076);
  assign n69132 = n27472 & n69077;
  assign n69133 = (n53905 & n69131) | (n53905 & n69132) | (n69131 & n69132);
  assign n69134 = n27472 | n69079;
  assign n69135 = n27472 | n69077;
  assign n69136 = (n53905 & n69134) | (n53905 & n69135) | (n69134 & n69135);
  assign n27475 = ~n69133 & n69136;
  assign n27476 = x152 & x186;
  assign n27477 = n27475 & n27476;
  assign n27478 = n27475 | n27476;
  assign n27479 = ~n27477 & n27478;
  assign n54330 = n27088 & n27479;
  assign n54331 = (n27479 & n54142) | (n27479 & n54330) | (n54142 & n54330);
  assign n54332 = n27088 | n27479;
  assign n54333 = n54142 | n54332;
  assign n27482 = ~n54331 & n54333;
  assign n27483 = x151 & x187;
  assign n27484 = n27482 & n27483;
  assign n27485 = n27482 | n27483;
  assign n27486 = ~n27484 & n27485;
  assign n27487 = n69075 & n27486;
  assign n27488 = n69075 | n27486;
  assign n27489 = ~n27487 & n27488;
  assign n27490 = x150 & x188;
  assign n27491 = n27489 & n27490;
  assign n27492 = n27489 | n27490;
  assign n27493 = ~n27491 & n27492;
  assign n54269 = n27102 | n27104;
  assign n54334 = n27493 & n54269;
  assign n54335 = n27102 & n27493;
  assign n54336 = (n54071 & n54334) | (n54071 & n54335) | (n54334 & n54335);
  assign n54337 = n27493 | n54269;
  assign n54338 = n27102 | n27493;
  assign n54339 = (n54071 & n54337) | (n54071 & n54338) | (n54337 & n54338);
  assign n27496 = ~n54336 & n54339;
  assign n27497 = x149 & x189;
  assign n27498 = n27496 & n27497;
  assign n27499 = n27496 | n27497;
  assign n27500 = ~n27498 & n27499;
  assign n54340 = n27109 & n27500;
  assign n54341 = (n27500 & n54152) | (n27500 & n54340) | (n54152 & n54340);
  assign n54342 = n27109 | n27500;
  assign n54343 = n54152 | n54342;
  assign n27503 = ~n54341 & n54343;
  assign n27504 = x148 & x190;
  assign n27505 = n27503 & n27504;
  assign n27506 = n27503 | n27504;
  assign n27507 = ~n27505 & n27506;
  assign n27508 = n69070 & n27507;
  assign n27509 = n69070 | n27507;
  assign n27510 = ~n27508 & n27509;
  assign n27511 = x147 & x191;
  assign n27512 = n27510 & n27511;
  assign n27513 = n27510 | n27511;
  assign n27514 = ~n27512 & n27513;
  assign n54264 = n27123 | n27125;
  assign n54344 = n27514 & n54264;
  assign n54345 = n27123 & n27514;
  assign n54346 = (n68973 & n54344) | (n68973 & n54345) | (n54344 & n54345);
  assign n54347 = n27514 | n54264;
  assign n54348 = n27123 | n27514;
  assign n54349 = (n68973 & n54347) | (n68973 & n54348) | (n54347 & n54348);
  assign n27517 = ~n54346 & n54349;
  assign n27518 = x146 & x192;
  assign n27519 = n27517 & n27518;
  assign n27520 = n27517 | n27518;
  assign n27521 = ~n27519 & n27520;
  assign n54350 = n27130 & n27521;
  assign n69137 = (n27521 & n54161) | (n27521 & n54350) | (n54161 & n54350);
  assign n69138 = (n27521 & n54160) | (n27521 & n54350) | (n54160 & n54350);
  assign n69139 = (n68868 & n69137) | (n68868 & n69138) | (n69137 & n69138);
  assign n54352 = n27130 | n27521;
  assign n69140 = n54161 | n54352;
  assign n69141 = n54160 | n54352;
  assign n69142 = (n68868 & n69140) | (n68868 & n69141) | (n69140 & n69141);
  assign n27524 = ~n69139 & n69142;
  assign n27525 = x145 & x193;
  assign n27526 = n27524 & n27525;
  assign n27527 = n27524 | n27525;
  assign n27528 = ~n27526 & n27527;
  assign n27529 = n69065 & n27528;
  assign n27530 = n69065 | n27528;
  assign n27531 = ~n27529 & n27530;
  assign n27532 = x144 & x194;
  assign n27533 = n27531 & n27532;
  assign n27534 = n27531 | n27532;
  assign n27535 = ~n27533 & n27534;
  assign n54259 = n27144 | n27146;
  assign n54354 = n27535 & n54259;
  assign n54355 = n27144 & n27535;
  assign n54356 = (n68968 & n54354) | (n68968 & n54355) | (n54354 & n54355);
  assign n54357 = n27535 | n54259;
  assign n54358 = n27144 | n27535;
  assign n54359 = (n68968 & n54357) | (n68968 & n54358) | (n54357 & n54358);
  assign n27538 = ~n54356 & n54359;
  assign n27539 = x143 & x195;
  assign n27540 = n27538 & n27539;
  assign n27541 = n27538 | n27539;
  assign n27542 = ~n27540 & n27541;
  assign n54360 = n27151 & n27542;
  assign n69143 = (n27542 & n54171) | (n27542 & n54360) | (n54171 & n54360);
  assign n69144 = (n27542 & n54170) | (n27542 & n54360) | (n54170 & n54360);
  assign n69145 = (n53887 & n69143) | (n53887 & n69144) | (n69143 & n69144);
  assign n54362 = n27151 | n27542;
  assign n69146 = n54171 | n54362;
  assign n69147 = n54170 | n54362;
  assign n69148 = (n53887 & n69146) | (n53887 & n69147) | (n69146 & n69147);
  assign n27545 = ~n69145 & n69148;
  assign n27546 = x142 & x196;
  assign n27547 = n27545 & n27546;
  assign n27548 = n27545 | n27546;
  assign n27549 = ~n27547 & n27548;
  assign n54257 = n27158 | n27160;
  assign n69149 = n27549 & n54257;
  assign n69059 = n26777 | n27158;
  assign n69060 = (n27158 & n27160) | (n27158 & n69059) | (n27160 & n69059);
  assign n69150 = n27549 & n69060;
  assign n69151 = (n68944 & n69149) | (n68944 & n69150) | (n69149 & n69150);
  assign n69152 = n27549 | n54257;
  assign n69153 = n27549 | n69060;
  assign n69154 = (n68944 & n69152) | (n68944 & n69153) | (n69152 & n69153);
  assign n27552 = ~n69151 & n69154;
  assign n27553 = x141 & x197;
  assign n27554 = n27552 & n27553;
  assign n27555 = n27552 | n27553;
  assign n27556 = ~n27554 & n27555;
  assign n54364 = n27165 & n27556;
  assign n69155 = (n27556 & n54180) | (n27556 & n54364) | (n54180 & n54364);
  assign n69156 = (n27167 & n27556) | (n27167 & n54364) | (n27556 & n54364);
  assign n69157 = (n53988 & n69155) | (n53988 & n69156) | (n69155 & n69156);
  assign n54366 = n27165 | n27556;
  assign n69158 = n54180 | n54366;
  assign n69159 = n27167 | n54366;
  assign n69160 = (n53988 & n69158) | (n53988 & n69159) | (n69158 & n69159);
  assign n27559 = ~n69157 & n69160;
  assign n27560 = x140 & x198;
  assign n27561 = n27559 & n27560;
  assign n27562 = n27559 | n27560;
  assign n27563 = ~n27561 & n27562;
  assign n54368 = n27172 & n27563;
  assign n54369 = (n27563 & n54185) | (n27563 & n54368) | (n54185 & n54368);
  assign n54370 = n27172 | n27563;
  assign n54371 = n54185 | n54370;
  assign n27566 = ~n54369 & n54371;
  assign n27567 = x139 & x199;
  assign n27568 = n27566 & n27567;
  assign n27569 = n27566 | n27567;
  assign n27570 = ~n27568 & n27569;
  assign n54372 = n27179 & n27570;
  assign n54373 = (n27570 & n54189) | (n27570 & n54372) | (n54189 & n54372);
  assign n54374 = n27179 | n27570;
  assign n54375 = n54189 | n54374;
  assign n27573 = ~n54373 & n54375;
  assign n27574 = x138 & x200;
  assign n27575 = n27573 & n27574;
  assign n27576 = n27573 | n27574;
  assign n27577 = ~n27575 & n27576;
  assign n54376 = n27186 & n27577;
  assign n54377 = (n27577 & n54193) | (n27577 & n54376) | (n54193 & n54376);
  assign n54378 = n27186 | n27577;
  assign n54379 = n54193 | n54378;
  assign n27580 = ~n54377 & n54379;
  assign n27581 = x137 & x201;
  assign n27582 = n27580 & n27581;
  assign n27583 = n27580 | n27581;
  assign n27584 = ~n27582 & n27583;
  assign n54380 = n27193 & n27584;
  assign n54381 = (n27584 & n54197) | (n27584 & n54380) | (n54197 & n54380);
  assign n54382 = n27193 | n27584;
  assign n54383 = n54197 | n54382;
  assign n27587 = ~n54381 & n54383;
  assign n27588 = x136 & x202;
  assign n27589 = n27587 & n27588;
  assign n27590 = n27587 | n27588;
  assign n27591 = ~n27589 & n27590;
  assign n54384 = n27200 & n27591;
  assign n54385 = (n27591 & n54201) | (n27591 & n54384) | (n54201 & n54384);
  assign n54386 = n27200 | n27591;
  assign n54387 = n54201 | n54386;
  assign n27594 = ~n54385 & n54387;
  assign n27595 = x135 & x203;
  assign n27596 = n27594 & n27595;
  assign n27597 = n27594 | n27595;
  assign n27598 = ~n27596 & n27597;
  assign n54388 = n27207 & n27598;
  assign n54389 = (n27598 & n54205) | (n27598 & n54388) | (n54205 & n54388);
  assign n54390 = n27207 | n27598;
  assign n54391 = n54205 | n54390;
  assign n27601 = ~n54389 & n54391;
  assign n27602 = x134 & x204;
  assign n27603 = n27601 & n27602;
  assign n27604 = n27601 | n27602;
  assign n27605 = ~n27603 & n27604;
  assign n54392 = n27214 & n27605;
  assign n54393 = (n27605 & n54209) | (n27605 & n54392) | (n54209 & n54392);
  assign n54394 = n27214 | n27605;
  assign n54395 = n54209 | n54394;
  assign n27608 = ~n54393 & n54395;
  assign n27609 = x133 & x205;
  assign n27610 = n27608 & n27609;
  assign n27611 = n27608 | n27609;
  assign n27612 = ~n27610 & n27611;
  assign n54396 = n27221 & n27612;
  assign n54397 = (n27612 & n54213) | (n27612 & n54396) | (n54213 & n54396);
  assign n54398 = n27221 | n27612;
  assign n54399 = n54213 | n54398;
  assign n27615 = ~n54397 & n54399;
  assign n27616 = x132 & x206;
  assign n27617 = n27615 & n27616;
  assign n27618 = n27615 | n27616;
  assign n27619 = ~n27617 & n27618;
  assign n54400 = n27228 & n27619;
  assign n54401 = (n27619 & n54217) | (n27619 & n54400) | (n54217 & n54400);
  assign n54402 = n27228 | n27619;
  assign n54403 = n54217 | n54402;
  assign n27622 = ~n54401 & n54403;
  assign n27623 = x131 & x207;
  assign n27624 = n27622 & n27623;
  assign n27625 = n27622 | n27623;
  assign n27626 = ~n27624 & n27625;
  assign n54404 = n27235 & n27626;
  assign n54405 = (n27626 & n54221) | (n27626 & n54404) | (n54221 & n54404);
  assign n54406 = n27235 | n27626;
  assign n54407 = n54221 | n54406;
  assign n27629 = ~n54405 & n54407;
  assign n27630 = x130 & x208;
  assign n27631 = n27629 & n27630;
  assign n27632 = n27629 | n27630;
  assign n27633 = ~n27631 & n27632;
  assign n54408 = n27242 & n27633;
  assign n54409 = (n27633 & n54226) | (n27633 & n54408) | (n54226 & n54408);
  assign n54410 = n27242 | n27633;
  assign n54411 = n54226 | n54410;
  assign n27636 = ~n54409 & n54411;
  assign n27637 = x129 & x209;
  assign n27638 = n27636 & n27637;
  assign n27639 = n27636 | n27637;
  assign n27640 = ~n27638 & n27639;
  assign n54254 = n27249 | n27251;
  assign n54412 = n27640 & n54254;
  assign n54413 = n27249 & n27640;
  assign n54414 = (n54054 & n54412) | (n54054 & n54413) | (n54412 & n54413);
  assign n54415 = n27640 | n54254;
  assign n54416 = n27249 | n27640;
  assign n54417 = (n54054 & n54415) | (n54054 & n54416) | (n54415 & n54416);
  assign n27643 = ~n54414 & n54417;
  assign n27644 = x128 & x210;
  assign n27645 = n27643 & n27644;
  assign n27646 = n27643 | n27644;
  assign n27647 = ~n27645 & n27646;
  assign n54252 = n27256 | n27258;
  assign n69161 = n27647 & n54252;
  assign n69162 = n27256 & n27647;
  assign n69163 = (n54052 & n69161) | (n54052 & n69162) | (n69161 & n69162);
  assign n69164 = n27647 | n54252;
  assign n69165 = n27256 | n27647;
  assign n69166 = (n54052 & n69164) | (n54052 & n69165) | (n69164 & n69165);
  assign n27650 = ~n69163 & n69166;
  assign n27651 = x127 & x211;
  assign n27652 = n27650 & n27651;
  assign n27653 = n27650 | n27651;
  assign n27654 = ~n27652 & n27653;
  assign n54250 = n27263 | n27265;
  assign n69167 = n27654 & n54250;
  assign n69168 = n27263 & n27654;
  assign n69169 = (n54050 & n69167) | (n54050 & n69168) | (n69167 & n69168);
  assign n69170 = n27654 | n54250;
  assign n69171 = n27263 | n27654;
  assign n69172 = (n54050 & n69170) | (n54050 & n69171) | (n69170 & n69171);
  assign n27657 = ~n69169 & n69172;
  assign n27658 = x126 & x212;
  assign n27659 = n27657 & n27658;
  assign n27660 = n27657 | n27658;
  assign n27661 = ~n27659 & n27660;
  assign n27662 = n54249 & n27661;
  assign n27663 = n54249 | n27661;
  assign n27664 = ~n27662 & n27663;
  assign n27665 = x125 & x213;
  assign n27666 = n27664 & n27665;
  assign n27667 = n27664 | n27665;
  assign n27668 = ~n27666 & n27667;
  assign n27669 = n54247 & n27668;
  assign n27670 = n54247 | n27668;
  assign n27671 = ~n27669 & n27670;
  assign n27672 = x124 & x214;
  assign n27673 = n27671 & n27672;
  assign n27674 = n27671 | n27672;
  assign n27675 = ~n27673 & n27674;
  assign n27676 = n54245 & n27675;
  assign n27677 = n54245 | n27675;
  assign n27678 = ~n27676 & n27677;
  assign n27679 = x123 & x215;
  assign n27680 = n27678 & n27679;
  assign n27681 = n27678 | n27679;
  assign n27682 = ~n27680 & n27681;
  assign n27683 = n54243 & n27682;
  assign n27684 = n54243 | n27682;
  assign n27685 = ~n27683 & n27684;
  assign n27686 = x122 & x216;
  assign n27687 = n27685 & n27686;
  assign n27688 = n27685 | n27686;
  assign n27689 = ~n27687 & n27688;
  assign n27690 = n27372 & n27689;
  assign n27691 = n27372 | n27689;
  assign n27692 = ~n27690 & n27691;
  assign n27693 = x121 & x217;
  assign n27694 = n27692 & n27693;
  assign n27695 = n27692 | n27693;
  assign n27696 = ~n27694 & n27695;
  assign n27697 = n27371 & n27696;
  assign n27698 = n27371 | n27696;
  assign n27699 = ~n27697 & n27698;
  assign n27700 = x120 & x218;
  assign n27701 = n27699 & n27700;
  assign n27702 = n27699 | n27700;
  assign n27703 = ~n27701 & n27702;
  assign n27704 = n69058 & n27703;
  assign n27705 = n69058 | n27703;
  assign n27706 = ~n27704 & n27705;
  assign n27707 = x119 & x219;
  assign n27708 = n27706 & n27707;
  assign n27709 = n27706 | n27707;
  assign n27710 = ~n27708 & n27709;
  assign n27711 = n54241 & n27710;
  assign n27712 = n54241 | n27710;
  assign n27713 = ~n27711 & n27712;
  assign n27714 = x118 & x220;
  assign n27715 = n27713 & n27714;
  assign n27716 = n27713 | n27714;
  assign n27717 = ~n27715 & n27716;
  assign n27718 = n54239 & n27717;
  assign n27719 = n54239 | n27717;
  assign n27720 = ~n27718 & n27719;
  assign n27721 = x117 & x221;
  assign n27722 = n27720 & n27721;
  assign n27723 = n27720 | n27721;
  assign n27724 = ~n27722 & n27723;
  assign n27725 = n54237 & n27724;
  assign n27726 = n54237 | n27724;
  assign n27727 = ~n27725 & n27726;
  assign n27728 = x116 & x222;
  assign n27729 = n27727 & n27728;
  assign n27730 = n27727 | n27728;
  assign n27731 = ~n27729 & n27730;
  assign n27732 = n54235 & n27731;
  assign n27733 = n54235 | n27731;
  assign n27734 = ~n27732 & n27733;
  assign n27735 = x115 & x223;
  assign n27736 = n27734 & n27735;
  assign n27737 = n27734 | n27735;
  assign n27738 = ~n27736 & n27737;
  assign n27739 = n54233 & n27738;
  assign n27740 = n54233 | n27738;
  assign n27741 = ~n27739 & n27740;
  assign n27742 = x114 & x224;
  assign n27743 = n27741 & n27742;
  assign n27744 = n27741 | n27742;
  assign n27745 = ~n27743 & n27744;
  assign n27746 = n54231 & n27745;
  assign n27747 = n54231 | n27745;
  assign n27748 = ~n27746 & n27747;
  assign n27749 = x113 & x225;
  assign n27750 = n27748 & n27749;
  assign n27751 = n27748 | n27749;
  assign n27752 = ~n27750 & n27751;
  assign n27753 = n27361 & n27752;
  assign n27754 = n27361 | n27752;
  assign n27755 = ~n27753 & n27754;
  assign n27756 = x112 & x226;
  assign n27757 = n27755 & n27756;
  assign n27758 = n27755 | n27756;
  assign n27759 = ~n27757 & n27758;
  assign n69173 = n27361 | n27749;
  assign n69174 = (n27361 & n27748) | (n27361 & n69173) | (n27748 & n69173);
  assign n54419 = (n27750 & n27752) | (n27750 & n69174) | (n27752 & n69174);
  assign n54420 = n27743 | n54231;
  assign n54421 = (n27743 & n27745) | (n27743 & n54420) | (n27745 & n54420);
  assign n54422 = n27736 | n54233;
  assign n54423 = (n27736 & n27738) | (n27736 & n54422) | (n27738 & n54422);
  assign n54424 = n27729 | n54235;
  assign n54425 = (n27729 & n27731) | (n27729 & n54424) | (n27731 & n54424);
  assign n54426 = n27722 | n54237;
  assign n54427 = (n27722 & n27724) | (n27722 & n54426) | (n27724 & n54426);
  assign n54428 = n27715 | n54239;
  assign n54429 = (n27715 & n27717) | (n27715 & n54428) | (n27717 & n54428);
  assign n54430 = n27708 | n54241;
  assign n54431 = (n27708 & n27710) | (n27708 & n54430) | (n27710 & n54430);
  assign n69175 = n27701 | n69058;
  assign n69176 = (n27701 & n27703) | (n27701 & n69175) | (n27703 & n69175);
  assign n27768 = n27694 | n27697;
  assign n54432 = n27687 | n27689;
  assign n54433 = (n27372 & n27687) | (n27372 & n54432) | (n27687 & n54432);
  assign n54434 = n27680 | n27682;
  assign n54435 = (n27680 & n54243) | (n27680 & n54434) | (n54243 & n54434);
  assign n54436 = n27673 | n27675;
  assign n54437 = (n27673 & n54245) | (n27673 & n54436) | (n54245 & n54436);
  assign n54438 = n27666 | n27668;
  assign n54439 = (n27666 & n54247) | (n27666 & n54438) | (n54247 & n54438);
  assign n54251 = (n27263 & n54050) | (n27263 & n54250) | (n54050 & n54250);
  assign n54253 = (n27256 & n54052) | (n27256 & n54252) | (n54052 & n54252);
  assign n54258 = (n68944 & n69060) | (n68944 & n54257) | (n69060 & n54257);
  assign n54449 = n27540 | n27542;
  assign n69177 = n27151 | n27540;
  assign n69178 = (n27540 & n27542) | (n27540 & n69177) | (n27542 & n69177);
  assign n69179 = (n54171 & n54449) | (n54171 & n69178) | (n54449 & n69178);
  assign n69180 = (n54170 & n54449) | (n54170 & n69178) | (n54449 & n69178);
  assign n69181 = (n53887 & n69179) | (n53887 & n69180) | (n69179 & n69180);
  assign n54454 = n27519 | n27521;
  assign n69182 = n27130 | n27519;
  assign n69183 = (n27519 & n27521) | (n27519 & n69182) | (n27521 & n69182);
  assign n69184 = (n54161 & n54454) | (n54161 & n69183) | (n54454 & n69183);
  assign n69185 = (n54160 & n54454) | (n54160 & n69183) | (n54454 & n69183);
  assign n69186 = (n68868 & n69184) | (n68868 & n69185) | (n69184 & n69185);
  assign n69191 = n27074 | n27463;
  assign n69192 = (n27463 & n27465) | (n27463 & n69191) | (n27465 & n69191);
  assign n69193 = n27463 | n27465;
  assign n69194 = (n27463 & n54277) | (n27463 & n69193) | (n54277 & n69193);
  assign n69195 = (n54077 & n69192) | (n54077 & n69194) | (n69192 & n69194);
  assign n69196 = (n68977 & n69192) | (n68977 & n69194) | (n69192 & n69194);
  assign n69197 = (n68766 & n69195) | (n68766 & n69196) | (n69195 & n69196);
  assign n27809 = x163 & x176;
  assign n27810 = x162 & x177;
  assign n27811 = n27809 & n27810;
  assign n27812 = n27809 | n27810;
  assign n27813 = ~n27811 & n27812;
  assign n69198 = n27414 | n27416;
  assign n69203 = (n27414 & n69088) | (n27414 & n69198) | (n69088 & n69198);
  assign n54488 = n27813 & n69203;
  assign n69200 = n27813 & n69198;
  assign n69201 = n27414 & n27813;
  assign n69202 = (n69086 & n69200) | (n69086 & n69201) | (n69200 & n69201);
  assign n69204 = (n53919 & n54488) | (n53919 & n69202) | (n54488 & n69202);
  assign n69205 = (n53918 & n54488) | (n53918 & n69202) | (n54488 & n69202);
  assign n69206 = (n68195 & n69204) | (n68195 & n69205) | (n69204 & n69205);
  assign n54491 = n27813 | n69203;
  assign n69207 = n27813 | n69198;
  assign n69208 = n27414 | n27813;
  assign n69209 = (n69086 & n69207) | (n69086 & n69208) | (n69207 & n69208);
  assign n69210 = (n53919 & n54491) | (n53919 & n69209) | (n54491 & n69209);
  assign n69211 = (n53918 & n54491) | (n53918 & n69209) | (n54491 & n69209);
  assign n69212 = (n68195 & n69210) | (n68195 & n69211) | (n69210 & n69211);
  assign n27816 = ~n69206 & n69212;
  assign n27817 = x161 & x178;
  assign n27818 = n27816 & n27817;
  assign n27819 = n27816 | n27817;
  assign n27820 = ~n27818 & n27819;
  assign n69213 = n27421 | n27423;
  assign n69215 = n27820 & n69213;
  assign n69216 = n27421 & n27820;
  assign n69217 = (n69096 & n69215) | (n69096 & n69216) | (n69215 & n69216);
  assign n69219 = (n69097 & n69215) | (n69097 & n69216) | (n69215 & n69216);
  assign n69220 = (n68795 & n69217) | (n68795 & n69219) | (n69217 & n69219);
  assign n69221 = (n68793 & n69217) | (n68793 & n69219) | (n69217 & n69219);
  assign n69222 = (n68389 & n69220) | (n68389 & n69221) | (n69220 & n69221);
  assign n69223 = n27820 | n69213;
  assign n69224 = n27421 | n27820;
  assign n69225 = (n69096 & n69223) | (n69096 & n69224) | (n69223 & n69224);
  assign n69226 = (n69097 & n69223) | (n69097 & n69224) | (n69223 & n69224);
  assign n69227 = (n68795 & n69225) | (n68795 & n69226) | (n69225 & n69226);
  assign n69228 = (n68793 & n69225) | (n68793 & n69226) | (n69225 & n69226);
  assign n69229 = (n68389 & n69227) | (n68389 & n69228) | (n69227 & n69228);
  assign n27823 = ~n69222 & n69229;
  assign n27824 = x160 & x179;
  assign n27825 = n27823 & n27824;
  assign n27826 = n27823 | n27824;
  assign n27827 = ~n27825 & n27826;
  assign n54499 = n27428 & n27827;
  assign n69230 = (n27827 & n54309) | (n27827 & n54499) | (n54309 & n54499);
  assign n69231 = (n27827 & n54499) | (n27827 & n69108) | (n54499 & n69108);
  assign n69232 = (n68776 & n69230) | (n68776 & n69231) | (n69230 & n69231);
  assign n54501 = n27428 | n27827;
  assign n69233 = n54309 | n54501;
  assign n69234 = n54501 | n69108;
  assign n69235 = (n68776 & n69233) | (n68776 & n69234) | (n69233 & n69234);
  assign n27830 = ~n69232 & n69235;
  assign n27831 = x159 & x180;
  assign n27832 = n27830 & n27831;
  assign n27833 = n27830 | n27831;
  assign n27834 = ~n27832 & n27833;
  assign n69236 = n27435 | n27437;
  assign n69237 = (n27435 & n54285) | (n27435 & n69236) | (n54285 & n69236);
  assign n54503 = n27834 & n69237;
  assign n69238 = n27046 | n27435;
  assign n69239 = (n27435 & n27437) | (n27435 & n69238) | (n27437 & n69238);
  assign n54504 = n27834 & n69239;
  assign n54505 = (n68982 & n54503) | (n68982 & n54504) | (n54503 & n54504);
  assign n54506 = n27834 | n69237;
  assign n54507 = n27834 | n69239;
  assign n54508 = (n68982 & n54506) | (n68982 & n54507) | (n54506 & n54507);
  assign n27837 = ~n54505 & n54508;
  assign n27838 = x158 & x181;
  assign n27839 = n27837 & n27838;
  assign n27840 = n27837 | n27838;
  assign n27841 = ~n27839 & n27840;
  assign n54476 = n27442 | n27444;
  assign n54509 = n27841 & n54476;
  assign n54510 = n27442 & n27841;
  assign n54511 = (n69084 & n54509) | (n69084 & n54510) | (n54509 & n54510);
  assign n54512 = n27841 | n54476;
  assign n54513 = n27442 | n27841;
  assign n54514 = (n69084 & n54512) | (n69084 & n54513) | (n54512 & n54513);
  assign n27844 = ~n54511 & n54514;
  assign n27845 = x157 & x182;
  assign n27846 = n27844 & n27845;
  assign n27847 = n27844 | n27845;
  assign n27848 = ~n27846 & n27847;
  assign n69240 = n27060 | n27449;
  assign n69241 = (n27449 & n27451) | (n27449 & n69240) | (n27451 & n69240);
  assign n54515 = n27848 & n69241;
  assign n54474 = n27449 | n27451;
  assign n54516 = n27848 & n54474;
  assign n69242 = (n54122 & n54515) | (n54122 & n54516) | (n54515 & n54516);
  assign n69243 = (n54123 & n54515) | (n54123 & n54516) | (n54515 & n54516);
  assign n69244 = (n53732 & n69242) | (n53732 & n69243) | (n69242 & n69243);
  assign n54518 = n27848 | n69241;
  assign n54519 = n27848 | n54474;
  assign n69245 = (n54122 & n54518) | (n54122 & n54519) | (n54518 & n54519);
  assign n69246 = (n54123 & n54518) | (n54123 & n54519) | (n54518 & n54519);
  assign n69247 = (n53732 & n69245) | (n53732 & n69246) | (n69245 & n69246);
  assign n27851 = ~n69244 & n69247;
  assign n27852 = x156 & x183;
  assign n27853 = n27851 & n27852;
  assign n27854 = n27851 | n27852;
  assign n27855 = ~n27853 & n27854;
  assign n54471 = n27456 | n27458;
  assign n54521 = n27855 & n54471;
  assign n54522 = n27456 & n27855;
  assign n69248 = (n54279 & n54521) | (n54279 & n54522) | (n54521 & n54522);
  assign n69249 = (n54521 & n54522) | (n54521 & n69081) | (n54522 & n69081);
  assign n69250 = (n68887 & n69248) | (n68887 & n69249) | (n69248 & n69249);
  assign n54524 = n27855 | n54471;
  assign n54525 = n27456 | n27855;
  assign n69251 = (n54279 & n54524) | (n54279 & n54525) | (n54524 & n54525);
  assign n69252 = (n54524 & n54525) | (n54524 & n69081) | (n54525 & n69081);
  assign n69253 = (n68887 & n69251) | (n68887 & n69252) | (n69251 & n69252);
  assign n27858 = ~n69250 & n69253;
  assign n27859 = x155 & x184;
  assign n27860 = n27858 & n27859;
  assign n27861 = n27858 | n27859;
  assign n27862 = ~n27860 & n27861;
  assign n27863 = n69197 & n27862;
  assign n27864 = n69197 | n27862;
  assign n27865 = ~n27863 & n27864;
  assign n27866 = x154 & x185;
  assign n27867 = n27865 & n27866;
  assign n27868 = n27865 | n27866;
  assign n27869 = ~n27867 & n27868;
  assign n54466 = n27470 | n27472;
  assign n54527 = n27869 & n54466;
  assign n54528 = n27470 & n27869;
  assign n69254 = (n54527 & n54528) | (n54527 & n69079) | (n54528 & n69079);
  assign n69255 = (n54527 & n54528) | (n54527 & n69077) | (n54528 & n69077);
  assign n69256 = (n53905 & n69254) | (n53905 & n69255) | (n69254 & n69255);
  assign n54530 = n27869 | n54466;
  assign n54531 = n27470 | n27869;
  assign n69257 = (n54530 & n54531) | (n54530 & n69079) | (n54531 & n69079);
  assign n69258 = (n54530 & n54531) | (n54530 & n69077) | (n54531 & n69077);
  assign n69259 = (n53905 & n69257) | (n53905 & n69258) | (n69257 & n69258);
  assign n27872 = ~n69256 & n69259;
  assign n27873 = x153 & x186;
  assign n27874 = n27872 & n27873;
  assign n27875 = n27872 | n27873;
  assign n27876 = ~n27874 & n27875;
  assign n54464 = n27477 | n27479;
  assign n69260 = n27876 & n54464;
  assign n69189 = n27088 | n27477;
  assign n69190 = (n27477 & n27479) | (n27477 & n69189) | (n27479 & n69189);
  assign n69261 = n27876 & n69190;
  assign n69262 = (n54142 & n69260) | (n54142 & n69261) | (n69260 & n69261);
  assign n69263 = n27876 | n54464;
  assign n69264 = n27876 | n69190;
  assign n69265 = (n54142 & n69263) | (n54142 & n69264) | (n69263 & n69264);
  assign n27879 = ~n69262 & n69265;
  assign n27880 = x152 & x187;
  assign n27881 = n27879 & n27880;
  assign n27882 = n27879 | n27880;
  assign n27883 = ~n27881 & n27882;
  assign n54461 = n27484 | n27486;
  assign n54533 = n27883 & n54461;
  assign n54534 = n27484 & n27883;
  assign n54535 = (n69075 & n54533) | (n69075 & n54534) | (n54533 & n54534);
  assign n54536 = n27883 | n54461;
  assign n54537 = n27484 | n27883;
  assign n54538 = (n69075 & n54536) | (n69075 & n54537) | (n54536 & n54537);
  assign n27886 = ~n54535 & n54538;
  assign n27887 = x151 & x188;
  assign n27888 = n27886 & n27887;
  assign n27889 = n27886 | n27887;
  assign n27890 = ~n27888 & n27889;
  assign n54539 = n27491 & n27890;
  assign n69266 = (n27890 & n54335) | (n27890 & n54539) | (n54335 & n54539);
  assign n69267 = (n27890 & n54334) | (n27890 & n54539) | (n54334 & n54539);
  assign n69268 = (n54071 & n69266) | (n54071 & n69267) | (n69266 & n69267);
  assign n54541 = n27491 | n27890;
  assign n69269 = n54335 | n54541;
  assign n69270 = n54334 | n54541;
  assign n69271 = (n54071 & n69269) | (n54071 & n69270) | (n69269 & n69270);
  assign n27893 = ~n69268 & n69271;
  assign n27894 = x150 & x189;
  assign n27895 = n27893 & n27894;
  assign n27896 = n27893 | n27894;
  assign n27897 = ~n27895 & n27896;
  assign n54459 = n27498 | n27500;
  assign n69272 = n27897 & n54459;
  assign n69187 = n27109 | n27498;
  assign n69188 = (n27498 & n27500) | (n27498 & n69187) | (n27500 & n69187);
  assign n69273 = n27897 & n69188;
  assign n69274 = (n54152 & n69272) | (n54152 & n69273) | (n69272 & n69273);
  assign n69275 = n27897 | n54459;
  assign n69276 = n27897 | n69188;
  assign n69277 = (n54152 & n69275) | (n54152 & n69276) | (n69275 & n69276);
  assign n27900 = ~n69274 & n69277;
  assign n27901 = x149 & x190;
  assign n27902 = n27900 & n27901;
  assign n27903 = n27900 | n27901;
  assign n27904 = ~n27902 & n27903;
  assign n54456 = n27505 | n27507;
  assign n54543 = n27904 & n54456;
  assign n54544 = n27505 & n27904;
  assign n54545 = (n69070 & n54543) | (n69070 & n54544) | (n54543 & n54544);
  assign n54546 = n27904 | n54456;
  assign n54547 = n27505 | n27904;
  assign n54548 = (n69070 & n54546) | (n69070 & n54547) | (n54546 & n54547);
  assign n27907 = ~n54545 & n54548;
  assign n27908 = x148 & x191;
  assign n27909 = n27907 & n27908;
  assign n27910 = n27907 | n27908;
  assign n27911 = ~n27909 & n27910;
  assign n54549 = n27512 & n27911;
  assign n69278 = (n27911 & n54345) | (n27911 & n54549) | (n54345 & n54549);
  assign n69279 = (n27911 & n54344) | (n27911 & n54549) | (n54344 & n54549);
  assign n69280 = (n68973 & n69278) | (n68973 & n69279) | (n69278 & n69279);
  assign n54551 = n27512 | n27911;
  assign n69281 = n54345 | n54551;
  assign n69282 = n54344 | n54551;
  assign n69283 = (n68973 & n69281) | (n68973 & n69282) | (n69281 & n69282);
  assign n27914 = ~n69280 & n69283;
  assign n27915 = x147 & x192;
  assign n27916 = n27914 & n27915;
  assign n27917 = n27914 | n27915;
  assign n27918 = ~n27916 & n27917;
  assign n27919 = n69186 & n27918;
  assign n27920 = n69186 | n27918;
  assign n27921 = ~n27919 & n27920;
  assign n27922 = x146 & x193;
  assign n27923 = n27921 & n27922;
  assign n27924 = n27921 | n27922;
  assign n27925 = ~n27923 & n27924;
  assign n54451 = n27526 | n27528;
  assign n54553 = n27925 & n54451;
  assign n54554 = n27526 & n27925;
  assign n54555 = (n69065 & n54553) | (n69065 & n54554) | (n54553 & n54554);
  assign n54556 = n27925 | n54451;
  assign n54557 = n27526 | n27925;
  assign n54558 = (n69065 & n54556) | (n69065 & n54557) | (n54556 & n54557);
  assign n27928 = ~n54555 & n54558;
  assign n27929 = x145 & x194;
  assign n27930 = n27928 & n27929;
  assign n27931 = n27928 | n27929;
  assign n27932 = ~n27930 & n27931;
  assign n54559 = n27533 & n27932;
  assign n69284 = (n27932 & n54355) | (n27932 & n54559) | (n54355 & n54559);
  assign n69285 = (n27932 & n54354) | (n27932 & n54559) | (n54354 & n54559);
  assign n69286 = (n68968 & n69284) | (n68968 & n69285) | (n69284 & n69285);
  assign n54561 = n27533 | n27932;
  assign n69287 = n54355 | n54561;
  assign n69288 = n54354 | n54561;
  assign n69289 = (n68968 & n69287) | (n68968 & n69288) | (n69287 & n69288);
  assign n27935 = ~n69286 & n69289;
  assign n27936 = x144 & x195;
  assign n27937 = n27935 & n27936;
  assign n27938 = n27935 | n27936;
  assign n27939 = ~n27937 & n27938;
  assign n27940 = n69181 & n27939;
  assign n27941 = n69181 | n27939;
  assign n27942 = ~n27940 & n27941;
  assign n27943 = x143 & x196;
  assign n27944 = n27942 & n27943;
  assign n27945 = n27942 | n27943;
  assign n27946 = ~n27944 & n27945;
  assign n54446 = n27547 | n27549;
  assign n54563 = n27946 & n54446;
  assign n54564 = n27547 & n27946;
  assign n54565 = (n54258 & n54563) | (n54258 & n54564) | (n54563 & n54564);
  assign n54566 = n27946 | n54446;
  assign n54567 = n27547 | n27946;
  assign n54568 = (n54258 & n54566) | (n54258 & n54567) | (n54566 & n54567);
  assign n27949 = ~n54565 & n54568;
  assign n27950 = x142 & x197;
  assign n27951 = n27949 & n27950;
  assign n27952 = n27949 | n27950;
  assign n27953 = ~n27951 & n27952;
  assign n54569 = n27554 & n27953;
  assign n54570 = (n27953 & n69157) | (n27953 & n54569) | (n69157 & n54569);
  assign n54571 = n27554 | n27953;
  assign n54572 = n69157 | n54571;
  assign n27956 = ~n54570 & n54572;
  assign n27957 = x141 & x198;
  assign n27958 = n27956 & n27957;
  assign n27959 = n27956 | n27957;
  assign n27960 = ~n27958 & n27959;
  assign n54573 = n27561 & n27960;
  assign n54574 = (n27960 & n54369) | (n27960 & n54573) | (n54369 & n54573);
  assign n54575 = n27561 | n27960;
  assign n54576 = n54369 | n54575;
  assign n27963 = ~n54574 & n54576;
  assign n27964 = x140 & x199;
  assign n27965 = n27963 & n27964;
  assign n27966 = n27963 | n27964;
  assign n27967 = ~n27965 & n27966;
  assign n54577 = n27568 & n27967;
  assign n54578 = (n27967 & n54373) | (n27967 & n54577) | (n54373 & n54577);
  assign n54579 = n27568 | n27967;
  assign n54580 = n54373 | n54579;
  assign n27970 = ~n54578 & n54580;
  assign n27971 = x139 & x200;
  assign n27972 = n27970 & n27971;
  assign n27973 = n27970 | n27971;
  assign n27974 = ~n27972 & n27973;
  assign n54581 = n27575 & n27974;
  assign n54582 = (n27974 & n54377) | (n27974 & n54581) | (n54377 & n54581);
  assign n54583 = n27575 | n27974;
  assign n54584 = n54377 | n54583;
  assign n27977 = ~n54582 & n54584;
  assign n27978 = x138 & x201;
  assign n27979 = n27977 & n27978;
  assign n27980 = n27977 | n27978;
  assign n27981 = ~n27979 & n27980;
  assign n54585 = n27582 & n27981;
  assign n54586 = (n27981 & n54381) | (n27981 & n54585) | (n54381 & n54585);
  assign n54587 = n27582 | n27981;
  assign n54588 = n54381 | n54587;
  assign n27984 = ~n54586 & n54588;
  assign n27985 = x137 & x202;
  assign n27986 = n27984 & n27985;
  assign n27987 = n27984 | n27985;
  assign n27988 = ~n27986 & n27987;
  assign n54589 = n27589 & n27988;
  assign n54590 = (n27988 & n54385) | (n27988 & n54589) | (n54385 & n54589);
  assign n54591 = n27589 | n27988;
  assign n54592 = n54385 | n54591;
  assign n27991 = ~n54590 & n54592;
  assign n27992 = x136 & x203;
  assign n27993 = n27991 & n27992;
  assign n27994 = n27991 | n27992;
  assign n27995 = ~n27993 & n27994;
  assign n54593 = n27596 & n27995;
  assign n54594 = (n27995 & n54389) | (n27995 & n54593) | (n54389 & n54593);
  assign n54595 = n27596 | n27995;
  assign n54596 = n54389 | n54595;
  assign n27998 = ~n54594 & n54596;
  assign n27999 = x135 & x204;
  assign n28000 = n27998 & n27999;
  assign n28001 = n27998 | n27999;
  assign n28002 = ~n28000 & n28001;
  assign n54597 = n27603 & n28002;
  assign n54598 = (n28002 & n54393) | (n28002 & n54597) | (n54393 & n54597);
  assign n54599 = n27603 | n28002;
  assign n54600 = n54393 | n54599;
  assign n28005 = ~n54598 & n54600;
  assign n28006 = x134 & x205;
  assign n28007 = n28005 & n28006;
  assign n28008 = n28005 | n28006;
  assign n28009 = ~n28007 & n28008;
  assign n54601 = n27610 & n28009;
  assign n54602 = (n28009 & n54397) | (n28009 & n54601) | (n54397 & n54601);
  assign n54603 = n27610 | n28009;
  assign n54604 = n54397 | n54603;
  assign n28012 = ~n54602 & n54604;
  assign n28013 = x133 & x206;
  assign n28014 = n28012 & n28013;
  assign n28015 = n28012 | n28013;
  assign n28016 = ~n28014 & n28015;
  assign n54605 = n27617 & n28016;
  assign n54606 = (n28016 & n54401) | (n28016 & n54605) | (n54401 & n54605);
  assign n54607 = n27617 | n28016;
  assign n54608 = n54401 | n54607;
  assign n28019 = ~n54606 & n54608;
  assign n28020 = x132 & x207;
  assign n28021 = n28019 & n28020;
  assign n28022 = n28019 | n28020;
  assign n28023 = ~n28021 & n28022;
  assign n54609 = n27624 & n28023;
  assign n54610 = (n28023 & n54405) | (n28023 & n54609) | (n54405 & n54609);
  assign n54611 = n27624 | n28023;
  assign n54612 = n54405 | n54611;
  assign n28026 = ~n54610 & n54612;
  assign n28027 = x131 & x208;
  assign n28028 = n28026 & n28027;
  assign n28029 = n28026 | n28027;
  assign n28030 = ~n28028 & n28029;
  assign n54613 = n27631 & n28030;
  assign n54614 = (n28030 & n54409) | (n28030 & n54613) | (n54409 & n54613);
  assign n54615 = n27631 | n28030;
  assign n54616 = n54409 | n54615;
  assign n28033 = ~n54614 & n54616;
  assign n28034 = x130 & x209;
  assign n28035 = n28033 & n28034;
  assign n28036 = n28033 | n28034;
  assign n28037 = ~n28035 & n28036;
  assign n54617 = n27638 & n28037;
  assign n54618 = (n28037 & n54414) | (n28037 & n54617) | (n54414 & n54617);
  assign n54619 = n27638 | n28037;
  assign n54620 = n54414 | n54619;
  assign n28040 = ~n54618 & n54620;
  assign n28041 = x129 & x210;
  assign n28042 = n28040 & n28041;
  assign n28043 = n28040 | n28041;
  assign n28044 = ~n28042 & n28043;
  assign n54444 = n27645 | n27647;
  assign n54621 = n28044 & n54444;
  assign n54622 = n27645 & n28044;
  assign n54623 = (n54253 & n54621) | (n54253 & n54622) | (n54621 & n54622);
  assign n54624 = n28044 | n54444;
  assign n54625 = n27645 | n28044;
  assign n54626 = (n54253 & n54624) | (n54253 & n54625) | (n54624 & n54625);
  assign n28047 = ~n54623 & n54626;
  assign n28048 = x128 & x211;
  assign n28049 = n28047 & n28048;
  assign n28050 = n28047 | n28048;
  assign n28051 = ~n28049 & n28050;
  assign n54442 = n27652 | n27654;
  assign n69290 = n28051 & n54442;
  assign n69291 = n27652 & n28051;
  assign n69292 = (n54251 & n69290) | (n54251 & n69291) | (n69290 & n69291);
  assign n69293 = n28051 | n54442;
  assign n69294 = n27652 | n28051;
  assign n69295 = (n54251 & n69293) | (n54251 & n69294) | (n69293 & n69294);
  assign n28054 = ~n69292 & n69295;
  assign n28055 = x127 & x212;
  assign n28056 = n28054 & n28055;
  assign n28057 = n28054 | n28055;
  assign n28058 = ~n28056 & n28057;
  assign n54440 = n27659 | n27661;
  assign n69296 = n28058 & n54440;
  assign n69297 = n27659 & n28058;
  assign n69298 = (n54249 & n69296) | (n54249 & n69297) | (n69296 & n69297);
  assign n69299 = n28058 | n54440;
  assign n69300 = n27659 | n28058;
  assign n69301 = (n54249 & n69299) | (n54249 & n69300) | (n69299 & n69300);
  assign n28061 = ~n69298 & n69301;
  assign n28062 = x126 & x213;
  assign n28063 = n28061 & n28062;
  assign n28064 = n28061 | n28062;
  assign n28065 = ~n28063 & n28064;
  assign n28066 = n54439 & n28065;
  assign n28067 = n54439 | n28065;
  assign n28068 = ~n28066 & n28067;
  assign n28069 = x125 & x214;
  assign n28070 = n28068 & n28069;
  assign n28071 = n28068 | n28069;
  assign n28072 = ~n28070 & n28071;
  assign n28073 = n54437 & n28072;
  assign n28074 = n54437 | n28072;
  assign n28075 = ~n28073 & n28074;
  assign n28076 = x124 & x215;
  assign n28077 = n28075 & n28076;
  assign n28078 = n28075 | n28076;
  assign n28079 = ~n28077 & n28078;
  assign n28080 = n54435 & n28079;
  assign n28081 = n54435 | n28079;
  assign n28082 = ~n28080 & n28081;
  assign n28083 = x123 & x216;
  assign n28084 = n28082 & n28083;
  assign n28085 = n28082 | n28083;
  assign n28086 = ~n28084 & n28085;
  assign n28087 = n54433 & n28086;
  assign n28088 = n54433 | n28086;
  assign n28089 = ~n28087 & n28088;
  assign n28090 = x122 & x217;
  assign n28091 = n28089 & n28090;
  assign n28092 = n28089 | n28090;
  assign n28093 = ~n28091 & n28092;
  assign n28094 = n27768 & n28093;
  assign n28095 = n27768 | n28093;
  assign n28096 = ~n28094 & n28095;
  assign n28097 = x121 & x218;
  assign n28098 = n28096 & n28097;
  assign n28099 = n28096 | n28097;
  assign n28100 = ~n28098 & n28099;
  assign n28101 = n69176 & n28100;
  assign n28102 = n69176 | n28100;
  assign n28103 = ~n28101 & n28102;
  assign n28104 = x120 & x219;
  assign n28105 = n28103 & n28104;
  assign n28106 = n28103 | n28104;
  assign n28107 = ~n28105 & n28106;
  assign n28108 = n54431 & n28107;
  assign n28109 = n54431 | n28107;
  assign n28110 = ~n28108 & n28109;
  assign n28111 = x119 & x220;
  assign n28112 = n28110 & n28111;
  assign n28113 = n28110 | n28111;
  assign n28114 = ~n28112 & n28113;
  assign n28115 = n54429 & n28114;
  assign n28116 = n54429 | n28114;
  assign n28117 = ~n28115 & n28116;
  assign n28118 = x118 & x221;
  assign n28119 = n28117 & n28118;
  assign n28120 = n28117 | n28118;
  assign n28121 = ~n28119 & n28120;
  assign n28122 = n54427 & n28121;
  assign n28123 = n54427 | n28121;
  assign n28124 = ~n28122 & n28123;
  assign n28125 = x117 & x222;
  assign n28126 = n28124 & n28125;
  assign n28127 = n28124 | n28125;
  assign n28128 = ~n28126 & n28127;
  assign n28129 = n54425 & n28128;
  assign n28130 = n54425 | n28128;
  assign n28131 = ~n28129 & n28130;
  assign n28132 = x116 & x223;
  assign n28133 = n28131 & n28132;
  assign n28134 = n28131 | n28132;
  assign n28135 = ~n28133 & n28134;
  assign n28136 = n54423 & n28135;
  assign n28137 = n54423 | n28135;
  assign n28138 = ~n28136 & n28137;
  assign n28139 = x115 & x224;
  assign n28140 = n28138 & n28139;
  assign n28141 = n28138 | n28139;
  assign n28142 = ~n28140 & n28141;
  assign n28143 = n54421 & n28142;
  assign n28144 = n54421 | n28142;
  assign n28145 = ~n28143 & n28144;
  assign n28146 = x114 & x225;
  assign n28147 = n28145 & n28146;
  assign n28148 = n28145 | n28146;
  assign n28149 = ~n28147 & n28148;
  assign n28150 = n54419 & n28149;
  assign n28151 = n54419 | n28149;
  assign n28152 = ~n28150 & n28151;
  assign n28153 = x113 & x226;
  assign n28154 = n28152 & n28153;
  assign n28155 = n28152 | n28153;
  assign n28156 = ~n28154 & n28155;
  assign n28157 = n27757 & n28156;
  assign n28158 = n27757 | n28156;
  assign n28159 = ~n28157 & n28158;
  assign n28160 = x112 & x227;
  assign n28161 = n28159 & n28160;
  assign n28162 = n28159 | n28160;
  assign n28163 = ~n28161 & n28162;
  assign n69302 = n27757 | n28153;
  assign n69303 = (n27757 & n28152) | (n27757 & n69302) | (n28152 & n69302);
  assign n54628 = (n28154 & n28156) | (n28154 & n69303) | (n28156 & n69303);
  assign n54629 = n28147 | n54419;
  assign n54630 = (n28147 & n28149) | (n28147 & n54629) | (n28149 & n54629);
  assign n54631 = n28140 | n54421;
  assign n54632 = (n28140 & n28142) | (n28140 & n54631) | (n28142 & n54631);
  assign n54633 = n28133 | n54423;
  assign n54634 = (n28133 & n28135) | (n28133 & n54633) | (n28135 & n54633);
  assign n54635 = n28126 | n54425;
  assign n54636 = (n28126 & n28128) | (n28126 & n54635) | (n28128 & n54635);
  assign n54637 = n28119 | n54427;
  assign n54638 = (n28119 & n28121) | (n28119 & n54637) | (n28121 & n54637);
  assign n54639 = n28112 | n54429;
  assign n54640 = (n28112 & n28114) | (n28112 & n54639) | (n28114 & n54639);
  assign n54641 = n28105 | n54431;
  assign n54642 = (n28105 & n28107) | (n28105 & n54641) | (n28107 & n54641);
  assign n69304 = n28098 | n69176;
  assign n69305 = (n28098 & n28100) | (n28098 & n69304) | (n28100 & n69304);
  assign n54643 = n28091 | n28093;
  assign n54644 = (n27768 & n28091) | (n27768 & n54643) | (n28091 & n54643);
  assign n54645 = n28084 | n28086;
  assign n54646 = (n28084 & n54433) | (n28084 & n54645) | (n54433 & n54645);
  assign n54647 = n28077 | n28079;
  assign n54648 = (n28077 & n54435) | (n28077 & n54647) | (n54435 & n54647);
  assign n54649 = n28070 | n28072;
  assign n54650 = (n28070 & n54437) | (n28070 & n54649) | (n54437 & n54649);
  assign n54441 = (n27659 & n54249) | (n27659 & n54440) | (n54249 & n54440);
  assign n54443 = (n27652 & n54251) | (n27652 & n54442) | (n54251 & n54442);
  assign n54663 = n27930 | n27932;
  assign n69308 = n27533 | n27930;
  assign n69309 = (n27930 & n27932) | (n27930 & n69308) | (n27932 & n69308);
  assign n69310 = (n54355 & n54663) | (n54355 & n69309) | (n54663 & n69309);
  assign n69311 = (n54354 & n54663) | (n54354 & n69309) | (n54663 & n69309);
  assign n69312 = (n68968 & n69310) | (n68968 & n69311) | (n69310 & n69311);
  assign n54668 = n27909 | n27911;
  assign n69313 = n27512 | n27909;
  assign n69314 = (n27909 & n27911) | (n27909 & n69313) | (n27911 & n69313);
  assign n69315 = (n54345 & n54668) | (n54345 & n69314) | (n54668 & n69314);
  assign n69316 = (n54344 & n54668) | (n54344 & n69314) | (n54668 & n69314);
  assign n69317 = (n68973 & n69315) | (n68973 & n69316) | (n69315 & n69316);
  assign n54460 = (n54152 & n69188) | (n54152 & n54459) | (n69188 & n54459);
  assign n54673 = n27888 | n27890;
  assign n69318 = n27491 | n27888;
  assign n69319 = (n27888 & n27890) | (n27888 & n69318) | (n27890 & n69318);
  assign n69320 = (n54335 & n54673) | (n54335 & n69319) | (n54673 & n69319);
  assign n69321 = (n54334 & n54673) | (n54334 & n69319) | (n54673 & n69319);
  assign n69322 = (n54071 & n69320) | (n54071 & n69321) | (n69320 & n69321);
  assign n54276 = (n53905 & n69077) | (n53905 & n69079) | (n69077 & n69079);
  assign n69325 = n27853 | n27855;
  assign n69326 = (n27853 & n54471) | (n27853 & n69325) | (n54471 & n69325);
  assign n69327 = n27456 | n27853;
  assign n69328 = (n27853 & n27855) | (n27853 & n69327) | (n27855 & n69327);
  assign n69329 = (n54279 & n69326) | (n54279 & n69328) | (n69326 & n69328);
  assign n69330 = (n69081 & n69326) | (n69081 & n69328) | (n69326 & n69328);
  assign n69331 = (n68887 & n69329) | (n68887 & n69330) | (n69329 & n69330);
  assign n28214 = x164 & x176;
  assign n28215 = x163 & x177;
  assign n28216 = n28214 & n28215;
  assign n28217 = n28214 | n28215;
  assign n28218 = ~n28216 & n28217;
  assign n69335 = n27811 & n28218;
  assign n69336 = (n28218 & n69202) | (n28218 & n69335) | (n69202 & n69335);
  assign n69337 = n27811 | n27813;
  assign n69339 = n28218 & n69337;
  assign n69340 = (n69203 & n69335) | (n69203 & n69339) | (n69335 & n69339);
  assign n69341 = (n53919 & n69336) | (n53919 & n69340) | (n69336 & n69340);
  assign n69342 = (n53918 & n69336) | (n53918 & n69340) | (n69336 & n69340);
  assign n69343 = (n68195 & n69341) | (n68195 & n69342) | (n69341 & n69342);
  assign n69344 = n27811 | n28218;
  assign n69345 = n69202 | n69344;
  assign n69346 = n28218 | n69337;
  assign n69347 = (n69203 & n69344) | (n69203 & n69346) | (n69344 & n69346);
  assign n69348 = (n53919 & n69345) | (n53919 & n69347) | (n69345 & n69347);
  assign n69349 = (n53918 & n69345) | (n53918 & n69347) | (n69345 & n69347);
  assign n69350 = (n68195 & n69348) | (n68195 & n69349) | (n69348 & n69349);
  assign n28221 = ~n69343 & n69350;
  assign n28222 = x162 & x178;
  assign n28223 = n28221 & n28222;
  assign n28224 = n28221 | n28222;
  assign n28225 = ~n28223 & n28224;
  assign n54703 = n27818 & n28225;
  assign n69351 = (n28225 & n54703) | (n28225 & n69221) | (n54703 & n69221);
  assign n69352 = (n28225 & n54703) | (n28225 & n69220) | (n54703 & n69220);
  assign n69353 = (n68389 & n69351) | (n68389 & n69352) | (n69351 & n69352);
  assign n54705 = n27818 | n28225;
  assign n69354 = n54705 | n69221;
  assign n69355 = n54705 | n69220;
  assign n69356 = (n68389 & n69354) | (n68389 & n69355) | (n69354 & n69355);
  assign n28228 = ~n69353 & n69356;
  assign n28229 = x161 & x179;
  assign n28230 = n28228 & n28229;
  assign n28231 = n28228 | n28229;
  assign n28232 = ~n28230 & n28231;
  assign n69357 = n27428 | n27825;
  assign n69358 = (n27825 & n27827) | (n27825 & n69357) | (n27827 & n69357);
  assign n54707 = n28232 & n69358;
  assign n54692 = n27825 | n27827;
  assign n54708 = n28232 & n54692;
  assign n69359 = (n54309 & n54707) | (n54309 & n54708) | (n54707 & n54708);
  assign n69360 = (n54707 & n54708) | (n54707 & n69108) | (n54708 & n69108);
  assign n69361 = (n68776 & n69359) | (n68776 & n69360) | (n69359 & n69360);
  assign n54710 = n28232 | n69358;
  assign n54711 = n28232 | n54692;
  assign n69362 = (n54309 & n54710) | (n54309 & n54711) | (n54710 & n54711);
  assign n69363 = (n54710 & n54711) | (n54710 & n69108) | (n54711 & n69108);
  assign n69364 = (n68776 & n69362) | (n68776 & n69363) | (n69362 & n69363);
  assign n28235 = ~n69361 & n69364;
  assign n28236 = x160 & x180;
  assign n28237 = n28235 & n28236;
  assign n28238 = n28235 | n28236;
  assign n28239 = ~n28237 & n28238;
  assign n69332 = n27832 | n27834;
  assign n69333 = (n27832 & n69237) | (n27832 & n69332) | (n69237 & n69332);
  assign n69365 = n28239 & n69333;
  assign n69334 = (n27832 & n69239) | (n27832 & n69332) | (n69239 & n69332);
  assign n69366 = n28239 & n69334;
  assign n69367 = (n68982 & n69365) | (n68982 & n69366) | (n69365 & n69366);
  assign n69368 = n28239 | n69333;
  assign n69369 = n28239 | n69334;
  assign n69370 = (n68982 & n69368) | (n68982 & n69369) | (n69368 & n69369);
  assign n28242 = ~n69367 & n69370;
  assign n28243 = x159 & x181;
  assign n28244 = n28242 & n28243;
  assign n28245 = n28242 | n28243;
  assign n28246 = ~n28244 & n28245;
  assign n69371 = n27839 | n27841;
  assign n69372 = (n27839 & n54476) | (n27839 & n69371) | (n54476 & n69371);
  assign n54713 = n28246 & n69372;
  assign n69373 = n27442 | n27839;
  assign n69374 = (n27839 & n27841) | (n27839 & n69373) | (n27841 & n69373);
  assign n54714 = n28246 & n69374;
  assign n54715 = (n69084 & n54713) | (n69084 & n54714) | (n54713 & n54714);
  assign n54716 = n28246 | n69372;
  assign n54717 = n28246 | n69374;
  assign n54718 = (n69084 & n54716) | (n69084 & n54717) | (n54716 & n54717);
  assign n28249 = ~n54715 & n54718;
  assign n28250 = x158 & x182;
  assign n28251 = n28249 & n28250;
  assign n28252 = n28249 | n28250;
  assign n28253 = ~n28251 & n28252;
  assign n54719 = n27846 & n28253;
  assign n54720 = (n28253 & n69244) | (n28253 & n54719) | (n69244 & n54719);
  assign n54721 = n27846 | n28253;
  assign n54722 = n69244 | n54721;
  assign n28256 = ~n54720 & n54722;
  assign n28257 = x157 & x183;
  assign n28258 = n28256 & n28257;
  assign n28259 = n28256 | n28257;
  assign n28260 = ~n28258 & n28259;
  assign n28261 = n69331 & n28260;
  assign n28262 = n69331 | n28260;
  assign n28263 = ~n28261 & n28262;
  assign n28264 = x156 & x184;
  assign n28265 = n28263 & n28264;
  assign n28266 = n28263 | n28264;
  assign n28267 = ~n28265 & n28266;
  assign n54680 = n27860 | n27862;
  assign n54723 = n28267 & n54680;
  assign n54724 = n27860 & n28267;
  assign n54725 = (n69197 & n54723) | (n69197 & n54724) | (n54723 & n54724);
  assign n54726 = n28267 | n54680;
  assign n54727 = n27860 | n28267;
  assign n54728 = (n69197 & n54726) | (n69197 & n54727) | (n54726 & n54727);
  assign n28270 = ~n54725 & n54728;
  assign n28271 = x155 & x185;
  assign n28272 = n28270 & n28271;
  assign n28273 = n28270 | n28271;
  assign n28274 = ~n28272 & n28273;
  assign n54678 = n27867 | n54527;
  assign n69375 = n28274 & n54678;
  assign n69323 = n27470 | n27867;
  assign n69324 = (n27867 & n27869) | (n27867 & n69323) | (n27869 & n69323);
  assign n69376 = n28274 & n69324;
  assign n69377 = (n54276 & n69375) | (n54276 & n69376) | (n69375 & n69376);
  assign n69378 = n28274 | n54678;
  assign n69379 = n28274 | n69324;
  assign n69380 = (n54276 & n69378) | (n54276 & n69379) | (n69378 & n69379);
  assign n28277 = ~n69377 & n69380;
  assign n28278 = x154 & x186;
  assign n28279 = n28277 & n28278;
  assign n28280 = n28277 | n28278;
  assign n28281 = ~n28279 & n28280;
  assign n54675 = n27874 | n27876;
  assign n54729 = n28281 & n54675;
  assign n54730 = n27874 & n28281;
  assign n69381 = (n54464 & n54729) | (n54464 & n54730) | (n54729 & n54730);
  assign n69382 = (n54729 & n54730) | (n54729 & n69190) | (n54730 & n69190);
  assign n69383 = (n54142 & n69381) | (n54142 & n69382) | (n69381 & n69382);
  assign n54732 = n28281 | n54675;
  assign n54733 = n27874 | n28281;
  assign n69384 = (n54464 & n54732) | (n54464 & n54733) | (n54732 & n54733);
  assign n69385 = (n54732 & n54733) | (n54732 & n69190) | (n54733 & n69190);
  assign n69386 = (n54142 & n69384) | (n54142 & n69385) | (n69384 & n69385);
  assign n28284 = ~n69383 & n69386;
  assign n28285 = x153 & x187;
  assign n28286 = n28284 & n28285;
  assign n28287 = n28284 | n28285;
  assign n28288 = ~n28286 & n28287;
  assign n54735 = n27881 & n28288;
  assign n54736 = (n28288 & n54535) | (n28288 & n54735) | (n54535 & n54735);
  assign n54737 = n27881 | n28288;
  assign n54738 = n54535 | n54737;
  assign n28291 = ~n54736 & n54738;
  assign n28292 = x152 & x188;
  assign n28293 = n28291 & n28292;
  assign n28294 = n28291 | n28292;
  assign n28295 = ~n28293 & n28294;
  assign n28296 = n69322 & n28295;
  assign n28297 = n69322 | n28295;
  assign n28298 = ~n28296 & n28297;
  assign n28299 = x151 & x189;
  assign n28300 = n28298 & n28299;
  assign n28301 = n28298 | n28299;
  assign n28302 = ~n28300 & n28301;
  assign n54670 = n27895 | n27897;
  assign n54739 = n28302 & n54670;
  assign n54740 = n27895 & n28302;
  assign n54741 = (n54460 & n54739) | (n54460 & n54740) | (n54739 & n54740);
  assign n54742 = n28302 | n54670;
  assign n54743 = n27895 | n28302;
  assign n54744 = (n54460 & n54742) | (n54460 & n54743) | (n54742 & n54743);
  assign n28305 = ~n54741 & n54744;
  assign n28306 = x150 & x190;
  assign n28307 = n28305 & n28306;
  assign n28308 = n28305 | n28306;
  assign n28309 = ~n28307 & n28308;
  assign n54745 = n27902 & n28309;
  assign n54746 = (n28309 & n54545) | (n28309 & n54745) | (n54545 & n54745);
  assign n54747 = n27902 | n28309;
  assign n54748 = n54545 | n54747;
  assign n28312 = ~n54746 & n54748;
  assign n28313 = x149 & x191;
  assign n28314 = n28312 & n28313;
  assign n28315 = n28312 | n28313;
  assign n28316 = ~n28314 & n28315;
  assign n28317 = n69317 & n28316;
  assign n28318 = n69317 | n28316;
  assign n28319 = ~n28317 & n28318;
  assign n28320 = x148 & x192;
  assign n28321 = n28319 & n28320;
  assign n28322 = n28319 | n28320;
  assign n28323 = ~n28321 & n28322;
  assign n54665 = n27916 | n27918;
  assign n54749 = n28323 & n54665;
  assign n54750 = n27916 & n28323;
  assign n54751 = (n69186 & n54749) | (n69186 & n54750) | (n54749 & n54750);
  assign n54752 = n28323 | n54665;
  assign n54753 = n27916 | n28323;
  assign n54754 = (n69186 & n54752) | (n69186 & n54753) | (n54752 & n54753);
  assign n28326 = ~n54751 & n54754;
  assign n28327 = x147 & x193;
  assign n28328 = n28326 & n28327;
  assign n28329 = n28326 | n28327;
  assign n28330 = ~n28328 & n28329;
  assign n54755 = n27923 & n28330;
  assign n69387 = (n28330 & n54554) | (n28330 & n54755) | (n54554 & n54755);
  assign n69388 = (n28330 & n54553) | (n28330 & n54755) | (n54553 & n54755);
  assign n69389 = (n69065 & n69387) | (n69065 & n69388) | (n69387 & n69388);
  assign n54757 = n27923 | n28330;
  assign n69390 = n54554 | n54757;
  assign n69391 = n54553 | n54757;
  assign n69392 = (n69065 & n69390) | (n69065 & n69391) | (n69390 & n69391);
  assign n28333 = ~n69389 & n69392;
  assign n28334 = x146 & x194;
  assign n28335 = n28333 & n28334;
  assign n28336 = n28333 | n28334;
  assign n28337 = ~n28335 & n28336;
  assign n28338 = n69312 & n28337;
  assign n28339 = n69312 | n28337;
  assign n28340 = ~n28338 & n28339;
  assign n28341 = x145 & x195;
  assign n28342 = n28340 & n28341;
  assign n28343 = n28340 | n28341;
  assign n28344 = ~n28342 & n28343;
  assign n54660 = n27937 | n27939;
  assign n54759 = n28344 & n54660;
  assign n54760 = n27937 & n28344;
  assign n54761 = (n69181 & n54759) | (n69181 & n54760) | (n54759 & n54760);
  assign n54762 = n28344 | n54660;
  assign n54763 = n27937 | n28344;
  assign n54764 = (n69181 & n54762) | (n69181 & n54763) | (n54762 & n54763);
  assign n28347 = ~n54761 & n54764;
  assign n28348 = x144 & x196;
  assign n28349 = n28347 & n28348;
  assign n28350 = n28347 | n28348;
  assign n28351 = ~n28349 & n28350;
  assign n54765 = n27944 & n28351;
  assign n69393 = (n28351 & n54564) | (n28351 & n54765) | (n54564 & n54765);
  assign n69394 = (n28351 & n54563) | (n28351 & n54765) | (n54563 & n54765);
  assign n69395 = (n54258 & n69393) | (n54258 & n69394) | (n69393 & n69394);
  assign n54767 = n27944 | n28351;
  assign n69396 = n54564 | n54767;
  assign n69397 = n54563 | n54767;
  assign n69398 = (n54258 & n69396) | (n54258 & n69397) | (n69396 & n69397);
  assign n28354 = ~n69395 & n69398;
  assign n28355 = x143 & x197;
  assign n28356 = n28354 & n28355;
  assign n28357 = n28354 | n28355;
  assign n28358 = ~n28356 & n28357;
  assign n54658 = n27951 | n27953;
  assign n69399 = n28358 & n54658;
  assign n69306 = n27554 | n27951;
  assign n69307 = (n27951 & n27953) | (n27951 & n69306) | (n27953 & n69306);
  assign n69400 = n28358 & n69307;
  assign n69401 = (n69157 & n69399) | (n69157 & n69400) | (n69399 & n69400);
  assign n69402 = n28358 | n54658;
  assign n69403 = n28358 | n69307;
  assign n69404 = (n69157 & n69402) | (n69157 & n69403) | (n69402 & n69403);
  assign n28361 = ~n69401 & n69404;
  assign n28362 = x142 & x198;
  assign n28363 = n28361 & n28362;
  assign n28364 = n28361 | n28362;
  assign n28365 = ~n28363 & n28364;
  assign n54769 = n27958 & n28365;
  assign n69405 = (n28365 & n54573) | (n28365 & n54769) | (n54573 & n54769);
  assign n69406 = (n27960 & n28365) | (n27960 & n54769) | (n28365 & n54769);
  assign n69407 = (n54369 & n69405) | (n54369 & n69406) | (n69405 & n69406);
  assign n54771 = n27958 | n28365;
  assign n69408 = n54573 | n54771;
  assign n69409 = n27960 | n54771;
  assign n69410 = (n54369 & n69408) | (n54369 & n69409) | (n69408 & n69409);
  assign n28368 = ~n69407 & n69410;
  assign n28369 = x141 & x199;
  assign n28370 = n28368 & n28369;
  assign n28371 = n28368 | n28369;
  assign n28372 = ~n28370 & n28371;
  assign n54773 = n27965 & n28372;
  assign n54774 = (n28372 & n54578) | (n28372 & n54773) | (n54578 & n54773);
  assign n54775 = n27965 | n28372;
  assign n54776 = n54578 | n54775;
  assign n28375 = ~n54774 & n54776;
  assign n28376 = x140 & x200;
  assign n28377 = n28375 & n28376;
  assign n28378 = n28375 | n28376;
  assign n28379 = ~n28377 & n28378;
  assign n54777 = n27972 & n28379;
  assign n54778 = (n28379 & n54582) | (n28379 & n54777) | (n54582 & n54777);
  assign n54779 = n27972 | n28379;
  assign n54780 = n54582 | n54779;
  assign n28382 = ~n54778 & n54780;
  assign n28383 = x139 & x201;
  assign n28384 = n28382 & n28383;
  assign n28385 = n28382 | n28383;
  assign n28386 = ~n28384 & n28385;
  assign n54781 = n27979 & n28386;
  assign n54782 = (n28386 & n54586) | (n28386 & n54781) | (n54586 & n54781);
  assign n54783 = n27979 | n28386;
  assign n54784 = n54586 | n54783;
  assign n28389 = ~n54782 & n54784;
  assign n28390 = x138 & x202;
  assign n28391 = n28389 & n28390;
  assign n28392 = n28389 | n28390;
  assign n28393 = ~n28391 & n28392;
  assign n54785 = n27986 & n28393;
  assign n54786 = (n28393 & n54590) | (n28393 & n54785) | (n54590 & n54785);
  assign n54787 = n27986 | n28393;
  assign n54788 = n54590 | n54787;
  assign n28396 = ~n54786 & n54788;
  assign n28397 = x137 & x203;
  assign n28398 = n28396 & n28397;
  assign n28399 = n28396 | n28397;
  assign n28400 = ~n28398 & n28399;
  assign n54789 = n27993 & n28400;
  assign n54790 = (n28400 & n54594) | (n28400 & n54789) | (n54594 & n54789);
  assign n54791 = n27993 | n28400;
  assign n54792 = n54594 | n54791;
  assign n28403 = ~n54790 & n54792;
  assign n28404 = x136 & x204;
  assign n28405 = n28403 & n28404;
  assign n28406 = n28403 | n28404;
  assign n28407 = ~n28405 & n28406;
  assign n54793 = n28000 & n28407;
  assign n54794 = (n28407 & n54598) | (n28407 & n54793) | (n54598 & n54793);
  assign n54795 = n28000 | n28407;
  assign n54796 = n54598 | n54795;
  assign n28410 = ~n54794 & n54796;
  assign n28411 = x135 & x205;
  assign n28412 = n28410 & n28411;
  assign n28413 = n28410 | n28411;
  assign n28414 = ~n28412 & n28413;
  assign n54797 = n28007 & n28414;
  assign n54798 = (n28414 & n54602) | (n28414 & n54797) | (n54602 & n54797);
  assign n54799 = n28007 | n28414;
  assign n54800 = n54602 | n54799;
  assign n28417 = ~n54798 & n54800;
  assign n28418 = x134 & x206;
  assign n28419 = n28417 & n28418;
  assign n28420 = n28417 | n28418;
  assign n28421 = ~n28419 & n28420;
  assign n54801 = n28014 & n28421;
  assign n54802 = (n28421 & n54606) | (n28421 & n54801) | (n54606 & n54801);
  assign n54803 = n28014 | n28421;
  assign n54804 = n54606 | n54803;
  assign n28424 = ~n54802 & n54804;
  assign n28425 = x133 & x207;
  assign n28426 = n28424 & n28425;
  assign n28427 = n28424 | n28425;
  assign n28428 = ~n28426 & n28427;
  assign n54805 = n28021 & n28428;
  assign n54806 = (n28428 & n54610) | (n28428 & n54805) | (n54610 & n54805);
  assign n54807 = n28021 | n28428;
  assign n54808 = n54610 | n54807;
  assign n28431 = ~n54806 & n54808;
  assign n28432 = x132 & x208;
  assign n28433 = n28431 & n28432;
  assign n28434 = n28431 | n28432;
  assign n28435 = ~n28433 & n28434;
  assign n54809 = n28028 & n28435;
  assign n54810 = (n28435 & n54614) | (n28435 & n54809) | (n54614 & n54809);
  assign n54811 = n28028 | n28435;
  assign n54812 = n54614 | n54811;
  assign n28438 = ~n54810 & n54812;
  assign n28439 = x131 & x209;
  assign n28440 = n28438 & n28439;
  assign n28441 = n28438 | n28439;
  assign n28442 = ~n28440 & n28441;
  assign n54813 = n28035 & n28442;
  assign n54814 = (n28442 & n54618) | (n28442 & n54813) | (n54618 & n54813);
  assign n54815 = n28035 | n28442;
  assign n54816 = n54618 | n54815;
  assign n28445 = ~n54814 & n54816;
  assign n28446 = x130 & x210;
  assign n28447 = n28445 & n28446;
  assign n28448 = n28445 | n28446;
  assign n28449 = ~n28447 & n28448;
  assign n54817 = n28042 & n28449;
  assign n54818 = (n28449 & n54623) | (n28449 & n54817) | (n54623 & n54817);
  assign n54819 = n28042 | n28449;
  assign n54820 = n54623 | n54819;
  assign n28452 = ~n54818 & n54820;
  assign n28453 = x129 & x211;
  assign n28454 = n28452 & n28453;
  assign n28455 = n28452 | n28453;
  assign n28456 = ~n28454 & n28455;
  assign n54655 = n28049 | n28051;
  assign n54821 = n28456 & n54655;
  assign n54822 = n28049 & n28456;
  assign n54823 = (n54443 & n54821) | (n54443 & n54822) | (n54821 & n54822);
  assign n54824 = n28456 | n54655;
  assign n54825 = n28049 | n28456;
  assign n54826 = (n54443 & n54824) | (n54443 & n54825) | (n54824 & n54825);
  assign n28459 = ~n54823 & n54826;
  assign n28460 = x128 & x212;
  assign n28461 = n28459 & n28460;
  assign n28462 = n28459 | n28460;
  assign n28463 = ~n28461 & n28462;
  assign n54653 = n28056 | n28058;
  assign n69411 = n28463 & n54653;
  assign n69412 = n28056 & n28463;
  assign n69413 = (n54441 & n69411) | (n54441 & n69412) | (n69411 & n69412);
  assign n69414 = n28463 | n54653;
  assign n69415 = n28056 | n28463;
  assign n69416 = (n54441 & n69414) | (n54441 & n69415) | (n69414 & n69415);
  assign n28466 = ~n69413 & n69416;
  assign n28467 = x127 & x213;
  assign n28468 = n28466 & n28467;
  assign n28469 = n28466 | n28467;
  assign n28470 = ~n28468 & n28469;
  assign n54651 = n28063 | n28065;
  assign n69417 = n28470 & n54651;
  assign n69418 = n28063 & n28470;
  assign n69419 = (n54439 & n69417) | (n54439 & n69418) | (n69417 & n69418);
  assign n69420 = n28470 | n54651;
  assign n69421 = n28063 | n28470;
  assign n69422 = (n54439 & n69420) | (n54439 & n69421) | (n69420 & n69421);
  assign n28473 = ~n69419 & n69422;
  assign n28474 = x126 & x214;
  assign n28475 = n28473 & n28474;
  assign n28476 = n28473 | n28474;
  assign n28477 = ~n28475 & n28476;
  assign n28478 = n54650 & n28477;
  assign n28479 = n54650 | n28477;
  assign n28480 = ~n28478 & n28479;
  assign n28481 = x125 & x215;
  assign n28482 = n28480 & n28481;
  assign n28483 = n28480 | n28481;
  assign n28484 = ~n28482 & n28483;
  assign n28485 = n54648 & n28484;
  assign n28486 = n54648 | n28484;
  assign n28487 = ~n28485 & n28486;
  assign n28488 = x124 & x216;
  assign n28489 = n28487 & n28488;
  assign n28490 = n28487 | n28488;
  assign n28491 = ~n28489 & n28490;
  assign n28492 = n54646 & n28491;
  assign n28493 = n54646 | n28491;
  assign n28494 = ~n28492 & n28493;
  assign n28495 = x123 & x217;
  assign n28496 = n28494 & n28495;
  assign n28497 = n28494 | n28495;
  assign n28498 = ~n28496 & n28497;
  assign n28499 = n54644 & n28498;
  assign n28500 = n54644 | n28498;
  assign n28501 = ~n28499 & n28500;
  assign n28502 = x122 & x218;
  assign n28503 = n28501 & n28502;
  assign n28504 = n28501 | n28502;
  assign n28505 = ~n28503 & n28504;
  assign n28506 = n69305 & n28505;
  assign n28507 = n69305 | n28505;
  assign n28508 = ~n28506 & n28507;
  assign n28509 = x121 & x219;
  assign n28510 = n28508 & n28509;
  assign n28511 = n28508 | n28509;
  assign n28512 = ~n28510 & n28511;
  assign n28513 = n54642 & n28512;
  assign n28514 = n54642 | n28512;
  assign n28515 = ~n28513 & n28514;
  assign n28516 = x120 & x220;
  assign n28517 = n28515 & n28516;
  assign n28518 = n28515 | n28516;
  assign n28519 = ~n28517 & n28518;
  assign n28520 = n54640 & n28519;
  assign n28521 = n54640 | n28519;
  assign n28522 = ~n28520 & n28521;
  assign n28523 = x119 & x221;
  assign n28524 = n28522 & n28523;
  assign n28525 = n28522 | n28523;
  assign n28526 = ~n28524 & n28525;
  assign n28527 = n54638 & n28526;
  assign n28528 = n54638 | n28526;
  assign n28529 = ~n28527 & n28528;
  assign n28530 = x118 & x222;
  assign n28531 = n28529 & n28530;
  assign n28532 = n28529 | n28530;
  assign n28533 = ~n28531 & n28532;
  assign n28534 = n54636 & n28533;
  assign n28535 = n54636 | n28533;
  assign n28536 = ~n28534 & n28535;
  assign n28537 = x117 & x223;
  assign n28538 = n28536 & n28537;
  assign n28539 = n28536 | n28537;
  assign n28540 = ~n28538 & n28539;
  assign n28541 = n54634 & n28540;
  assign n28542 = n54634 | n28540;
  assign n28543 = ~n28541 & n28542;
  assign n28544 = x116 & x224;
  assign n28545 = n28543 & n28544;
  assign n28546 = n28543 | n28544;
  assign n28547 = ~n28545 & n28546;
  assign n28548 = n54632 & n28547;
  assign n28549 = n54632 | n28547;
  assign n28550 = ~n28548 & n28549;
  assign n28551 = x115 & x225;
  assign n28552 = n28550 & n28551;
  assign n28553 = n28550 | n28551;
  assign n28554 = ~n28552 & n28553;
  assign n28555 = n54630 & n28554;
  assign n28556 = n54630 | n28554;
  assign n28557 = ~n28555 & n28556;
  assign n28558 = x114 & x226;
  assign n28559 = n28557 & n28558;
  assign n28560 = n28557 | n28558;
  assign n28561 = ~n28559 & n28560;
  assign n28562 = n54628 & n28561;
  assign n28563 = n54628 | n28561;
  assign n28564 = ~n28562 & n28563;
  assign n28565 = x113 & x227;
  assign n28566 = n28564 & n28565;
  assign n28567 = n28564 | n28565;
  assign n28568 = ~n28566 & n28567;
  assign n28569 = n28161 & n28568;
  assign n28570 = n28161 | n28568;
  assign n28571 = ~n28569 & n28570;
  assign n28572 = x112 & x228;
  assign n28573 = n28571 & n28572;
  assign n28574 = n28571 | n28572;
  assign n28575 = ~n28573 & n28574;
  assign n54827 = n28161 | n28566;
  assign n54828 = (n28566 & n28568) | (n28566 & n54827) | (n28568 & n54827);
  assign n54829 = n28559 | n54628;
  assign n54830 = (n28559 & n28561) | (n28559 & n54829) | (n28561 & n54829);
  assign n54831 = n28552 | n54630;
  assign n54832 = (n28552 & n28554) | (n28552 & n54831) | (n28554 & n54831);
  assign n54833 = n28545 | n54632;
  assign n54834 = (n28545 & n28547) | (n28545 & n54833) | (n28547 & n54833);
  assign n54835 = n28538 | n54634;
  assign n54836 = (n28538 & n28540) | (n28538 & n54835) | (n28540 & n54835);
  assign n54837 = n28531 | n54636;
  assign n54838 = (n28531 & n28533) | (n28531 & n54837) | (n28533 & n54837);
  assign n54839 = n28524 | n54638;
  assign n54840 = (n28524 & n28526) | (n28524 & n54839) | (n28526 & n54839);
  assign n54841 = n28517 | n54640;
  assign n54842 = (n28517 & n28519) | (n28517 & n54841) | (n28519 & n54841);
  assign n54843 = n28510 | n54642;
  assign n54844 = (n28510 & n28512) | (n28510 & n54843) | (n28512 & n54843);
  assign n54845 = n28503 | n28505;
  assign n54846 = (n69305 & n28503) | (n69305 & n54845) | (n28503 & n54845);
  assign n54847 = n28496 | n28498;
  assign n54848 = (n28496 & n54644) | (n28496 & n54847) | (n54644 & n54847);
  assign n54849 = n28489 | n28491;
  assign n54850 = (n28489 & n54646) | (n28489 & n54849) | (n54646 & n54849);
  assign n54851 = n28482 | n28484;
  assign n54852 = (n28482 & n54648) | (n28482 & n54851) | (n54648 & n54851);
  assign n54652 = (n28063 & n54439) | (n28063 & n54651) | (n54439 & n54651);
  assign n54654 = (n28056 & n54441) | (n28056 & n54653) | (n54441 & n54653);
  assign n54659 = (n69157 & n69307) | (n69157 & n54658) | (n69307 & n54658);
  assign n54862 = n28349 | n28351;
  assign n69423 = n27944 | n28349;
  assign n69424 = (n28349 & n28351) | (n28349 & n69423) | (n28351 & n69423);
  assign n69425 = (n54564 & n54862) | (n54564 & n69424) | (n54862 & n69424);
  assign n69426 = (n54563 & n54862) | (n54563 & n69424) | (n54862 & n69424);
  assign n69427 = (n54258 & n69425) | (n54258 & n69426) | (n69425 & n69426);
  assign n54867 = n28328 | n28330;
  assign n69428 = n27923 | n28328;
  assign n69429 = (n28328 & n28330) | (n28328 & n69428) | (n28330 & n69428);
  assign n69430 = (n54554 & n54867) | (n54554 & n69429) | (n54867 & n69429);
  assign n69431 = (n54553 & n54867) | (n54553 & n69429) | (n54867 & n69429);
  assign n69432 = (n69065 & n69430) | (n69065 & n69431) | (n69430 & n69431);
  assign n54465 = (n54142 & n69190) | (n54142 & n54464) | (n69190 & n54464);
  assign n28627 = x165 & x176;
  assign n28628 = x164 & x177;
  assign n28629 = n28627 & n28628;
  assign n28630 = n28627 | n28628;
  assign n28631 = ~n28629 & n28630;
  assign n69441 = n28216 | n69335;
  assign n69444 = n28631 & n69441;
  assign n69442 = n28216 | n28218;
  assign n69445 = n28631 & n69442;
  assign n69446 = (n69202 & n69444) | (n69202 & n69445) | (n69444 & n69445);
  assign n69447 = n28216 & n28631;
  assign n69448 = (n28631 & n69340) | (n28631 & n69447) | (n69340 & n69447);
  assign n69449 = (n53919 & n69446) | (n53919 & n69448) | (n69446 & n69448);
  assign n69450 = (n53918 & n69446) | (n53918 & n69448) | (n69446 & n69448);
  assign n69451 = (n68195 & n69449) | (n68195 & n69450) | (n69449 & n69450);
  assign n69452 = n28631 | n69441;
  assign n69453 = n28631 | n69442;
  assign n69454 = (n69202 & n69452) | (n69202 & n69453) | (n69452 & n69453);
  assign n69455 = n28216 | n28631;
  assign n69456 = n69340 | n69455;
  assign n69457 = (n53919 & n69454) | (n53919 & n69456) | (n69454 & n69456);
  assign n69458 = (n53918 & n69454) | (n53918 & n69456) | (n69454 & n69456);
  assign n69459 = (n68195 & n69457) | (n68195 & n69458) | (n69457 & n69458);
  assign n28634 = ~n69451 & n69459;
  assign n28635 = x163 & x178;
  assign n28636 = n28634 & n28635;
  assign n28637 = n28634 | n28635;
  assign n28638 = ~n28636 & n28637;
  assign n69460 = n27818 | n28223;
  assign n69461 = (n28223 & n28225) | (n28223 & n69460) | (n28225 & n69460);
  assign n54909 = n28638 & n69461;
  assign n54898 = n28223 | n28225;
  assign n54910 = n28638 & n54898;
  assign n69462 = (n54909 & n54910) | (n54909 & n69221) | (n54910 & n69221);
  assign n69463 = (n54909 & n54910) | (n54909 & n69220) | (n54910 & n69220);
  assign n69464 = (n68389 & n69462) | (n68389 & n69463) | (n69462 & n69463);
  assign n54912 = n28638 | n69461;
  assign n54913 = n28638 | n54898;
  assign n69465 = (n54912 & n54913) | (n54912 & n69221) | (n54913 & n69221);
  assign n69466 = (n54912 & n54913) | (n54912 & n69220) | (n54913 & n69220);
  assign n69467 = (n68389 & n69465) | (n68389 & n69466) | (n69465 & n69466);
  assign n28641 = ~n69464 & n69467;
  assign n28642 = x162 & x179;
  assign n28643 = n28641 & n28642;
  assign n28644 = n28641 | n28642;
  assign n28645 = ~n28643 & n28644;
  assign n69468 = n28230 | n28232;
  assign n69469 = (n28230 & n69358) | (n28230 & n69468) | (n69358 & n69468);
  assign n54915 = n28645 & n69469;
  assign n69470 = (n28230 & n54692) | (n28230 & n69468) | (n54692 & n69468);
  assign n54916 = n28645 & n69470;
  assign n69471 = (n54309 & n54915) | (n54309 & n54916) | (n54915 & n54916);
  assign n69472 = (n54915 & n54916) | (n54915 & n69108) | (n54916 & n69108);
  assign n69473 = (n68776 & n69471) | (n68776 & n69472) | (n69471 & n69472);
  assign n54918 = n28645 | n69469;
  assign n54919 = n28645 | n69470;
  assign n69474 = (n54309 & n54918) | (n54309 & n54919) | (n54918 & n54919);
  assign n69475 = (n54918 & n54919) | (n54918 & n69108) | (n54919 & n69108);
  assign n69476 = (n68776 & n69474) | (n68776 & n69475) | (n69474 & n69475);
  assign n28648 = ~n69473 & n69476;
  assign n28649 = x161 & x180;
  assign n28650 = n28648 & n28649;
  assign n28651 = n28648 | n28649;
  assign n28652 = ~n28650 & n28651;
  assign n54892 = n28237 | n28239;
  assign n54921 = n28652 & n54892;
  assign n54922 = n28237 & n28652;
  assign n69477 = (n54921 & n54922) | (n54921 & n69333) | (n54922 & n69333);
  assign n69478 = (n54921 & n54922) | (n54921 & n69334) | (n54922 & n69334);
  assign n69479 = (n68982 & n69477) | (n68982 & n69478) | (n69477 & n69478);
  assign n54924 = n28652 | n54892;
  assign n54925 = n28237 | n28652;
  assign n69480 = (n54924 & n54925) | (n54924 & n69333) | (n54925 & n69333);
  assign n69481 = (n54924 & n54925) | (n54924 & n69334) | (n54925 & n69334);
  assign n69482 = (n68982 & n69480) | (n68982 & n69481) | (n69480 & n69481);
  assign n28655 = ~n69479 & n69482;
  assign n28656 = x160 & x181;
  assign n28657 = n28655 & n28656;
  assign n28658 = n28655 | n28656;
  assign n28659 = ~n28657 & n28658;
  assign n54927 = n28244 & n28659;
  assign n69483 = (n28659 & n54713) | (n28659 & n54927) | (n54713 & n54927);
  assign n69484 = (n28659 & n54714) | (n28659 & n54927) | (n54714 & n54927);
  assign n69485 = (n69084 & n69483) | (n69084 & n69484) | (n69483 & n69484);
  assign n54929 = n28244 | n28659;
  assign n69486 = n54713 | n54929;
  assign n69487 = n54714 | n54929;
  assign n69488 = (n69084 & n69486) | (n69084 & n69487) | (n69486 & n69487);
  assign n28662 = ~n69485 & n69488;
  assign n28663 = x159 & x182;
  assign n28664 = n28662 & n28663;
  assign n28665 = n28662 | n28663;
  assign n28666 = ~n28664 & n28665;
  assign n69489 = n27846 | n28251;
  assign n69490 = (n28251 & n28253) | (n28251 & n69489) | (n28253 & n69489);
  assign n54931 = n28666 & n69490;
  assign n54890 = n28251 | n28253;
  assign n54932 = n28666 & n54890;
  assign n54933 = (n69244 & n54931) | (n69244 & n54932) | (n54931 & n54932);
  assign n54934 = n28666 | n69490;
  assign n54935 = n28666 | n54890;
  assign n54936 = (n69244 & n54934) | (n69244 & n54935) | (n54934 & n54935);
  assign n28669 = ~n54933 & n54936;
  assign n28670 = x158 & x183;
  assign n28671 = n28669 & n28670;
  assign n28672 = n28669 | n28670;
  assign n28673 = ~n28671 & n28672;
  assign n54887 = n28258 | n28260;
  assign n54937 = n28673 & n54887;
  assign n54938 = n28258 & n28673;
  assign n54939 = (n69331 & n54937) | (n69331 & n54938) | (n54937 & n54938);
  assign n54940 = n28673 | n54887;
  assign n54941 = n28258 | n28673;
  assign n54942 = (n69331 & n54940) | (n69331 & n54941) | (n54940 & n54941);
  assign n28676 = ~n54939 & n54942;
  assign n28677 = x157 & x184;
  assign n28678 = n28676 & n28677;
  assign n28679 = n28676 | n28677;
  assign n28680 = ~n28678 & n28679;
  assign n54885 = n28265 | n54723;
  assign n69491 = n28680 & n54885;
  assign n69439 = n27860 | n28265;
  assign n69440 = (n28265 & n28267) | (n28265 & n69439) | (n28267 & n69439);
  assign n69492 = n28680 & n69440;
  assign n69493 = (n69197 & n69491) | (n69197 & n69492) | (n69491 & n69492);
  assign n69494 = n28680 | n54885;
  assign n69495 = n28680 | n69440;
  assign n69496 = (n69197 & n69494) | (n69197 & n69495) | (n69494 & n69495);
  assign n28683 = ~n69493 & n69496;
  assign n28684 = x156 & x185;
  assign n28685 = n28683 & n28684;
  assign n28686 = n28683 | n28684;
  assign n28687 = ~n28685 & n28686;
  assign n54882 = n28272 | n28274;
  assign n54943 = n28687 & n54882;
  assign n54944 = n28272 & n28687;
  assign n69497 = (n54678 & n54943) | (n54678 & n54944) | (n54943 & n54944);
  assign n69498 = (n54943 & n54944) | (n54943 & n69324) | (n54944 & n69324);
  assign n69499 = (n54276 & n69497) | (n54276 & n69498) | (n69497 & n69498);
  assign n54946 = n28687 | n54882;
  assign n54947 = n28272 | n28687;
  assign n69500 = (n54678 & n54946) | (n54678 & n54947) | (n54946 & n54947);
  assign n69501 = (n54946 & n54947) | (n54946 & n69324) | (n54947 & n69324);
  assign n69502 = (n54276 & n69500) | (n54276 & n69501) | (n69500 & n69501);
  assign n28690 = ~n69499 & n69502;
  assign n28691 = x155 & x186;
  assign n28692 = n28690 & n28691;
  assign n28693 = n28690 | n28691;
  assign n28694 = ~n28692 & n28693;
  assign n54880 = n28279 | n54729;
  assign n69503 = n28694 & n54880;
  assign n69437 = n27874 | n28279;
  assign n69438 = (n28279 & n28281) | (n28279 & n69437) | (n28281 & n69437);
  assign n69504 = n28694 & n69438;
  assign n69505 = (n54465 & n69503) | (n54465 & n69504) | (n69503 & n69504);
  assign n69506 = n28694 | n54880;
  assign n69507 = n28694 | n69438;
  assign n69508 = (n54465 & n69506) | (n54465 & n69507) | (n69506 & n69507);
  assign n28697 = ~n69505 & n69508;
  assign n28698 = x154 & x187;
  assign n28699 = n28697 & n28698;
  assign n28700 = n28697 | n28698;
  assign n28701 = ~n28699 & n28700;
  assign n54877 = n28286 | n28288;
  assign n69509 = n28701 & n54877;
  assign n69435 = n27881 | n28286;
  assign n69436 = (n28286 & n28288) | (n28286 & n69435) | (n28288 & n69435);
  assign n69510 = n28701 & n69436;
  assign n69511 = (n54535 & n69509) | (n54535 & n69510) | (n69509 & n69510);
  assign n69512 = n28701 | n54877;
  assign n69513 = n28701 | n69436;
  assign n69514 = (n54535 & n69512) | (n54535 & n69513) | (n69512 & n69513);
  assign n28704 = ~n69511 & n69514;
  assign n28705 = x153 & x188;
  assign n28706 = n28704 & n28705;
  assign n28707 = n28704 | n28705;
  assign n28708 = ~n28706 & n28707;
  assign n54874 = n28293 | n28295;
  assign n54949 = n28708 & n54874;
  assign n54950 = n28293 & n28708;
  assign n54951 = (n69322 & n54949) | (n69322 & n54950) | (n54949 & n54950);
  assign n54952 = n28708 | n54874;
  assign n54953 = n28293 | n28708;
  assign n54954 = (n69322 & n54952) | (n69322 & n54953) | (n54952 & n54953);
  assign n28711 = ~n54951 & n54954;
  assign n28712 = x152 & x189;
  assign n28713 = n28711 & n28712;
  assign n28714 = n28711 | n28712;
  assign n28715 = ~n28713 & n28714;
  assign n54955 = n28300 & n28715;
  assign n69515 = (n28715 & n54740) | (n28715 & n54955) | (n54740 & n54955);
  assign n69516 = (n28715 & n54739) | (n28715 & n54955) | (n54739 & n54955);
  assign n69517 = (n54460 & n69515) | (n54460 & n69516) | (n69515 & n69516);
  assign n54957 = n28300 | n28715;
  assign n69518 = n54740 | n54957;
  assign n69519 = n54739 | n54957;
  assign n69520 = (n54460 & n69518) | (n54460 & n69519) | (n69518 & n69519);
  assign n28718 = ~n69517 & n69520;
  assign n28719 = x151 & x190;
  assign n28720 = n28718 & n28719;
  assign n28721 = n28718 | n28719;
  assign n28722 = ~n28720 & n28721;
  assign n54872 = n28307 | n28309;
  assign n69521 = n28722 & n54872;
  assign n69433 = n27902 | n28307;
  assign n69434 = (n28307 & n28309) | (n28307 & n69433) | (n28309 & n69433);
  assign n69522 = n28722 & n69434;
  assign n69523 = (n54545 & n69521) | (n54545 & n69522) | (n69521 & n69522);
  assign n69524 = n28722 | n54872;
  assign n69525 = n28722 | n69434;
  assign n69526 = (n54545 & n69524) | (n54545 & n69525) | (n69524 & n69525);
  assign n28725 = ~n69523 & n69526;
  assign n28726 = x150 & x191;
  assign n28727 = n28725 & n28726;
  assign n28728 = n28725 | n28726;
  assign n28729 = ~n28727 & n28728;
  assign n54869 = n28314 | n28316;
  assign n54959 = n28729 & n54869;
  assign n54960 = n28314 & n28729;
  assign n54961 = (n69317 & n54959) | (n69317 & n54960) | (n54959 & n54960);
  assign n54962 = n28729 | n54869;
  assign n54963 = n28314 | n28729;
  assign n54964 = (n69317 & n54962) | (n69317 & n54963) | (n54962 & n54963);
  assign n28732 = ~n54961 & n54964;
  assign n28733 = x149 & x192;
  assign n28734 = n28732 & n28733;
  assign n28735 = n28732 | n28733;
  assign n28736 = ~n28734 & n28735;
  assign n54965 = n28321 & n28736;
  assign n69527 = (n28736 & n54750) | (n28736 & n54965) | (n54750 & n54965);
  assign n69528 = (n28736 & n54749) | (n28736 & n54965) | (n54749 & n54965);
  assign n69529 = (n69186 & n69527) | (n69186 & n69528) | (n69527 & n69528);
  assign n54967 = n28321 | n28736;
  assign n69530 = n54750 | n54967;
  assign n69531 = n54749 | n54967;
  assign n69532 = (n69186 & n69530) | (n69186 & n69531) | (n69530 & n69531);
  assign n28739 = ~n69529 & n69532;
  assign n28740 = x148 & x193;
  assign n28741 = n28739 & n28740;
  assign n28742 = n28739 | n28740;
  assign n28743 = ~n28741 & n28742;
  assign n28744 = n69432 & n28743;
  assign n28745 = n69432 | n28743;
  assign n28746 = ~n28744 & n28745;
  assign n28747 = x147 & x194;
  assign n28748 = n28746 & n28747;
  assign n28749 = n28746 | n28747;
  assign n28750 = ~n28748 & n28749;
  assign n54864 = n28335 | n28337;
  assign n54969 = n28750 & n54864;
  assign n54970 = n28335 & n28750;
  assign n54971 = (n69312 & n54969) | (n69312 & n54970) | (n54969 & n54970);
  assign n54972 = n28750 | n54864;
  assign n54973 = n28335 | n28750;
  assign n54974 = (n69312 & n54972) | (n69312 & n54973) | (n54972 & n54973);
  assign n28753 = ~n54971 & n54974;
  assign n28754 = x146 & x195;
  assign n28755 = n28753 & n28754;
  assign n28756 = n28753 | n28754;
  assign n28757 = ~n28755 & n28756;
  assign n54975 = n28342 & n28757;
  assign n69533 = (n28757 & n54760) | (n28757 & n54975) | (n54760 & n54975);
  assign n69534 = (n28757 & n54759) | (n28757 & n54975) | (n54759 & n54975);
  assign n69535 = (n69181 & n69533) | (n69181 & n69534) | (n69533 & n69534);
  assign n54977 = n28342 | n28757;
  assign n69536 = n54760 | n54977;
  assign n69537 = n54759 | n54977;
  assign n69538 = (n69181 & n69536) | (n69181 & n69537) | (n69536 & n69537);
  assign n28760 = ~n69535 & n69538;
  assign n28761 = x145 & x196;
  assign n28762 = n28760 & n28761;
  assign n28763 = n28760 | n28761;
  assign n28764 = ~n28762 & n28763;
  assign n28765 = n69427 & n28764;
  assign n28766 = n69427 | n28764;
  assign n28767 = ~n28765 & n28766;
  assign n28768 = x144 & x197;
  assign n28769 = n28767 & n28768;
  assign n28770 = n28767 | n28768;
  assign n28771 = ~n28769 & n28770;
  assign n54859 = n28356 | n28358;
  assign n54979 = n28771 & n54859;
  assign n54980 = n28356 & n28771;
  assign n54981 = (n54659 & n54979) | (n54659 & n54980) | (n54979 & n54980);
  assign n54982 = n28771 | n54859;
  assign n54983 = n28356 | n28771;
  assign n54984 = (n54659 & n54982) | (n54659 & n54983) | (n54982 & n54983);
  assign n28774 = ~n54981 & n54984;
  assign n28775 = x143 & x198;
  assign n28776 = n28774 & n28775;
  assign n28777 = n28774 | n28775;
  assign n28778 = ~n28776 & n28777;
  assign n54985 = n28363 & n28778;
  assign n54986 = (n28778 & n69407) | (n28778 & n54985) | (n69407 & n54985);
  assign n54987 = n28363 | n28778;
  assign n54988 = n69407 | n54987;
  assign n28781 = ~n54986 & n54988;
  assign n28782 = x142 & x199;
  assign n28783 = n28781 & n28782;
  assign n28784 = n28781 | n28782;
  assign n28785 = ~n28783 & n28784;
  assign n54989 = n28370 & n28785;
  assign n54990 = (n28785 & n54774) | (n28785 & n54989) | (n54774 & n54989);
  assign n54991 = n28370 | n28785;
  assign n54992 = n54774 | n54991;
  assign n28788 = ~n54990 & n54992;
  assign n28789 = x141 & x200;
  assign n28790 = n28788 & n28789;
  assign n28791 = n28788 | n28789;
  assign n28792 = ~n28790 & n28791;
  assign n54993 = n28377 & n28792;
  assign n54994 = (n28792 & n54778) | (n28792 & n54993) | (n54778 & n54993);
  assign n54995 = n28377 | n28792;
  assign n54996 = n54778 | n54995;
  assign n28795 = ~n54994 & n54996;
  assign n28796 = x140 & x201;
  assign n28797 = n28795 & n28796;
  assign n28798 = n28795 | n28796;
  assign n28799 = ~n28797 & n28798;
  assign n54997 = n28384 & n28799;
  assign n54998 = (n28799 & n54782) | (n28799 & n54997) | (n54782 & n54997);
  assign n54999 = n28384 | n28799;
  assign n55000 = n54782 | n54999;
  assign n28802 = ~n54998 & n55000;
  assign n28803 = x139 & x202;
  assign n28804 = n28802 & n28803;
  assign n28805 = n28802 | n28803;
  assign n28806 = ~n28804 & n28805;
  assign n55001 = n28391 & n28806;
  assign n55002 = (n28806 & n54786) | (n28806 & n55001) | (n54786 & n55001);
  assign n55003 = n28391 | n28806;
  assign n55004 = n54786 | n55003;
  assign n28809 = ~n55002 & n55004;
  assign n28810 = x138 & x203;
  assign n28811 = n28809 & n28810;
  assign n28812 = n28809 | n28810;
  assign n28813 = ~n28811 & n28812;
  assign n55005 = n28398 & n28813;
  assign n55006 = (n28813 & n54790) | (n28813 & n55005) | (n54790 & n55005);
  assign n55007 = n28398 | n28813;
  assign n55008 = n54790 | n55007;
  assign n28816 = ~n55006 & n55008;
  assign n28817 = x137 & x204;
  assign n28818 = n28816 & n28817;
  assign n28819 = n28816 | n28817;
  assign n28820 = ~n28818 & n28819;
  assign n55009 = n28405 & n28820;
  assign n55010 = (n28820 & n54794) | (n28820 & n55009) | (n54794 & n55009);
  assign n55011 = n28405 | n28820;
  assign n55012 = n54794 | n55011;
  assign n28823 = ~n55010 & n55012;
  assign n28824 = x136 & x205;
  assign n28825 = n28823 & n28824;
  assign n28826 = n28823 | n28824;
  assign n28827 = ~n28825 & n28826;
  assign n55013 = n28412 & n28827;
  assign n55014 = (n28827 & n54798) | (n28827 & n55013) | (n54798 & n55013);
  assign n55015 = n28412 | n28827;
  assign n55016 = n54798 | n55015;
  assign n28830 = ~n55014 & n55016;
  assign n28831 = x135 & x206;
  assign n28832 = n28830 & n28831;
  assign n28833 = n28830 | n28831;
  assign n28834 = ~n28832 & n28833;
  assign n55017 = n28419 & n28834;
  assign n55018 = (n28834 & n54802) | (n28834 & n55017) | (n54802 & n55017);
  assign n55019 = n28419 | n28834;
  assign n55020 = n54802 | n55019;
  assign n28837 = ~n55018 & n55020;
  assign n28838 = x134 & x207;
  assign n28839 = n28837 & n28838;
  assign n28840 = n28837 | n28838;
  assign n28841 = ~n28839 & n28840;
  assign n55021 = n28426 & n28841;
  assign n55022 = (n28841 & n54806) | (n28841 & n55021) | (n54806 & n55021);
  assign n55023 = n28426 | n28841;
  assign n55024 = n54806 | n55023;
  assign n28844 = ~n55022 & n55024;
  assign n28845 = x133 & x208;
  assign n28846 = n28844 & n28845;
  assign n28847 = n28844 | n28845;
  assign n28848 = ~n28846 & n28847;
  assign n55025 = n28433 & n28848;
  assign n55026 = (n28848 & n54810) | (n28848 & n55025) | (n54810 & n55025);
  assign n55027 = n28433 | n28848;
  assign n55028 = n54810 | n55027;
  assign n28851 = ~n55026 & n55028;
  assign n28852 = x132 & x209;
  assign n28853 = n28851 & n28852;
  assign n28854 = n28851 | n28852;
  assign n28855 = ~n28853 & n28854;
  assign n55029 = n28440 & n28855;
  assign n55030 = (n28855 & n54814) | (n28855 & n55029) | (n54814 & n55029);
  assign n55031 = n28440 | n28855;
  assign n55032 = n54814 | n55031;
  assign n28858 = ~n55030 & n55032;
  assign n28859 = x131 & x210;
  assign n28860 = n28858 & n28859;
  assign n28861 = n28858 | n28859;
  assign n28862 = ~n28860 & n28861;
  assign n55033 = n28447 & n28862;
  assign n55034 = (n28862 & n54818) | (n28862 & n55033) | (n54818 & n55033);
  assign n55035 = n28447 | n28862;
  assign n55036 = n54818 | n55035;
  assign n28865 = ~n55034 & n55036;
  assign n28866 = x130 & x211;
  assign n28867 = n28865 & n28866;
  assign n28868 = n28865 | n28866;
  assign n28869 = ~n28867 & n28868;
  assign n55037 = n28454 & n28869;
  assign n55038 = (n28869 & n54823) | (n28869 & n55037) | (n54823 & n55037);
  assign n55039 = n28454 | n28869;
  assign n55040 = n54823 | n55039;
  assign n28872 = ~n55038 & n55040;
  assign n28873 = x129 & x212;
  assign n28874 = n28872 & n28873;
  assign n28875 = n28872 | n28873;
  assign n28876 = ~n28874 & n28875;
  assign n54857 = n28461 | n28463;
  assign n55041 = n28876 & n54857;
  assign n55042 = n28461 & n28876;
  assign n55043 = (n54654 & n55041) | (n54654 & n55042) | (n55041 & n55042);
  assign n55044 = n28876 | n54857;
  assign n55045 = n28461 | n28876;
  assign n55046 = (n54654 & n55044) | (n54654 & n55045) | (n55044 & n55045);
  assign n28879 = ~n55043 & n55046;
  assign n28880 = x128 & x213;
  assign n28881 = n28879 & n28880;
  assign n28882 = n28879 | n28880;
  assign n28883 = ~n28881 & n28882;
  assign n54855 = n28468 | n28470;
  assign n69539 = n28883 & n54855;
  assign n69540 = n28468 & n28883;
  assign n69541 = (n54652 & n69539) | (n54652 & n69540) | (n69539 & n69540);
  assign n69542 = n28883 | n54855;
  assign n69543 = n28468 | n28883;
  assign n69544 = (n54652 & n69542) | (n54652 & n69543) | (n69542 & n69543);
  assign n28886 = ~n69541 & n69544;
  assign n28887 = x127 & x214;
  assign n28888 = n28886 & n28887;
  assign n28889 = n28886 | n28887;
  assign n28890 = ~n28888 & n28889;
  assign n54853 = n28475 | n28477;
  assign n69545 = n28890 & n54853;
  assign n69546 = n28475 & n28890;
  assign n69547 = (n54650 & n69545) | (n54650 & n69546) | (n69545 & n69546);
  assign n69548 = n28890 | n54853;
  assign n69549 = n28475 | n28890;
  assign n69550 = (n54650 & n69548) | (n54650 & n69549) | (n69548 & n69549);
  assign n28893 = ~n69547 & n69550;
  assign n28894 = x126 & x215;
  assign n28895 = n28893 & n28894;
  assign n28896 = n28893 | n28894;
  assign n28897 = ~n28895 & n28896;
  assign n28898 = n54852 & n28897;
  assign n28899 = n54852 | n28897;
  assign n28900 = ~n28898 & n28899;
  assign n28901 = x125 & x216;
  assign n28902 = n28900 & n28901;
  assign n28903 = n28900 | n28901;
  assign n28904 = ~n28902 & n28903;
  assign n28905 = n54850 & n28904;
  assign n28906 = n54850 | n28904;
  assign n28907 = ~n28905 & n28906;
  assign n28908 = x124 & x217;
  assign n28909 = n28907 & n28908;
  assign n28910 = n28907 | n28908;
  assign n28911 = ~n28909 & n28910;
  assign n28912 = n54848 & n28911;
  assign n28913 = n54848 | n28911;
  assign n28914 = ~n28912 & n28913;
  assign n28915 = x123 & x218;
  assign n28916 = n28914 & n28915;
  assign n28917 = n28914 | n28915;
  assign n28918 = ~n28916 & n28917;
  assign n28919 = n54846 & n28918;
  assign n28920 = n54846 | n28918;
  assign n28921 = ~n28919 & n28920;
  assign n28922 = x122 & x219;
  assign n28923 = n28921 & n28922;
  assign n28924 = n28921 | n28922;
  assign n28925 = ~n28923 & n28924;
  assign n28926 = n54844 & n28925;
  assign n28927 = n54844 | n28925;
  assign n28928 = ~n28926 & n28927;
  assign n28929 = x121 & x220;
  assign n28930 = n28928 & n28929;
  assign n28931 = n28928 | n28929;
  assign n28932 = ~n28930 & n28931;
  assign n28933 = n54842 & n28932;
  assign n28934 = n54842 | n28932;
  assign n28935 = ~n28933 & n28934;
  assign n28936 = x120 & x221;
  assign n28937 = n28935 & n28936;
  assign n28938 = n28935 | n28936;
  assign n28939 = ~n28937 & n28938;
  assign n28940 = n54840 & n28939;
  assign n28941 = n54840 | n28939;
  assign n28942 = ~n28940 & n28941;
  assign n28943 = x119 & x222;
  assign n28944 = n28942 & n28943;
  assign n28945 = n28942 | n28943;
  assign n28946 = ~n28944 & n28945;
  assign n28947 = n54838 & n28946;
  assign n28948 = n54838 | n28946;
  assign n28949 = ~n28947 & n28948;
  assign n28950 = x118 & x223;
  assign n28951 = n28949 & n28950;
  assign n28952 = n28949 | n28950;
  assign n28953 = ~n28951 & n28952;
  assign n28954 = n54836 & n28953;
  assign n28955 = n54836 | n28953;
  assign n28956 = ~n28954 & n28955;
  assign n28957 = x117 & x224;
  assign n28958 = n28956 & n28957;
  assign n28959 = n28956 | n28957;
  assign n28960 = ~n28958 & n28959;
  assign n28961 = n54834 & n28960;
  assign n28962 = n54834 | n28960;
  assign n28963 = ~n28961 & n28962;
  assign n28964 = x116 & x225;
  assign n28965 = n28963 & n28964;
  assign n28966 = n28963 | n28964;
  assign n28967 = ~n28965 & n28966;
  assign n28968 = n54832 & n28967;
  assign n28969 = n54832 | n28967;
  assign n28970 = ~n28968 & n28969;
  assign n28971 = x115 & x226;
  assign n28972 = n28970 & n28971;
  assign n28973 = n28970 | n28971;
  assign n28974 = ~n28972 & n28973;
  assign n28975 = n54830 & n28974;
  assign n28976 = n54830 | n28974;
  assign n28977 = ~n28975 & n28976;
  assign n28978 = x114 & x227;
  assign n28979 = n28977 & n28978;
  assign n28980 = n28977 | n28978;
  assign n28981 = ~n28979 & n28980;
  assign n28982 = n54828 & n28981;
  assign n28983 = n54828 | n28981;
  assign n28984 = ~n28982 & n28983;
  assign n28985 = x113 & x228;
  assign n28986 = n28984 & n28985;
  assign n28987 = n28984 | n28985;
  assign n28988 = ~n28986 & n28987;
  assign n28989 = n28573 & n28988;
  assign n28990 = n28573 | n28988;
  assign n28991 = ~n28989 & n28990;
  assign n28992 = x112 & x229;
  assign n28993 = n28991 & n28992;
  assign n28994 = n28991 | n28992;
  assign n28995 = ~n28993 & n28994;
  assign n69551 = n28573 | n28985;
  assign n69552 = (n28573 & n28984) | (n28573 & n69551) | (n28984 & n69551);
  assign n55048 = (n28986 & n28988) | (n28986 & n69552) | (n28988 & n69552);
  assign n69553 = n28979 | n54828;
  assign n69554 = (n28979 & n28981) | (n28979 & n69553) | (n28981 & n69553);
  assign n28998 = n28972 | n28975;
  assign n28999 = n28965 | n28968;
  assign n29000 = n28958 | n28961;
  assign n29001 = n28951 | n28954;
  assign n29002 = n28944 | n28947;
  assign n29003 = n28937 | n28940;
  assign n29004 = n28930 | n28933;
  assign n29005 = n28923 | n28926;
  assign n55049 = n28916 | n28918;
  assign n55050 = (n28916 & n54846) | (n28916 & n55049) | (n54846 & n55049);
  assign n55051 = n28909 | n28911;
  assign n55052 = (n28909 & n54848) | (n28909 & n55051) | (n54848 & n55051);
  assign n55053 = n28902 | n28904;
  assign n55054 = (n28902 & n54850) | (n28902 & n55053) | (n54850 & n55053);
  assign n54854 = (n28475 & n54650) | (n28475 & n54853) | (n54650 & n54853);
  assign n54856 = (n28468 & n54652) | (n28468 & n54855) | (n54652 & n54855);
  assign n55067 = n28755 | n28757;
  assign n69557 = n28342 | n28755;
  assign n69558 = (n28755 & n28757) | (n28755 & n69557) | (n28757 & n69557);
  assign n69559 = (n54760 & n55067) | (n54760 & n69558) | (n55067 & n69558);
  assign n69560 = (n54759 & n55067) | (n54759 & n69558) | (n55067 & n69558);
  assign n69561 = (n69181 & n69559) | (n69181 & n69560) | (n69559 & n69560);
  assign n55072 = n28734 | n28736;
  assign n69562 = n28321 | n28734;
  assign n69563 = (n28734 & n28736) | (n28734 & n69562) | (n28736 & n69562);
  assign n69564 = (n54750 & n55072) | (n54750 & n69563) | (n55072 & n69563);
  assign n69565 = (n54749 & n55072) | (n54749 & n69563) | (n55072 & n69563);
  assign n69566 = (n69186 & n69564) | (n69186 & n69565) | (n69564 & n69565);
  assign n54873 = (n54545 & n69434) | (n54545 & n54872) | (n69434 & n54872);
  assign n55077 = n28713 | n28715;
  assign n69567 = n28300 | n28713;
  assign n69568 = (n28713 & n28715) | (n28713 & n69567) | (n28715 & n69567);
  assign n69569 = (n54740 & n55077) | (n54740 & n69568) | (n55077 & n69568);
  assign n69570 = (n54739 & n55077) | (n54739 & n69568) | (n55077 & n69568);
  assign n69571 = (n54460 & n69569) | (n54460 & n69570) | (n69569 & n69570);
  assign n54878 = (n54535 & n69436) | (n54535 & n54877) | (n69436 & n54877);
  assign n69572 = n28272 | n28685;
  assign n69573 = (n28685 & n28687) | (n28685 & n69572) | (n28687 & n69572);
  assign n69574 = n28685 | n28687;
  assign n69575 = (n28685 & n54882) | (n28685 & n69574) | (n54882 & n69574);
  assign n69576 = (n54678 & n69573) | (n54678 & n69575) | (n69573 & n69575);
  assign n69577 = (n69324 & n69573) | (n69324 & n69575) | (n69573 & n69575);
  assign n69578 = (n54276 & n69576) | (n54276 & n69577) | (n69576 & n69577);
  assign n29048 = x166 & x176;
  assign n29049 = x165 & x177;
  assign n29050 = n29048 & n29049;
  assign n29051 = n29048 | n29049;
  assign n29052 = ~n29050 & n29051;
  assign n69592 = n28629 & n29052;
  assign n69593 = (n29052 & n69446) | (n29052 & n69592) | (n69446 & n69592);
  assign n69594 = n28629 | n69447;
  assign n69597 = n29052 & n69594;
  assign n69595 = n28629 | n28631;
  assign n69598 = n29052 & n69595;
  assign n69599 = (n69340 & n69597) | (n69340 & n69598) | (n69597 & n69598);
  assign n69600 = (n53919 & n69593) | (n53919 & n69599) | (n69593 & n69599);
  assign n69601 = (n53918 & n69593) | (n53918 & n69599) | (n69593 & n69599);
  assign n69602 = (n68195 & n69600) | (n68195 & n69601) | (n69600 & n69601);
  assign n69603 = n28629 | n29052;
  assign n69604 = n69446 | n69603;
  assign n69605 = n29052 | n69594;
  assign n69606 = n29052 | n69595;
  assign n69607 = (n69340 & n69605) | (n69340 & n69606) | (n69605 & n69606);
  assign n69608 = (n53919 & n69604) | (n53919 & n69607) | (n69604 & n69607);
  assign n69609 = (n53918 & n69604) | (n53918 & n69607) | (n69604 & n69607);
  assign n69610 = (n68195 & n69608) | (n68195 & n69609) | (n69608 & n69609);
  assign n29055 = ~n69602 & n69610;
  assign n29056 = x164 & x178;
  assign n29057 = n29055 & n29056;
  assign n29058 = n29055 | n29056;
  assign n29059 = ~n29057 & n29058;
  assign n69611 = n28636 | n28638;
  assign n69612 = (n28636 & n69461) | (n28636 & n69611) | (n69461 & n69611);
  assign n55115 = n29059 & n69612;
  assign n69613 = (n28636 & n54898) | (n28636 & n69611) | (n54898 & n69611);
  assign n55116 = n29059 & n69613;
  assign n69614 = (n55115 & n55116) | (n55115 & n69221) | (n55116 & n69221);
  assign n69615 = (n55115 & n55116) | (n55115 & n69220) | (n55116 & n69220);
  assign n69616 = (n68389 & n69614) | (n68389 & n69615) | (n69614 & n69615);
  assign n55118 = n29059 | n69612;
  assign n55119 = n29059 | n69613;
  assign n69617 = (n55118 & n55119) | (n55118 & n69221) | (n55119 & n69221);
  assign n69618 = (n55118 & n55119) | (n55118 & n69220) | (n55119 & n69220);
  assign n69619 = (n68389 & n69617) | (n68389 & n69618) | (n69617 & n69618);
  assign n29062 = ~n69616 & n69619;
  assign n29063 = x163 & x179;
  assign n29064 = n29062 & n29063;
  assign n29065 = n29062 | n29063;
  assign n29066 = ~n29064 & n29065;
  assign n69586 = n28643 | n28645;
  assign n69587 = (n28643 & n69469) | (n28643 & n69586) | (n69469 & n69586);
  assign n69588 = (n28643 & n69470) | (n28643 & n69586) | (n69470 & n69586);
  assign n69590 = (n69108 & n69587) | (n69108 & n69588) | (n69587 & n69588);
  assign n69620 = n29066 & n69590;
  assign n69589 = (n54309 & n69587) | (n54309 & n69588) | (n69587 & n69588);
  assign n69621 = n29066 & n69589;
  assign n69622 = (n68776 & n69620) | (n68776 & n69621) | (n69620 & n69621);
  assign n69623 = n29066 | n69590;
  assign n69624 = n29066 | n69589;
  assign n69625 = (n68776 & n69623) | (n68776 & n69624) | (n69623 & n69624);
  assign n29069 = ~n69622 & n69625;
  assign n29070 = x162 & x180;
  assign n29071 = n29069 & n29070;
  assign n29072 = n29069 | n29070;
  assign n29073 = ~n29071 & n29072;
  assign n69626 = n28650 | n28652;
  assign n69627 = (n28650 & n54892) | (n28650 & n69626) | (n54892 & n69626);
  assign n55121 = n29073 & n69627;
  assign n69628 = n28237 | n28650;
  assign n69629 = (n28650 & n28652) | (n28650 & n69628) | (n28652 & n69628);
  assign n55122 = n29073 & n69629;
  assign n69630 = (n55121 & n55122) | (n55121 & n69333) | (n55122 & n69333);
  assign n69631 = (n55121 & n55122) | (n55121 & n69334) | (n55122 & n69334);
  assign n69632 = (n68982 & n69630) | (n68982 & n69631) | (n69630 & n69631);
  assign n55124 = n29073 | n69627;
  assign n55125 = n29073 | n69629;
  assign n69633 = (n55124 & n55125) | (n55124 & n69333) | (n55125 & n69333);
  assign n69634 = (n55124 & n55125) | (n55124 & n69334) | (n55125 & n69334);
  assign n69635 = (n68982 & n69633) | (n68982 & n69634) | (n69633 & n69634);
  assign n29076 = ~n69632 & n69635;
  assign n29077 = x161 & x181;
  assign n29078 = n29076 & n29077;
  assign n29079 = n29076 | n29077;
  assign n29080 = ~n29078 & n29079;
  assign n69636 = n28244 | n28657;
  assign n69637 = (n28657 & n28659) | (n28657 & n69636) | (n28659 & n69636);
  assign n55127 = n29080 & n69637;
  assign n55095 = n28657 | n28659;
  assign n55128 = n29080 & n55095;
  assign n69638 = (n54713 & n55127) | (n54713 & n55128) | (n55127 & n55128);
  assign n69639 = (n54714 & n55127) | (n54714 & n55128) | (n55127 & n55128);
  assign n69640 = (n69084 & n69638) | (n69084 & n69639) | (n69638 & n69639);
  assign n55130 = n29080 | n69637;
  assign n55131 = n29080 | n55095;
  assign n69641 = (n54713 & n55130) | (n54713 & n55131) | (n55130 & n55131);
  assign n69642 = (n54714 & n55130) | (n54714 & n55131) | (n55130 & n55131);
  assign n69643 = (n69084 & n69641) | (n69084 & n69642) | (n69641 & n69642);
  assign n29083 = ~n69640 & n69643;
  assign n29084 = x160 & x182;
  assign n29085 = n29083 & n29084;
  assign n29086 = n29083 | n29084;
  assign n29087 = ~n29085 & n29086;
  assign n69583 = n28664 | n28666;
  assign n69585 = (n28664 & n54890) | (n28664 & n69583) | (n54890 & n69583);
  assign n69644 = n29087 & n69585;
  assign n69584 = (n28664 & n69490) | (n28664 & n69583) | (n69490 & n69583);
  assign n69645 = n29087 & n69584;
  assign n69646 = (n69244 & n69644) | (n69244 & n69645) | (n69644 & n69645);
  assign n69647 = n29087 | n69585;
  assign n69648 = n29087 | n69584;
  assign n69649 = (n69244 & n69647) | (n69244 & n69648) | (n69647 & n69648);
  assign n29090 = ~n69646 & n69649;
  assign n29091 = x159 & x183;
  assign n29092 = n29090 & n29091;
  assign n29093 = n29090 | n29091;
  assign n29094 = ~n29092 & n29093;
  assign n69579 = n28671 | n28673;
  assign n69580 = (n28671 & n54887) | (n28671 & n69579) | (n54887 & n69579);
  assign n69650 = n29094 & n69580;
  assign n69581 = n28258 | n28671;
  assign n69582 = (n28671 & n28673) | (n28671 & n69581) | (n28673 & n69581);
  assign n69651 = n29094 & n69582;
  assign n69652 = (n69331 & n69650) | (n69331 & n69651) | (n69650 & n69651);
  assign n69653 = n29094 | n69580;
  assign n69654 = n29094 | n69582;
  assign n69655 = (n69331 & n69653) | (n69331 & n69654) | (n69653 & n69654);
  assign n29097 = ~n69652 & n69655;
  assign n29098 = x158 & x184;
  assign n29099 = n29097 & n29098;
  assign n29100 = n29097 | n29098;
  assign n29101 = ~n29099 & n29100;
  assign n55086 = n28678 | n28680;
  assign n55133 = n29101 & n55086;
  assign n55134 = n28678 & n29101;
  assign n69656 = (n54885 & n55133) | (n54885 & n55134) | (n55133 & n55134);
  assign n69657 = (n55133 & n55134) | (n55133 & n69440) | (n55134 & n69440);
  assign n69658 = (n69197 & n69656) | (n69197 & n69657) | (n69656 & n69657);
  assign n55136 = n29101 | n55086;
  assign n55137 = n28678 | n29101;
  assign n69659 = (n54885 & n55136) | (n54885 & n55137) | (n55136 & n55137);
  assign n69660 = (n55136 & n55137) | (n55136 & n69440) | (n55137 & n69440);
  assign n69661 = (n69197 & n69659) | (n69197 & n69660) | (n69659 & n69660);
  assign n29104 = ~n69658 & n69661;
  assign n29105 = x157 & x185;
  assign n29106 = n29104 & n29105;
  assign n29107 = n29104 | n29105;
  assign n29108 = ~n29106 & n29107;
  assign n29109 = n69578 & n29108;
  assign n29110 = n69578 | n29108;
  assign n29111 = ~n29109 & n29110;
  assign n29112 = x156 & x186;
  assign n29113 = n29111 & n29112;
  assign n29114 = n29111 | n29112;
  assign n29115 = ~n29113 & n29114;
  assign n55081 = n28692 | n28694;
  assign n55139 = n29115 & n55081;
  assign n55140 = n28692 & n29115;
  assign n69662 = (n54880 & n55139) | (n54880 & n55140) | (n55139 & n55140);
  assign n69663 = (n55139 & n55140) | (n55139 & n69438) | (n55140 & n69438);
  assign n69664 = (n54465 & n69662) | (n54465 & n69663) | (n69662 & n69663);
  assign n55142 = n29115 | n55081;
  assign n55143 = n28692 | n29115;
  assign n69665 = (n54880 & n55142) | (n54880 & n55143) | (n55142 & n55143);
  assign n69666 = (n55142 & n55143) | (n55142 & n69438) | (n55143 & n69438);
  assign n69667 = (n54465 & n69665) | (n54465 & n69666) | (n69665 & n69666);
  assign n29118 = ~n69664 & n69667;
  assign n29119 = x155 & x187;
  assign n29120 = n29118 & n29119;
  assign n29121 = n29118 | n29119;
  assign n29122 = ~n29120 & n29121;
  assign n55079 = n28699 | n28701;
  assign n55145 = n29122 & n55079;
  assign n55146 = n28699 & n29122;
  assign n55147 = (n54878 & n55145) | (n54878 & n55146) | (n55145 & n55146);
  assign n55148 = n29122 | n55079;
  assign n55149 = n28699 | n29122;
  assign n55150 = (n54878 & n55148) | (n54878 & n55149) | (n55148 & n55149);
  assign n29125 = ~n55147 & n55150;
  assign n29126 = x154 & x188;
  assign n29127 = n29125 & n29126;
  assign n29128 = n29125 | n29126;
  assign n29129 = ~n29127 & n29128;
  assign n55151 = n28706 & n29129;
  assign n55152 = (n29129 & n54951) | (n29129 & n55151) | (n54951 & n55151);
  assign n55153 = n28706 | n29129;
  assign n55154 = n54951 | n55153;
  assign n29132 = ~n55152 & n55154;
  assign n29133 = x153 & x189;
  assign n29134 = n29132 & n29133;
  assign n29135 = n29132 | n29133;
  assign n29136 = ~n29134 & n29135;
  assign n29137 = n69571 & n29136;
  assign n29138 = n69571 | n29136;
  assign n29139 = ~n29137 & n29138;
  assign n29140 = x152 & x190;
  assign n29141 = n29139 & n29140;
  assign n29142 = n29139 | n29140;
  assign n29143 = ~n29141 & n29142;
  assign n55074 = n28720 | n28722;
  assign n55155 = n29143 & n55074;
  assign n55156 = n28720 & n29143;
  assign n55157 = (n54873 & n55155) | (n54873 & n55156) | (n55155 & n55156);
  assign n55158 = n29143 | n55074;
  assign n55159 = n28720 | n29143;
  assign n55160 = (n54873 & n55158) | (n54873 & n55159) | (n55158 & n55159);
  assign n29146 = ~n55157 & n55160;
  assign n29147 = x151 & x191;
  assign n29148 = n29146 & n29147;
  assign n29149 = n29146 | n29147;
  assign n29150 = ~n29148 & n29149;
  assign n55161 = n28727 & n29150;
  assign n55162 = (n29150 & n54961) | (n29150 & n55161) | (n54961 & n55161);
  assign n55163 = n28727 | n29150;
  assign n55164 = n54961 | n55163;
  assign n29153 = ~n55162 & n55164;
  assign n29154 = x150 & x192;
  assign n29155 = n29153 & n29154;
  assign n29156 = n29153 | n29154;
  assign n29157 = ~n29155 & n29156;
  assign n29158 = n69566 & n29157;
  assign n29159 = n69566 | n29157;
  assign n29160 = ~n29158 & n29159;
  assign n29161 = x149 & x193;
  assign n29162 = n29160 & n29161;
  assign n29163 = n29160 | n29161;
  assign n29164 = ~n29162 & n29163;
  assign n55069 = n28741 | n28743;
  assign n55165 = n29164 & n55069;
  assign n55166 = n28741 & n29164;
  assign n55167 = (n69432 & n55165) | (n69432 & n55166) | (n55165 & n55166);
  assign n55168 = n29164 | n55069;
  assign n55169 = n28741 | n29164;
  assign n55170 = (n69432 & n55168) | (n69432 & n55169) | (n55168 & n55169);
  assign n29167 = ~n55167 & n55170;
  assign n29168 = x148 & x194;
  assign n29169 = n29167 & n29168;
  assign n29170 = n29167 | n29168;
  assign n29171 = ~n29169 & n29170;
  assign n55171 = n28748 & n29171;
  assign n69668 = (n29171 & n54970) | (n29171 & n55171) | (n54970 & n55171);
  assign n69669 = (n29171 & n54969) | (n29171 & n55171) | (n54969 & n55171);
  assign n69670 = (n69312 & n69668) | (n69312 & n69669) | (n69668 & n69669);
  assign n55173 = n28748 | n29171;
  assign n69671 = n54970 | n55173;
  assign n69672 = n54969 | n55173;
  assign n69673 = (n69312 & n69671) | (n69312 & n69672) | (n69671 & n69672);
  assign n29174 = ~n69670 & n69673;
  assign n29175 = x147 & x195;
  assign n29176 = n29174 & n29175;
  assign n29177 = n29174 | n29175;
  assign n29178 = ~n29176 & n29177;
  assign n29179 = n69561 & n29178;
  assign n29180 = n69561 | n29178;
  assign n29181 = ~n29179 & n29180;
  assign n29182 = x146 & x196;
  assign n29183 = n29181 & n29182;
  assign n29184 = n29181 | n29182;
  assign n29185 = ~n29183 & n29184;
  assign n55064 = n28762 | n28764;
  assign n55175 = n29185 & n55064;
  assign n55176 = n28762 & n29185;
  assign n55177 = (n69427 & n55175) | (n69427 & n55176) | (n55175 & n55176);
  assign n55178 = n29185 | n55064;
  assign n55179 = n28762 | n29185;
  assign n55180 = (n69427 & n55178) | (n69427 & n55179) | (n55178 & n55179);
  assign n29188 = ~n55177 & n55180;
  assign n29189 = x145 & x197;
  assign n29190 = n29188 & n29189;
  assign n29191 = n29188 | n29189;
  assign n29192 = ~n29190 & n29191;
  assign n55181 = n28769 & n29192;
  assign n69674 = (n29192 & n54980) | (n29192 & n55181) | (n54980 & n55181);
  assign n69675 = (n29192 & n54979) | (n29192 & n55181) | (n54979 & n55181);
  assign n69676 = (n54659 & n69674) | (n54659 & n69675) | (n69674 & n69675);
  assign n55183 = n28769 | n29192;
  assign n69677 = n54980 | n55183;
  assign n69678 = n54979 | n55183;
  assign n69679 = (n54659 & n69677) | (n54659 & n69678) | (n69677 & n69678);
  assign n29195 = ~n69676 & n69679;
  assign n29196 = x144 & x198;
  assign n29197 = n29195 & n29196;
  assign n29198 = n29195 | n29196;
  assign n29199 = ~n29197 & n29198;
  assign n55062 = n28776 | n28778;
  assign n69680 = n29199 & n55062;
  assign n69555 = n28363 | n28776;
  assign n69556 = (n28776 & n28778) | (n28776 & n69555) | (n28778 & n69555);
  assign n69681 = n29199 & n69556;
  assign n69682 = (n69407 & n69680) | (n69407 & n69681) | (n69680 & n69681);
  assign n69683 = n29199 | n55062;
  assign n69684 = n29199 | n69556;
  assign n69685 = (n69407 & n69683) | (n69407 & n69684) | (n69683 & n69684);
  assign n29202 = ~n69682 & n69685;
  assign n29203 = x143 & x199;
  assign n29204 = n29202 & n29203;
  assign n29205 = n29202 | n29203;
  assign n29206 = ~n29204 & n29205;
  assign n55185 = n28783 & n29206;
  assign n69686 = (n29206 & n54989) | (n29206 & n55185) | (n54989 & n55185);
  assign n69687 = (n28785 & n29206) | (n28785 & n55185) | (n29206 & n55185);
  assign n69688 = (n54774 & n69686) | (n54774 & n69687) | (n69686 & n69687);
  assign n55187 = n28783 | n29206;
  assign n69689 = n54989 | n55187;
  assign n69690 = n28785 | n55187;
  assign n69691 = (n54774 & n69689) | (n54774 & n69690) | (n69689 & n69690);
  assign n29209 = ~n69688 & n69691;
  assign n29210 = x142 & x200;
  assign n29211 = n29209 & n29210;
  assign n29212 = n29209 | n29210;
  assign n29213 = ~n29211 & n29212;
  assign n55189 = n28790 & n29213;
  assign n55190 = (n29213 & n54994) | (n29213 & n55189) | (n54994 & n55189);
  assign n55191 = n28790 | n29213;
  assign n55192 = n54994 | n55191;
  assign n29216 = ~n55190 & n55192;
  assign n29217 = x141 & x201;
  assign n29218 = n29216 & n29217;
  assign n29219 = n29216 | n29217;
  assign n29220 = ~n29218 & n29219;
  assign n55193 = n28797 & n29220;
  assign n55194 = (n29220 & n54998) | (n29220 & n55193) | (n54998 & n55193);
  assign n55195 = n28797 | n29220;
  assign n55196 = n54998 | n55195;
  assign n29223 = ~n55194 & n55196;
  assign n29224 = x140 & x202;
  assign n29225 = n29223 & n29224;
  assign n29226 = n29223 | n29224;
  assign n29227 = ~n29225 & n29226;
  assign n55197 = n28804 & n29227;
  assign n55198 = (n29227 & n55002) | (n29227 & n55197) | (n55002 & n55197);
  assign n55199 = n28804 | n29227;
  assign n55200 = n55002 | n55199;
  assign n29230 = ~n55198 & n55200;
  assign n29231 = x139 & x203;
  assign n29232 = n29230 & n29231;
  assign n29233 = n29230 | n29231;
  assign n29234 = ~n29232 & n29233;
  assign n55201 = n28811 & n29234;
  assign n55202 = (n29234 & n55006) | (n29234 & n55201) | (n55006 & n55201);
  assign n55203 = n28811 | n29234;
  assign n55204 = n55006 | n55203;
  assign n29237 = ~n55202 & n55204;
  assign n29238 = x138 & x204;
  assign n29239 = n29237 & n29238;
  assign n29240 = n29237 | n29238;
  assign n29241 = ~n29239 & n29240;
  assign n55205 = n28818 & n29241;
  assign n55206 = (n29241 & n55010) | (n29241 & n55205) | (n55010 & n55205);
  assign n55207 = n28818 | n29241;
  assign n55208 = n55010 | n55207;
  assign n29244 = ~n55206 & n55208;
  assign n29245 = x137 & x205;
  assign n29246 = n29244 & n29245;
  assign n29247 = n29244 | n29245;
  assign n29248 = ~n29246 & n29247;
  assign n55209 = n28825 & n29248;
  assign n55210 = (n29248 & n55014) | (n29248 & n55209) | (n55014 & n55209);
  assign n55211 = n28825 | n29248;
  assign n55212 = n55014 | n55211;
  assign n29251 = ~n55210 & n55212;
  assign n29252 = x136 & x206;
  assign n29253 = n29251 & n29252;
  assign n29254 = n29251 | n29252;
  assign n29255 = ~n29253 & n29254;
  assign n55213 = n28832 & n29255;
  assign n55214 = (n29255 & n55018) | (n29255 & n55213) | (n55018 & n55213);
  assign n55215 = n28832 | n29255;
  assign n55216 = n55018 | n55215;
  assign n29258 = ~n55214 & n55216;
  assign n29259 = x135 & x207;
  assign n29260 = n29258 & n29259;
  assign n29261 = n29258 | n29259;
  assign n29262 = ~n29260 & n29261;
  assign n55217 = n28839 & n29262;
  assign n55218 = (n29262 & n55022) | (n29262 & n55217) | (n55022 & n55217);
  assign n55219 = n28839 | n29262;
  assign n55220 = n55022 | n55219;
  assign n29265 = ~n55218 & n55220;
  assign n29266 = x134 & x208;
  assign n29267 = n29265 & n29266;
  assign n29268 = n29265 | n29266;
  assign n29269 = ~n29267 & n29268;
  assign n55221 = n28846 & n29269;
  assign n55222 = (n29269 & n55026) | (n29269 & n55221) | (n55026 & n55221);
  assign n55223 = n28846 | n29269;
  assign n55224 = n55026 | n55223;
  assign n29272 = ~n55222 & n55224;
  assign n29273 = x133 & x209;
  assign n29274 = n29272 & n29273;
  assign n29275 = n29272 | n29273;
  assign n29276 = ~n29274 & n29275;
  assign n55225 = n28853 & n29276;
  assign n55226 = (n29276 & n55030) | (n29276 & n55225) | (n55030 & n55225);
  assign n55227 = n28853 | n29276;
  assign n55228 = n55030 | n55227;
  assign n29279 = ~n55226 & n55228;
  assign n29280 = x132 & x210;
  assign n29281 = n29279 & n29280;
  assign n29282 = n29279 | n29280;
  assign n29283 = ~n29281 & n29282;
  assign n55229 = n28860 & n29283;
  assign n55230 = (n29283 & n55034) | (n29283 & n55229) | (n55034 & n55229);
  assign n55231 = n28860 | n29283;
  assign n55232 = n55034 | n55231;
  assign n29286 = ~n55230 & n55232;
  assign n29287 = x131 & x211;
  assign n29288 = n29286 & n29287;
  assign n29289 = n29286 | n29287;
  assign n29290 = ~n29288 & n29289;
  assign n55233 = n28867 & n29290;
  assign n55234 = (n29290 & n55038) | (n29290 & n55233) | (n55038 & n55233);
  assign n55235 = n28867 | n29290;
  assign n55236 = n55038 | n55235;
  assign n29293 = ~n55234 & n55236;
  assign n29294 = x130 & x212;
  assign n29295 = n29293 & n29294;
  assign n29296 = n29293 | n29294;
  assign n29297 = ~n29295 & n29296;
  assign n55237 = n28874 & n29297;
  assign n55238 = (n29297 & n55043) | (n29297 & n55237) | (n55043 & n55237);
  assign n55239 = n28874 | n29297;
  assign n55240 = n55043 | n55239;
  assign n29300 = ~n55238 & n55240;
  assign n29301 = x129 & x213;
  assign n29302 = n29300 & n29301;
  assign n29303 = n29300 | n29301;
  assign n29304 = ~n29302 & n29303;
  assign n55059 = n28881 | n28883;
  assign n55241 = n29304 & n55059;
  assign n55242 = n28881 & n29304;
  assign n55243 = (n54856 & n55241) | (n54856 & n55242) | (n55241 & n55242);
  assign n55244 = n29304 | n55059;
  assign n55245 = n28881 | n29304;
  assign n55246 = (n54856 & n55244) | (n54856 & n55245) | (n55244 & n55245);
  assign n29307 = ~n55243 & n55246;
  assign n29308 = x128 & x214;
  assign n29309 = n29307 & n29308;
  assign n29310 = n29307 | n29308;
  assign n29311 = ~n29309 & n29310;
  assign n55057 = n28888 | n28890;
  assign n69692 = n29311 & n55057;
  assign n69693 = n28888 & n29311;
  assign n69694 = (n54854 & n69692) | (n54854 & n69693) | (n69692 & n69693);
  assign n69695 = n29311 | n55057;
  assign n69696 = n28888 | n29311;
  assign n69697 = (n54854 & n69695) | (n54854 & n69696) | (n69695 & n69696);
  assign n29314 = ~n69694 & n69697;
  assign n29315 = x127 & x215;
  assign n29316 = n29314 & n29315;
  assign n29317 = n29314 | n29315;
  assign n29318 = ~n29316 & n29317;
  assign n55055 = n28895 | n28897;
  assign n69698 = n29318 & n55055;
  assign n69699 = n28895 & n29318;
  assign n69700 = (n54852 & n69698) | (n54852 & n69699) | (n69698 & n69699);
  assign n69701 = n29318 | n55055;
  assign n69702 = n28895 | n29318;
  assign n69703 = (n54852 & n69701) | (n54852 & n69702) | (n69701 & n69702);
  assign n29321 = ~n69700 & n69703;
  assign n29322 = x126 & x216;
  assign n29323 = n29321 & n29322;
  assign n29324 = n29321 | n29322;
  assign n29325 = ~n29323 & n29324;
  assign n29326 = n55054 & n29325;
  assign n29327 = n55054 | n29325;
  assign n29328 = ~n29326 & n29327;
  assign n29329 = x125 & x217;
  assign n29330 = n29328 & n29329;
  assign n29331 = n29328 | n29329;
  assign n29332 = ~n29330 & n29331;
  assign n29333 = n55052 & n29332;
  assign n29334 = n55052 | n29332;
  assign n29335 = ~n29333 & n29334;
  assign n29336 = x124 & x218;
  assign n29337 = n29335 & n29336;
  assign n29338 = n29335 | n29336;
  assign n29339 = ~n29337 & n29338;
  assign n29340 = n55050 & n29339;
  assign n29341 = n55050 | n29339;
  assign n29342 = ~n29340 & n29341;
  assign n29343 = x123 & x219;
  assign n29344 = n29342 & n29343;
  assign n29345 = n29342 | n29343;
  assign n29346 = ~n29344 & n29345;
  assign n29347 = n29005 & n29346;
  assign n29348 = n29005 | n29346;
  assign n29349 = ~n29347 & n29348;
  assign n29350 = x122 & x220;
  assign n29351 = n29349 & n29350;
  assign n29352 = n29349 | n29350;
  assign n29353 = ~n29351 & n29352;
  assign n29354 = n29004 & n29353;
  assign n29355 = n29004 | n29353;
  assign n29356 = ~n29354 & n29355;
  assign n29357 = x121 & x221;
  assign n29358 = n29356 & n29357;
  assign n29359 = n29356 | n29357;
  assign n29360 = ~n29358 & n29359;
  assign n29361 = n29003 & n29360;
  assign n29362 = n29003 | n29360;
  assign n29363 = ~n29361 & n29362;
  assign n29364 = x120 & x222;
  assign n29365 = n29363 & n29364;
  assign n29366 = n29363 | n29364;
  assign n29367 = ~n29365 & n29366;
  assign n29368 = n29002 & n29367;
  assign n29369 = n29002 | n29367;
  assign n29370 = ~n29368 & n29369;
  assign n29371 = x119 & x223;
  assign n29372 = n29370 & n29371;
  assign n29373 = n29370 | n29371;
  assign n29374 = ~n29372 & n29373;
  assign n29375 = n29001 & n29374;
  assign n29376 = n29001 | n29374;
  assign n29377 = ~n29375 & n29376;
  assign n29378 = x118 & x224;
  assign n29379 = n29377 & n29378;
  assign n29380 = n29377 | n29378;
  assign n29381 = ~n29379 & n29380;
  assign n29382 = n29000 & n29381;
  assign n29383 = n29000 | n29381;
  assign n29384 = ~n29382 & n29383;
  assign n29385 = x117 & x225;
  assign n29386 = n29384 & n29385;
  assign n29387 = n29384 | n29385;
  assign n29388 = ~n29386 & n29387;
  assign n29389 = n28999 & n29388;
  assign n29390 = n28999 | n29388;
  assign n29391 = ~n29389 & n29390;
  assign n29392 = x116 & x226;
  assign n29393 = n29391 & n29392;
  assign n29394 = n29391 | n29392;
  assign n29395 = ~n29393 & n29394;
  assign n29396 = n28998 & n29395;
  assign n29397 = n28998 | n29395;
  assign n29398 = ~n29396 & n29397;
  assign n29399 = x115 & x227;
  assign n29400 = n29398 & n29399;
  assign n29401 = n29398 | n29399;
  assign n29402 = ~n29400 & n29401;
  assign n29403 = n69554 & n29402;
  assign n29404 = n69554 | n29402;
  assign n29405 = ~n29403 & n29404;
  assign n29406 = x114 & x228;
  assign n29407 = n29405 & n29406;
  assign n29408 = n29405 | n29406;
  assign n29409 = ~n29407 & n29408;
  assign n29410 = n55048 & n29409;
  assign n29411 = n55048 | n29409;
  assign n29412 = ~n29410 & n29411;
  assign n29413 = x113 & x229;
  assign n29414 = n29412 & n29413;
  assign n29415 = n29412 | n29413;
  assign n29416 = ~n29414 & n29415;
  assign n29417 = n28993 & n29416;
  assign n29418 = n28993 | n29416;
  assign n29419 = ~n29417 & n29418;
  assign n29420 = x112 & x230;
  assign n29421 = n29419 & n29420;
  assign n29422 = n29419 | n29420;
  assign n29423 = ~n29421 & n29422;
  assign n69704 = n28993 | n29413;
  assign n69705 = (n28993 & n29412) | (n28993 & n69704) | (n29412 & n69704);
  assign n55248 = (n29414 & n29416) | (n29414 & n69705) | (n29416 & n69705);
  assign n55249 = n29407 | n55048;
  assign n55250 = (n29407 & n29409) | (n29407 & n55249) | (n29409 & n55249);
  assign n69706 = n29400 | n69554;
  assign n69707 = (n29400 & n29402) | (n29400 & n69706) | (n29402 & n69706);
  assign n29427 = n29393 | n29396;
  assign n29428 = n29386 | n29389;
  assign n29429 = n29379 | n29382;
  assign n29430 = n29372 | n29375;
  assign n29431 = n29365 | n29368;
  assign n29432 = n29358 | n29361;
  assign n29433 = n29351 | n29354;
  assign n55251 = n29344 | n29346;
  assign n55252 = (n29005 & n29344) | (n29005 & n55251) | (n29344 & n55251);
  assign n55253 = n29337 | n29339;
  assign n55254 = (n29337 & n55050) | (n29337 & n55253) | (n55050 & n55253);
  assign n55255 = n29330 | n29332;
  assign n55256 = (n29330 & n55052) | (n29330 & n55255) | (n55052 & n55255);
  assign n55056 = (n28895 & n54852) | (n28895 & n55055) | (n54852 & n55055);
  assign n55058 = (n28888 & n54854) | (n28888 & n55057) | (n54854 & n55057);
  assign n55063 = (n69407 & n69556) | (n69407 & n55062) | (n69556 & n55062);
  assign n55266 = n29190 | n29192;
  assign n69708 = n28769 | n29190;
  assign n69709 = (n29190 & n29192) | (n29190 & n69708) | (n29192 & n69708);
  assign n69710 = (n54980 & n55266) | (n54980 & n69709) | (n55266 & n69709);
  assign n69711 = (n54979 & n55266) | (n54979 & n69709) | (n55266 & n69709);
  assign n69712 = (n54659 & n69710) | (n54659 & n69711) | (n69710 & n69711);
  assign n55271 = n29169 | n29171;
  assign n69713 = n28748 | n29169;
  assign n69714 = (n29169 & n29171) | (n29169 & n69713) | (n29171 & n69713);
  assign n69715 = (n54970 & n55271) | (n54970 & n69714) | (n55271 & n69714);
  assign n69716 = (n54969 & n55271) | (n54969 & n69714) | (n55271 & n69714);
  assign n69717 = (n69312 & n69715) | (n69312 & n69716) | (n69715 & n69716);
  assign n54881 = (n54465 & n69438) | (n54465 & n54880) | (n69438 & n54880);
  assign n69724 = n28678 | n29099;
  assign n69725 = (n29099 & n29101) | (n29099 & n69724) | (n29101 & n69724);
  assign n69726 = n29099 | n29101;
  assign n69727 = (n29099 & n55086) | (n29099 & n69726) | (n55086 & n69726);
  assign n69728 = (n54885 & n69725) | (n54885 & n69727) | (n69725 & n69727);
  assign n69729 = (n69440 & n69725) | (n69440 & n69727) | (n69725 & n69727);
  assign n69730 = (n69197 & n69728) | (n69197 & n69729) | (n69728 & n69729);
  assign n69731 = n29078 | n29080;
  assign n69732 = (n29078 & n69637) | (n29078 & n69731) | (n69637 & n69731);
  assign n69733 = (n29078 & n55095) | (n29078 & n69731) | (n55095 & n69731);
  assign n69734 = (n54713 & n69732) | (n54713 & n69733) | (n69732 & n69733);
  assign n69735 = (n54714 & n69732) | (n54714 & n69733) | (n69732 & n69733);
  assign n69736 = (n69084 & n69734) | (n69084 & n69735) | (n69734 & n69735);
  assign n29477 = x167 & x176;
  assign n29478 = x166 & x177;
  assign n29479 = n29477 & n29478;
  assign n29480 = n29477 | n29478;
  assign n29481 = ~n29479 & n29480;
  assign n55307 = n29050 | n69599;
  assign n69743 = n29050 | n69592;
  assign n69744 = n29050 | n29052;
  assign n69745 = (n69446 & n69743) | (n69446 & n69744) | (n69743 & n69744);
  assign n69747 = (n53918 & n55307) | (n53918 & n69745) | (n55307 & n69745);
  assign n69749 = n29481 & n69747;
  assign n69746 = (n53919 & n55307) | (n53919 & n69745) | (n55307 & n69745);
  assign n69750 = n29481 & n69746;
  assign n69751 = (n68195 & n69749) | (n68195 & n69750) | (n69749 & n69750);
  assign n69752 = n29481 | n69747;
  assign n69753 = n29481 | n69746;
  assign n69754 = (n68195 & n69752) | (n68195 & n69753) | (n69752 & n69753);
  assign n29484 = ~n69751 & n69754;
  assign n29485 = x165 & x178;
  assign n29486 = n29484 & n29485;
  assign n29487 = n29484 | n29485;
  assign n29488 = ~n29486 & n29487;
  assign n69755 = n29057 | n29059;
  assign n69757 = n29488 & n69755;
  assign n69758 = n29057 & n29488;
  assign n69759 = (n69612 & n69757) | (n69612 & n69758) | (n69757 & n69758);
  assign n69761 = (n69613 & n69757) | (n69613 & n69758) | (n69757 & n69758);
  assign n69762 = (n69221 & n69759) | (n69221 & n69761) | (n69759 & n69761);
  assign n69763 = (n69220 & n69759) | (n69220 & n69761) | (n69759 & n69761);
  assign n69764 = (n68389 & n69762) | (n68389 & n69763) | (n69762 & n69763);
  assign n69765 = n29488 | n69755;
  assign n69766 = n29057 | n29488;
  assign n69767 = (n69612 & n69765) | (n69612 & n69766) | (n69765 & n69766);
  assign n69768 = (n69613 & n69765) | (n69613 & n69766) | (n69765 & n69766);
  assign n69769 = (n69221 & n69767) | (n69221 & n69768) | (n69767 & n69768);
  assign n69770 = (n69220 & n69767) | (n69220 & n69768) | (n69767 & n69768);
  assign n69771 = (n68389 & n69769) | (n68389 & n69770) | (n69769 & n69770);
  assign n29491 = ~n69764 & n69771;
  assign n29492 = x164 & x179;
  assign n29493 = n29491 & n29492;
  assign n29494 = n29491 | n29492;
  assign n29495 = ~n29493 & n29494;
  assign n55301 = n29064 | n29066;
  assign n55315 = n29495 & n55301;
  assign n55316 = n29064 & n29495;
  assign n69772 = (n55315 & n55316) | (n55315 & n69590) | (n55316 & n69590);
  assign n69773 = (n55315 & n55316) | (n55315 & n69589) | (n55316 & n69589);
  assign n69774 = (n68776 & n69772) | (n68776 & n69773) | (n69772 & n69773);
  assign n55318 = n29495 | n55301;
  assign n55319 = n29064 | n29495;
  assign n69775 = (n55318 & n55319) | (n55318 & n69590) | (n55319 & n69590);
  assign n69776 = (n55318 & n55319) | (n55318 & n69589) | (n55319 & n69589);
  assign n69777 = (n68776 & n69775) | (n68776 & n69776) | (n69775 & n69776);
  assign n29498 = ~n69774 & n69777;
  assign n29499 = x163 & x180;
  assign n29500 = n29498 & n29499;
  assign n29501 = n29498 | n29499;
  assign n29502 = ~n29500 & n29501;
  assign n69737 = n29071 | n29073;
  assign n69738 = (n29071 & n69627) | (n29071 & n69737) | (n69627 & n69737);
  assign n69739 = (n29071 & n69629) | (n29071 & n69737) | (n69629 & n69737);
  assign n69741 = (n69334 & n69738) | (n69334 & n69739) | (n69738 & n69739);
  assign n69778 = n29502 & n69741;
  assign n69740 = (n69333 & n69738) | (n69333 & n69739) | (n69738 & n69739);
  assign n69779 = n29502 & n69740;
  assign n69780 = (n68982 & n69778) | (n68982 & n69779) | (n69778 & n69779);
  assign n69781 = n29502 | n69741;
  assign n69782 = n29502 | n69740;
  assign n69783 = (n68982 & n69781) | (n68982 & n69782) | (n69781 & n69782);
  assign n29505 = ~n69780 & n69783;
  assign n29506 = x162 & x181;
  assign n29507 = n29505 & n29506;
  assign n29508 = n29505 | n29506;
  assign n29509 = ~n29507 & n29508;
  assign n29510 = n69736 & n29509;
  assign n29511 = n69736 | n29509;
  assign n29512 = ~n29510 & n29511;
  assign n29513 = x161 & x182;
  assign n29514 = n29512 & n29513;
  assign n29515 = n29512 | n29513;
  assign n29516 = ~n29514 & n29515;
  assign n55293 = n29085 | n29087;
  assign n55321 = n29516 & n55293;
  assign n55322 = n29085 & n29516;
  assign n69784 = (n55321 & n55322) | (n55321 & n69585) | (n55322 & n69585);
  assign n69785 = (n55321 & n55322) | (n55321 & n69584) | (n55322 & n69584);
  assign n69786 = (n69244 & n69784) | (n69244 & n69785) | (n69784 & n69785);
  assign n55324 = n29516 | n55293;
  assign n55325 = n29085 | n29516;
  assign n69787 = (n55324 & n55325) | (n55324 & n69585) | (n55325 & n69585);
  assign n69788 = (n55324 & n55325) | (n55324 & n69584) | (n55325 & n69584);
  assign n69789 = (n69244 & n69787) | (n69244 & n69788) | (n69787 & n69788);
  assign n29519 = ~n69786 & n69789;
  assign n29520 = x160 & x183;
  assign n29521 = n29519 & n29520;
  assign n29522 = n29519 | n29520;
  assign n29523 = ~n29521 & n29522;
  assign n55291 = n29092 | n29094;
  assign n55327 = n29523 & n55291;
  assign n55328 = n29092 & n29523;
  assign n69790 = (n55327 & n55328) | (n55327 & n69580) | (n55328 & n69580);
  assign n69791 = (n55327 & n55328) | (n55327 & n69582) | (n55328 & n69582);
  assign n69792 = (n69331 & n69790) | (n69331 & n69791) | (n69790 & n69791);
  assign n55330 = n29523 | n55291;
  assign n55331 = n29092 | n29523;
  assign n69793 = (n55330 & n55331) | (n55330 & n69580) | (n55331 & n69580);
  assign n69794 = (n55330 & n55331) | (n55330 & n69582) | (n55331 & n69582);
  assign n69795 = (n69331 & n69793) | (n69331 & n69794) | (n69793 & n69794);
  assign n29526 = ~n69792 & n69795;
  assign n29527 = x159 & x184;
  assign n29528 = n29526 & n29527;
  assign n29529 = n29526 | n29527;
  assign n29530 = ~n29528 & n29529;
  assign n29531 = n69730 & n29530;
  assign n29532 = n69730 | n29530;
  assign n29533 = ~n29531 & n29532;
  assign n29534 = x158 & x185;
  assign n29535 = n29533 & n29534;
  assign n29536 = n29533 | n29534;
  assign n29537 = ~n29535 & n29536;
  assign n55286 = n29106 | n29108;
  assign n55333 = n29537 & n55286;
  assign n55334 = n29106 & n29537;
  assign n55335 = (n69578 & n55333) | (n69578 & n55334) | (n55333 & n55334);
  assign n55336 = n29537 | n55286;
  assign n55337 = n29106 | n29537;
  assign n55338 = (n69578 & n55336) | (n69578 & n55337) | (n55336 & n55337);
  assign n29540 = ~n55335 & n55338;
  assign n29541 = x157 & x186;
  assign n29542 = n29540 & n29541;
  assign n29543 = n29540 | n29541;
  assign n29544 = ~n29542 & n29543;
  assign n55284 = n29113 | n55139;
  assign n69796 = n29544 & n55284;
  assign n69722 = n28692 | n29113;
  assign n69723 = (n29113 & n29115) | (n29113 & n69722) | (n29115 & n69722);
  assign n69797 = n29544 & n69723;
  assign n69798 = (n54881 & n69796) | (n54881 & n69797) | (n69796 & n69797);
  assign n69799 = n29544 | n55284;
  assign n69800 = n29544 | n69723;
  assign n69801 = (n54881 & n69799) | (n54881 & n69800) | (n69799 & n69800);
  assign n29547 = ~n69798 & n69801;
  assign n29548 = x156 & x187;
  assign n29549 = n29547 & n29548;
  assign n29550 = n29547 | n29548;
  assign n29551 = ~n29549 & n29550;
  assign n55339 = n29120 & n29551;
  assign n69802 = (n29551 & n55145) | (n29551 & n55339) | (n55145 & n55339);
  assign n69803 = (n29551 & n55146) | (n29551 & n55339) | (n55146 & n55339);
  assign n69804 = (n54878 & n69802) | (n54878 & n69803) | (n69802 & n69803);
  assign n55341 = n29120 | n29551;
  assign n69805 = n55145 | n55341;
  assign n69806 = n55146 | n55341;
  assign n69807 = (n54878 & n69805) | (n54878 & n69806) | (n69805 & n69806);
  assign n29554 = ~n69804 & n69807;
  assign n29555 = x155 & x188;
  assign n29556 = n29554 & n29555;
  assign n29557 = n29554 | n29555;
  assign n29558 = ~n29556 & n29557;
  assign n55281 = n29127 | n29129;
  assign n69808 = n29558 & n55281;
  assign n69720 = n28706 | n29127;
  assign n69721 = (n29127 & n29129) | (n29127 & n69720) | (n29129 & n69720);
  assign n69809 = n29558 & n69721;
  assign n69810 = (n54951 & n69808) | (n54951 & n69809) | (n69808 & n69809);
  assign n69811 = n29558 | n55281;
  assign n69812 = n29558 | n69721;
  assign n69813 = (n54951 & n69811) | (n54951 & n69812) | (n69811 & n69812);
  assign n29561 = ~n69810 & n69813;
  assign n29562 = x154 & x189;
  assign n29563 = n29561 & n29562;
  assign n29564 = n29561 | n29562;
  assign n29565 = ~n29563 & n29564;
  assign n55278 = n29134 | n29136;
  assign n55343 = n29565 & n55278;
  assign n55344 = n29134 & n29565;
  assign n55345 = (n69571 & n55343) | (n69571 & n55344) | (n55343 & n55344);
  assign n55346 = n29565 | n55278;
  assign n55347 = n29134 | n29565;
  assign n55348 = (n69571 & n55346) | (n69571 & n55347) | (n55346 & n55347);
  assign n29568 = ~n55345 & n55348;
  assign n29569 = x153 & x190;
  assign n29570 = n29568 & n29569;
  assign n29571 = n29568 | n29569;
  assign n29572 = ~n29570 & n29571;
  assign n55349 = n29141 & n29572;
  assign n69814 = (n29572 & n55156) | (n29572 & n55349) | (n55156 & n55349);
  assign n69815 = (n29572 & n55155) | (n29572 & n55349) | (n55155 & n55349);
  assign n69816 = (n54873 & n69814) | (n54873 & n69815) | (n69814 & n69815);
  assign n55351 = n29141 | n29572;
  assign n69817 = n55156 | n55351;
  assign n69818 = n55155 | n55351;
  assign n69819 = (n54873 & n69817) | (n54873 & n69818) | (n69817 & n69818);
  assign n29575 = ~n69816 & n69819;
  assign n29576 = x152 & x191;
  assign n29577 = n29575 & n29576;
  assign n29578 = n29575 | n29576;
  assign n29579 = ~n29577 & n29578;
  assign n55276 = n29148 | n29150;
  assign n69820 = n29579 & n55276;
  assign n69718 = n28727 | n29148;
  assign n69719 = (n29148 & n29150) | (n29148 & n69718) | (n29150 & n69718);
  assign n69821 = n29579 & n69719;
  assign n69822 = (n54961 & n69820) | (n54961 & n69821) | (n69820 & n69821);
  assign n69823 = n29579 | n55276;
  assign n69824 = n29579 | n69719;
  assign n69825 = (n54961 & n69823) | (n54961 & n69824) | (n69823 & n69824);
  assign n29582 = ~n69822 & n69825;
  assign n29583 = x151 & x192;
  assign n29584 = n29582 & n29583;
  assign n29585 = n29582 | n29583;
  assign n29586 = ~n29584 & n29585;
  assign n55273 = n29155 | n29157;
  assign n55353 = n29586 & n55273;
  assign n55354 = n29155 & n29586;
  assign n55355 = (n69566 & n55353) | (n69566 & n55354) | (n55353 & n55354);
  assign n55356 = n29586 | n55273;
  assign n55357 = n29155 | n29586;
  assign n55358 = (n69566 & n55356) | (n69566 & n55357) | (n55356 & n55357);
  assign n29589 = ~n55355 & n55358;
  assign n29590 = x150 & x193;
  assign n29591 = n29589 & n29590;
  assign n29592 = n29589 | n29590;
  assign n29593 = ~n29591 & n29592;
  assign n55359 = n29162 & n29593;
  assign n69826 = (n29593 & n55166) | (n29593 & n55359) | (n55166 & n55359);
  assign n69827 = (n29593 & n55165) | (n29593 & n55359) | (n55165 & n55359);
  assign n69828 = (n69432 & n69826) | (n69432 & n69827) | (n69826 & n69827);
  assign n55361 = n29162 | n29593;
  assign n69829 = n55166 | n55361;
  assign n69830 = n55165 | n55361;
  assign n69831 = (n69432 & n69829) | (n69432 & n69830) | (n69829 & n69830);
  assign n29596 = ~n69828 & n69831;
  assign n29597 = x149 & x194;
  assign n29598 = n29596 & n29597;
  assign n29599 = n29596 | n29597;
  assign n29600 = ~n29598 & n29599;
  assign n29601 = n69717 & n29600;
  assign n29602 = n69717 | n29600;
  assign n29603 = ~n29601 & n29602;
  assign n29604 = x148 & x195;
  assign n29605 = n29603 & n29604;
  assign n29606 = n29603 | n29604;
  assign n29607 = ~n29605 & n29606;
  assign n55268 = n29176 | n29178;
  assign n55363 = n29607 & n55268;
  assign n55364 = n29176 & n29607;
  assign n55365 = (n69561 & n55363) | (n69561 & n55364) | (n55363 & n55364);
  assign n55366 = n29607 | n55268;
  assign n55367 = n29176 | n29607;
  assign n55368 = (n69561 & n55366) | (n69561 & n55367) | (n55366 & n55367);
  assign n29610 = ~n55365 & n55368;
  assign n29611 = x147 & x196;
  assign n29612 = n29610 & n29611;
  assign n29613 = n29610 | n29611;
  assign n29614 = ~n29612 & n29613;
  assign n55369 = n29183 & n29614;
  assign n69832 = (n29614 & n55176) | (n29614 & n55369) | (n55176 & n55369);
  assign n69833 = (n29614 & n55175) | (n29614 & n55369) | (n55175 & n55369);
  assign n69834 = (n69427 & n69832) | (n69427 & n69833) | (n69832 & n69833);
  assign n55371 = n29183 | n29614;
  assign n69835 = n55176 | n55371;
  assign n69836 = n55175 | n55371;
  assign n69837 = (n69427 & n69835) | (n69427 & n69836) | (n69835 & n69836);
  assign n29617 = ~n69834 & n69837;
  assign n29618 = x146 & x197;
  assign n29619 = n29617 & n29618;
  assign n29620 = n29617 | n29618;
  assign n29621 = ~n29619 & n29620;
  assign n29622 = n69712 & n29621;
  assign n29623 = n69712 | n29621;
  assign n29624 = ~n29622 & n29623;
  assign n29625 = x145 & x198;
  assign n29626 = n29624 & n29625;
  assign n29627 = n29624 | n29625;
  assign n29628 = ~n29626 & n29627;
  assign n55263 = n29197 | n29199;
  assign n55373 = n29628 & n55263;
  assign n55374 = n29197 & n29628;
  assign n55375 = (n55063 & n55373) | (n55063 & n55374) | (n55373 & n55374);
  assign n55376 = n29628 | n55263;
  assign n55377 = n29197 | n29628;
  assign n55378 = (n55063 & n55376) | (n55063 & n55377) | (n55376 & n55377);
  assign n29631 = ~n55375 & n55378;
  assign n29632 = x144 & x199;
  assign n29633 = n29631 & n29632;
  assign n29634 = n29631 | n29632;
  assign n29635 = ~n29633 & n29634;
  assign n55379 = n29204 & n29635;
  assign n55380 = (n29635 & n69688) | (n29635 & n55379) | (n69688 & n55379);
  assign n55381 = n29204 | n29635;
  assign n55382 = n69688 | n55381;
  assign n29638 = ~n55380 & n55382;
  assign n29639 = x143 & x200;
  assign n29640 = n29638 & n29639;
  assign n29641 = n29638 | n29639;
  assign n29642 = ~n29640 & n29641;
  assign n55383 = n29211 & n29642;
  assign n55384 = (n29642 & n55190) | (n29642 & n55383) | (n55190 & n55383);
  assign n55385 = n29211 | n29642;
  assign n55386 = n55190 | n55385;
  assign n29645 = ~n55384 & n55386;
  assign n29646 = x142 & x201;
  assign n29647 = n29645 & n29646;
  assign n29648 = n29645 | n29646;
  assign n29649 = ~n29647 & n29648;
  assign n55387 = n29218 & n29649;
  assign n55388 = (n29649 & n55194) | (n29649 & n55387) | (n55194 & n55387);
  assign n55389 = n29218 | n29649;
  assign n55390 = n55194 | n55389;
  assign n29652 = ~n55388 & n55390;
  assign n29653 = x141 & x202;
  assign n29654 = n29652 & n29653;
  assign n29655 = n29652 | n29653;
  assign n29656 = ~n29654 & n29655;
  assign n55391 = n29225 & n29656;
  assign n55392 = (n29656 & n55198) | (n29656 & n55391) | (n55198 & n55391);
  assign n55393 = n29225 | n29656;
  assign n55394 = n55198 | n55393;
  assign n29659 = ~n55392 & n55394;
  assign n29660 = x140 & x203;
  assign n29661 = n29659 & n29660;
  assign n29662 = n29659 | n29660;
  assign n29663 = ~n29661 & n29662;
  assign n55395 = n29232 & n29663;
  assign n55396 = (n29663 & n55202) | (n29663 & n55395) | (n55202 & n55395);
  assign n55397 = n29232 | n29663;
  assign n55398 = n55202 | n55397;
  assign n29666 = ~n55396 & n55398;
  assign n29667 = x139 & x204;
  assign n29668 = n29666 & n29667;
  assign n29669 = n29666 | n29667;
  assign n29670 = ~n29668 & n29669;
  assign n55399 = n29239 & n29670;
  assign n55400 = (n29670 & n55206) | (n29670 & n55399) | (n55206 & n55399);
  assign n55401 = n29239 | n29670;
  assign n55402 = n55206 | n55401;
  assign n29673 = ~n55400 & n55402;
  assign n29674 = x138 & x205;
  assign n29675 = n29673 & n29674;
  assign n29676 = n29673 | n29674;
  assign n29677 = ~n29675 & n29676;
  assign n55403 = n29246 & n29677;
  assign n55404 = (n29677 & n55210) | (n29677 & n55403) | (n55210 & n55403);
  assign n55405 = n29246 | n29677;
  assign n55406 = n55210 | n55405;
  assign n29680 = ~n55404 & n55406;
  assign n29681 = x137 & x206;
  assign n29682 = n29680 & n29681;
  assign n29683 = n29680 | n29681;
  assign n29684 = ~n29682 & n29683;
  assign n55407 = n29253 & n29684;
  assign n55408 = (n29684 & n55214) | (n29684 & n55407) | (n55214 & n55407);
  assign n55409 = n29253 | n29684;
  assign n55410 = n55214 | n55409;
  assign n29687 = ~n55408 & n55410;
  assign n29688 = x136 & x207;
  assign n29689 = n29687 & n29688;
  assign n29690 = n29687 | n29688;
  assign n29691 = ~n29689 & n29690;
  assign n55411 = n29260 & n29691;
  assign n55412 = (n29691 & n55218) | (n29691 & n55411) | (n55218 & n55411);
  assign n55413 = n29260 | n29691;
  assign n55414 = n55218 | n55413;
  assign n29694 = ~n55412 & n55414;
  assign n29695 = x135 & x208;
  assign n29696 = n29694 & n29695;
  assign n29697 = n29694 | n29695;
  assign n29698 = ~n29696 & n29697;
  assign n55415 = n29267 & n29698;
  assign n55416 = (n29698 & n55222) | (n29698 & n55415) | (n55222 & n55415);
  assign n55417 = n29267 | n29698;
  assign n55418 = n55222 | n55417;
  assign n29701 = ~n55416 & n55418;
  assign n29702 = x134 & x209;
  assign n29703 = n29701 & n29702;
  assign n29704 = n29701 | n29702;
  assign n29705 = ~n29703 & n29704;
  assign n55419 = n29274 & n29705;
  assign n55420 = (n29705 & n55226) | (n29705 & n55419) | (n55226 & n55419);
  assign n55421 = n29274 | n29705;
  assign n55422 = n55226 | n55421;
  assign n29708 = ~n55420 & n55422;
  assign n29709 = x133 & x210;
  assign n29710 = n29708 & n29709;
  assign n29711 = n29708 | n29709;
  assign n29712 = ~n29710 & n29711;
  assign n55423 = n29281 & n29712;
  assign n55424 = (n29712 & n55230) | (n29712 & n55423) | (n55230 & n55423);
  assign n55425 = n29281 | n29712;
  assign n55426 = n55230 | n55425;
  assign n29715 = ~n55424 & n55426;
  assign n29716 = x132 & x211;
  assign n29717 = n29715 & n29716;
  assign n29718 = n29715 | n29716;
  assign n29719 = ~n29717 & n29718;
  assign n55427 = n29288 & n29719;
  assign n55428 = (n29719 & n55234) | (n29719 & n55427) | (n55234 & n55427);
  assign n55429 = n29288 | n29719;
  assign n55430 = n55234 | n55429;
  assign n29722 = ~n55428 & n55430;
  assign n29723 = x131 & x212;
  assign n29724 = n29722 & n29723;
  assign n29725 = n29722 | n29723;
  assign n29726 = ~n29724 & n29725;
  assign n55431 = n29295 & n29726;
  assign n55432 = (n29726 & n55238) | (n29726 & n55431) | (n55238 & n55431);
  assign n55433 = n29295 | n29726;
  assign n55434 = n55238 | n55433;
  assign n29729 = ~n55432 & n55434;
  assign n29730 = x130 & x213;
  assign n29731 = n29729 & n29730;
  assign n29732 = n29729 | n29730;
  assign n29733 = ~n29731 & n29732;
  assign n55435 = n29302 & n29733;
  assign n55436 = (n29733 & n55243) | (n29733 & n55435) | (n55243 & n55435);
  assign n55437 = n29302 | n29733;
  assign n55438 = n55243 | n55437;
  assign n29736 = ~n55436 & n55438;
  assign n29737 = x129 & x214;
  assign n29738 = n29736 & n29737;
  assign n29739 = n29736 | n29737;
  assign n29740 = ~n29738 & n29739;
  assign n55261 = n29309 | n29311;
  assign n55439 = n29740 & n55261;
  assign n55440 = n29309 & n29740;
  assign n55441 = (n55058 & n55439) | (n55058 & n55440) | (n55439 & n55440);
  assign n55442 = n29740 | n55261;
  assign n55443 = n29309 | n29740;
  assign n55444 = (n55058 & n55442) | (n55058 & n55443) | (n55442 & n55443);
  assign n29743 = ~n55441 & n55444;
  assign n29744 = x128 & x215;
  assign n29745 = n29743 & n29744;
  assign n29746 = n29743 | n29744;
  assign n29747 = ~n29745 & n29746;
  assign n55259 = n29316 | n29318;
  assign n69838 = n29747 & n55259;
  assign n69839 = n29316 & n29747;
  assign n69840 = (n55056 & n69838) | (n55056 & n69839) | (n69838 & n69839);
  assign n69841 = n29747 | n55259;
  assign n69842 = n29316 | n29747;
  assign n69843 = (n55056 & n69841) | (n55056 & n69842) | (n69841 & n69842);
  assign n29750 = ~n69840 & n69843;
  assign n29751 = x127 & x216;
  assign n29752 = n29750 & n29751;
  assign n29753 = n29750 | n29751;
  assign n29754 = ~n29752 & n29753;
  assign n55257 = n29323 | n29325;
  assign n69844 = n29754 & n55257;
  assign n69845 = n29323 & n29754;
  assign n69846 = (n55054 & n69844) | (n55054 & n69845) | (n69844 & n69845);
  assign n69847 = n29754 | n55257;
  assign n69848 = n29323 | n29754;
  assign n69849 = (n55054 & n69847) | (n55054 & n69848) | (n69847 & n69848);
  assign n29757 = ~n69846 & n69849;
  assign n29758 = x126 & x217;
  assign n29759 = n29757 & n29758;
  assign n29760 = n29757 | n29758;
  assign n29761 = ~n29759 & n29760;
  assign n29762 = n55256 & n29761;
  assign n29763 = n55256 | n29761;
  assign n29764 = ~n29762 & n29763;
  assign n29765 = x125 & x218;
  assign n29766 = n29764 & n29765;
  assign n29767 = n29764 | n29765;
  assign n29768 = ~n29766 & n29767;
  assign n29769 = n55254 & n29768;
  assign n29770 = n55254 | n29768;
  assign n29771 = ~n29769 & n29770;
  assign n29772 = x124 & x219;
  assign n29773 = n29771 & n29772;
  assign n29774 = n29771 | n29772;
  assign n29775 = ~n29773 & n29774;
  assign n29776 = n55252 & n29775;
  assign n29777 = n55252 | n29775;
  assign n29778 = ~n29776 & n29777;
  assign n29779 = x123 & x220;
  assign n29780 = n29778 & n29779;
  assign n29781 = n29778 | n29779;
  assign n29782 = ~n29780 & n29781;
  assign n29783 = n29433 & n29782;
  assign n29784 = n29433 | n29782;
  assign n29785 = ~n29783 & n29784;
  assign n29786 = x122 & x221;
  assign n29787 = n29785 & n29786;
  assign n29788 = n29785 | n29786;
  assign n29789 = ~n29787 & n29788;
  assign n29790 = n29432 & n29789;
  assign n29791 = n29432 | n29789;
  assign n29792 = ~n29790 & n29791;
  assign n29793 = x121 & x222;
  assign n29794 = n29792 & n29793;
  assign n29795 = n29792 | n29793;
  assign n29796 = ~n29794 & n29795;
  assign n29797 = n29431 & n29796;
  assign n29798 = n29431 | n29796;
  assign n29799 = ~n29797 & n29798;
  assign n29800 = x120 & x223;
  assign n29801 = n29799 & n29800;
  assign n29802 = n29799 | n29800;
  assign n29803 = ~n29801 & n29802;
  assign n29804 = n29430 & n29803;
  assign n29805 = n29430 | n29803;
  assign n29806 = ~n29804 & n29805;
  assign n29807 = x119 & x224;
  assign n29808 = n29806 & n29807;
  assign n29809 = n29806 | n29807;
  assign n29810 = ~n29808 & n29809;
  assign n29811 = n29429 & n29810;
  assign n29812 = n29429 | n29810;
  assign n29813 = ~n29811 & n29812;
  assign n29814 = x118 & x225;
  assign n29815 = n29813 & n29814;
  assign n29816 = n29813 | n29814;
  assign n29817 = ~n29815 & n29816;
  assign n29818 = n29428 & n29817;
  assign n29819 = n29428 | n29817;
  assign n29820 = ~n29818 & n29819;
  assign n29821 = x117 & x226;
  assign n29822 = n29820 & n29821;
  assign n29823 = n29820 | n29821;
  assign n29824 = ~n29822 & n29823;
  assign n29825 = n29427 & n29824;
  assign n29826 = n29427 | n29824;
  assign n29827 = ~n29825 & n29826;
  assign n29828 = x116 & x227;
  assign n29829 = n29827 & n29828;
  assign n29830 = n29827 | n29828;
  assign n29831 = ~n29829 & n29830;
  assign n29832 = n69707 & n29831;
  assign n29833 = n69707 | n29831;
  assign n29834 = ~n29832 & n29833;
  assign n29835 = x115 & x228;
  assign n29836 = n29834 & n29835;
  assign n29837 = n29834 | n29835;
  assign n29838 = ~n29836 & n29837;
  assign n29839 = n55250 & n29838;
  assign n29840 = n55250 | n29838;
  assign n29841 = ~n29839 & n29840;
  assign n29842 = x114 & x229;
  assign n29843 = n29841 & n29842;
  assign n29844 = n29841 | n29842;
  assign n29845 = ~n29843 & n29844;
  assign n29846 = n55248 & n29845;
  assign n29847 = n55248 | n29845;
  assign n29848 = ~n29846 & n29847;
  assign n29849 = x113 & x230;
  assign n29850 = n29848 & n29849;
  assign n29851 = n29848 | n29849;
  assign n29852 = ~n29850 & n29851;
  assign n29853 = n29421 & n29852;
  assign n29854 = n29421 | n29852;
  assign n29855 = ~n29853 & n29854;
  assign n29856 = x112 & x231;
  assign n29857 = n29855 & n29856;
  assign n29858 = n29855 | n29856;
  assign n29859 = ~n29857 & n29858;
  assign n69850 = n29421 | n29849;
  assign n69851 = (n29421 & n29848) | (n29421 & n69850) | (n29848 & n69850);
  assign n55446 = (n29850 & n29852) | (n29850 & n69851) | (n29852 & n69851);
  assign n55447 = n29843 | n55248;
  assign n55448 = (n29843 & n29845) | (n29843 & n55447) | (n29845 & n55447);
  assign n55449 = n29836 | n55250;
  assign n55450 = (n29836 & n29838) | (n29836 & n55449) | (n29838 & n55449);
  assign n69852 = n29829 | n69707;
  assign n69853 = (n29829 & n29831) | (n29829 & n69852) | (n29831 & n69852);
  assign n29864 = n29822 | n29825;
  assign n29865 = n29815 | n29818;
  assign n29866 = n29808 | n29811;
  assign n29867 = n29801 | n29804;
  assign n29868 = n29794 | n29797;
  assign n29869 = n29787 | n29790;
  assign n55451 = n29780 | n29782;
  assign n55452 = (n29433 & n29780) | (n29433 & n55451) | (n29780 & n55451);
  assign n55453 = n29773 | n29775;
  assign n55454 = (n29773 & n55252) | (n29773 & n55453) | (n55252 & n55453);
  assign n55455 = n29766 | n29768;
  assign n55456 = (n29766 & n55254) | (n29766 & n55455) | (n55254 & n55455);
  assign n55258 = (n29323 & n55054) | (n29323 & n55257) | (n55054 & n55257);
  assign n55260 = (n29316 & n55056) | (n29316 & n55259) | (n55056 & n55259);
  assign n55469 = n29612 | n29614;
  assign n69856 = n29183 | n29612;
  assign n69857 = (n29612 & n29614) | (n29612 & n69856) | (n29614 & n69856);
  assign n69858 = (n55176 & n55469) | (n55176 & n69857) | (n55469 & n69857);
  assign n69859 = (n55175 & n55469) | (n55175 & n69857) | (n55469 & n69857);
  assign n69860 = (n69427 & n69858) | (n69427 & n69859) | (n69858 & n69859);
  assign n55474 = n29591 | n29593;
  assign n69861 = n29162 | n29591;
  assign n69862 = (n29591 & n29593) | (n29591 & n69861) | (n29593 & n69861);
  assign n69863 = (n55166 & n55474) | (n55166 & n69862) | (n55474 & n69862);
  assign n69864 = (n55165 & n55474) | (n55165 & n69862) | (n55474 & n69862);
  assign n69865 = (n69432 & n69863) | (n69432 & n69864) | (n69863 & n69864);
  assign n55277 = (n54961 & n69719) | (n54961 & n55276) | (n69719 & n55276);
  assign n55479 = n29570 | n29572;
  assign n69866 = n29141 | n29570;
  assign n69867 = (n29570 & n29572) | (n29570 & n69866) | (n29572 & n69866);
  assign n69868 = (n55156 & n55479) | (n55156 & n69867) | (n55479 & n69867);
  assign n69869 = (n55155 & n55479) | (n55155 & n69867) | (n55479 & n69867);
  assign n69870 = (n54873 & n69868) | (n54873 & n69869) | (n69868 & n69869);
  assign n55282 = (n54951 & n69721) | (n54951 & n55281) | (n69721 & n55281);
  assign n55484 = n29549 | n29551;
  assign n69871 = n29120 | n29549;
  assign n69872 = (n29549 & n29551) | (n29549 & n69871) | (n29551 & n69871);
  assign n69873 = (n55145 & n55484) | (n55145 & n69872) | (n55484 & n69872);
  assign n69874 = (n55146 & n55484) | (n55146 & n69872) | (n55484 & n69872);
  assign n69875 = (n54878 & n69873) | (n54878 & n69874) | (n69873 & n69874);
  assign n69878 = n29521 | n29523;
  assign n69879 = (n29521 & n55291) | (n29521 & n69878) | (n55291 & n69878);
  assign n69880 = n29092 | n29521;
  assign n69881 = (n29521 & n29523) | (n29521 & n69880) | (n29523 & n69880);
  assign n69882 = (n69580 & n69879) | (n69580 & n69881) | (n69879 & n69881);
  assign n69883 = (n69582 & n69879) | (n69582 & n69881) | (n69879 & n69881);
  assign n69884 = (n69331 & n69882) | (n69331 & n69883) | (n69882 & n69883);
  assign n55506 = n29486 | n69759;
  assign n55507 = n29486 | n69761;
  assign n69885 = (n55506 & n55507) | (n55506 & n69221) | (n55507 & n69221);
  assign n69886 = (n55506 & n55507) | (n55506 & n69220) | (n55507 & n69220);
  assign n69887 = (n68389 & n69885) | (n68389 & n69886) | (n69885 & n69886);
  assign n29914 = x168 & x176;
  assign n29915 = x167 & x177;
  assign n29916 = n29914 & n29915;
  assign n29917 = n29914 | n29915;
  assign n29918 = ~n29916 & n29917;
  assign n55509 = n29479 | n29481;
  assign n55511 = n29918 & n55509;
  assign n55512 = n29479 & n29918;
  assign n69888 = (n55511 & n55512) | (n55511 & n69747) | (n55512 & n69747);
  assign n69889 = (n55511 & n55512) | (n55511 & n69746) | (n55512 & n69746);
  assign n69890 = (n68195 & n69888) | (n68195 & n69889) | (n69888 & n69889);
  assign n55514 = n29918 | n55509;
  assign n55515 = n29479 | n29918;
  assign n69891 = (n55514 & n55515) | (n55514 & n69747) | (n55515 & n69747);
  assign n69892 = (n55514 & n55515) | (n55514 & n69746) | (n55515 & n69746);
  assign n69893 = (n68195 & n69891) | (n68195 & n69892) | (n69891 & n69892);
  assign n29921 = ~n69890 & n69893;
  assign n29922 = x166 & x178;
  assign n29923 = n29921 & n29922;
  assign n29924 = n29921 | n29922;
  assign n29925 = ~n29923 & n29924;
  assign n29926 = n69887 & n29925;
  assign n29927 = n69887 | n29925;
  assign n29928 = ~n29926 & n29927;
  assign n29929 = x165 & x179;
  assign n29930 = n29928 & n29929;
  assign n29931 = n29928 | n29929;
  assign n29932 = ~n29930 & n29931;
  assign n69894 = n29493 | n29495;
  assign n69895 = (n29493 & n55301) | (n29493 & n69894) | (n55301 & n69894);
  assign n55517 = n29932 & n69895;
  assign n69896 = n29064 | n29493;
  assign n69897 = (n29493 & n29495) | (n29493 & n69896) | (n29495 & n69896);
  assign n55518 = n29932 & n69897;
  assign n69898 = (n55517 & n55518) | (n55517 & n69590) | (n55518 & n69590);
  assign n69899 = (n55517 & n55518) | (n55517 & n69589) | (n55518 & n69589);
  assign n69900 = (n68776 & n69898) | (n68776 & n69899) | (n69898 & n69899);
  assign n55520 = n29932 | n69895;
  assign n55521 = n29932 | n69897;
  assign n69901 = (n55520 & n55521) | (n55520 & n69590) | (n55521 & n69590);
  assign n69902 = (n55520 & n55521) | (n55520 & n69589) | (n55521 & n69589);
  assign n69903 = (n68776 & n69901) | (n68776 & n69902) | (n69901 & n69902);
  assign n29935 = ~n69900 & n69903;
  assign n29936 = x164 & x180;
  assign n29937 = n29935 & n29936;
  assign n29938 = n29935 | n29936;
  assign n29939 = ~n29937 & n29938;
  assign n55501 = n29500 | n29502;
  assign n55523 = n29939 & n55501;
  assign n55524 = n29500 & n29939;
  assign n69904 = (n55523 & n55524) | (n55523 & n69741) | (n55524 & n69741);
  assign n69905 = (n55523 & n55524) | (n55523 & n69740) | (n55524 & n69740);
  assign n69906 = (n68982 & n69904) | (n68982 & n69905) | (n69904 & n69905);
  assign n55526 = n29939 | n55501;
  assign n55527 = n29500 | n29939;
  assign n69907 = (n55526 & n55527) | (n55526 & n69741) | (n55527 & n69741);
  assign n69908 = (n55526 & n55527) | (n55526 & n69740) | (n55527 & n69740);
  assign n69909 = (n68982 & n69907) | (n68982 & n69908) | (n69907 & n69908);
  assign n29942 = ~n69906 & n69909;
  assign n29943 = x163 & x181;
  assign n29944 = n29942 & n29943;
  assign n29945 = n29942 | n29943;
  assign n29946 = ~n29944 & n29945;
  assign n55499 = n29507 | n29509;
  assign n55529 = n29946 & n55499;
  assign n55530 = n29507 & n29946;
  assign n55531 = (n69736 & n55529) | (n69736 & n55530) | (n55529 & n55530);
  assign n55532 = n29946 | n55499;
  assign n55533 = n29507 | n29946;
  assign n55534 = (n69736 & n55532) | (n69736 & n55533) | (n55532 & n55533);
  assign n29949 = ~n55531 & n55534;
  assign n29950 = x162 & x182;
  assign n29951 = n29949 & n29950;
  assign n29952 = n29949 | n29950;
  assign n29953 = ~n29951 & n29952;
  assign n69912 = n29085 | n29514;
  assign n69913 = (n29514 & n29516) | (n29514 & n69912) | (n29516 & n69912);
  assign n55536 = n29953 & n69913;
  assign n69910 = n29514 & n29953;
  assign n69911 = (n29953 & n55321) | (n29953 & n69910) | (n55321 & n69910);
  assign n69914 = (n55536 & n69585) | (n55536 & n69911) | (n69585 & n69911);
  assign n69915 = (n55536 & n69584) | (n55536 & n69911) | (n69584 & n69911);
  assign n69916 = (n69244 & n69914) | (n69244 & n69915) | (n69914 & n69915);
  assign n55539 = n29953 | n69913;
  assign n69917 = n29514 | n29953;
  assign n69918 = n55321 | n69917;
  assign n69919 = (n55539 & n69585) | (n55539 & n69918) | (n69585 & n69918);
  assign n69920 = (n55539 & n69584) | (n55539 & n69918) | (n69584 & n69918);
  assign n69921 = (n69244 & n69919) | (n69244 & n69920) | (n69919 & n69920);
  assign n29956 = ~n69916 & n69921;
  assign n29957 = x161 & x183;
  assign n29958 = n29956 & n29957;
  assign n29959 = n29956 | n29957;
  assign n29960 = ~n29958 & n29959;
  assign n29961 = n69884 & n29960;
  assign n29962 = n69884 | n29960;
  assign n29963 = ~n29961 & n29962;
  assign n29964 = x160 & x184;
  assign n29965 = n29963 & n29964;
  assign n29966 = n29963 | n29964;
  assign n29967 = ~n29965 & n29966;
  assign n55491 = n29528 | n29530;
  assign n55541 = n29967 & n55491;
  assign n55542 = n29528 & n29967;
  assign n55543 = (n69730 & n55541) | (n69730 & n55542) | (n55541 & n55542);
  assign n55544 = n29967 | n55491;
  assign n55545 = n29528 | n29967;
  assign n55546 = (n69730 & n55544) | (n69730 & n55545) | (n55544 & n55545);
  assign n29970 = ~n55543 & n55546;
  assign n29971 = x159 & x185;
  assign n29972 = n29970 & n29971;
  assign n29973 = n29970 | n29971;
  assign n29974 = ~n29972 & n29973;
  assign n55489 = n29535 | n55333;
  assign n69922 = n29974 & n55489;
  assign n69876 = n29106 | n29535;
  assign n69877 = (n29535 & n29537) | (n29535 & n69876) | (n29537 & n69876);
  assign n69923 = n29974 & n69877;
  assign n69924 = (n69578 & n69922) | (n69578 & n69923) | (n69922 & n69923);
  assign n69925 = n29974 | n55489;
  assign n69926 = n29974 | n69877;
  assign n69927 = (n69578 & n69925) | (n69578 & n69926) | (n69925 & n69926);
  assign n29977 = ~n69924 & n69927;
  assign n29978 = x158 & x186;
  assign n29979 = n29977 & n29978;
  assign n29980 = n29977 | n29978;
  assign n29981 = ~n29979 & n29980;
  assign n55486 = n29542 | n29544;
  assign n55547 = n29981 & n55486;
  assign n55548 = n29542 & n29981;
  assign n69928 = (n55284 & n55547) | (n55284 & n55548) | (n55547 & n55548);
  assign n69929 = (n55547 & n55548) | (n55547 & n69723) | (n55548 & n69723);
  assign n69930 = (n54881 & n69928) | (n54881 & n69929) | (n69928 & n69929);
  assign n55550 = n29981 | n55486;
  assign n55551 = n29542 | n29981;
  assign n69931 = (n55284 & n55550) | (n55284 & n55551) | (n55550 & n55551);
  assign n69932 = (n55550 & n55551) | (n55550 & n69723) | (n55551 & n69723);
  assign n69933 = (n54881 & n69931) | (n54881 & n69932) | (n69931 & n69932);
  assign n29984 = ~n69930 & n69933;
  assign n29985 = x157 & x187;
  assign n29986 = n29984 & n29985;
  assign n29987 = n29984 | n29985;
  assign n29988 = ~n29986 & n29987;
  assign n29989 = n69875 & n29988;
  assign n29990 = n69875 | n29988;
  assign n29991 = ~n29989 & n29990;
  assign n29992 = x156 & x188;
  assign n29993 = n29991 & n29992;
  assign n29994 = n29991 | n29992;
  assign n29995 = ~n29993 & n29994;
  assign n55481 = n29556 | n29558;
  assign n55553 = n29995 & n55481;
  assign n55554 = n29556 & n29995;
  assign n55555 = (n55282 & n55553) | (n55282 & n55554) | (n55553 & n55554);
  assign n55556 = n29995 | n55481;
  assign n55557 = n29556 | n29995;
  assign n55558 = (n55282 & n55556) | (n55282 & n55557) | (n55556 & n55557);
  assign n29998 = ~n55555 & n55558;
  assign n29999 = x155 & x189;
  assign n30000 = n29998 & n29999;
  assign n30001 = n29998 | n29999;
  assign n30002 = ~n30000 & n30001;
  assign n55559 = n29563 & n30002;
  assign n55560 = (n30002 & n55345) | (n30002 & n55559) | (n55345 & n55559);
  assign n55561 = n29563 | n30002;
  assign n55562 = n55345 | n55561;
  assign n30005 = ~n55560 & n55562;
  assign n30006 = x154 & x190;
  assign n30007 = n30005 & n30006;
  assign n30008 = n30005 | n30006;
  assign n30009 = ~n30007 & n30008;
  assign n30010 = n69870 & n30009;
  assign n30011 = n69870 | n30009;
  assign n30012 = ~n30010 & n30011;
  assign n30013 = x153 & x191;
  assign n30014 = n30012 & n30013;
  assign n30015 = n30012 | n30013;
  assign n30016 = ~n30014 & n30015;
  assign n55476 = n29577 | n29579;
  assign n55563 = n30016 & n55476;
  assign n55564 = n29577 & n30016;
  assign n55565 = (n55277 & n55563) | (n55277 & n55564) | (n55563 & n55564);
  assign n55566 = n30016 | n55476;
  assign n55567 = n29577 | n30016;
  assign n55568 = (n55277 & n55566) | (n55277 & n55567) | (n55566 & n55567);
  assign n30019 = ~n55565 & n55568;
  assign n30020 = x152 & x192;
  assign n30021 = n30019 & n30020;
  assign n30022 = n30019 | n30020;
  assign n30023 = ~n30021 & n30022;
  assign n55569 = n29584 & n30023;
  assign n55570 = (n30023 & n55355) | (n30023 & n55569) | (n55355 & n55569);
  assign n55571 = n29584 | n30023;
  assign n55572 = n55355 | n55571;
  assign n30026 = ~n55570 & n55572;
  assign n30027 = x151 & x193;
  assign n30028 = n30026 & n30027;
  assign n30029 = n30026 | n30027;
  assign n30030 = ~n30028 & n30029;
  assign n30031 = n69865 & n30030;
  assign n30032 = n69865 | n30030;
  assign n30033 = ~n30031 & n30032;
  assign n30034 = x150 & x194;
  assign n30035 = n30033 & n30034;
  assign n30036 = n30033 | n30034;
  assign n30037 = ~n30035 & n30036;
  assign n55471 = n29598 | n29600;
  assign n55573 = n30037 & n55471;
  assign n55574 = n29598 & n30037;
  assign n55575 = (n69717 & n55573) | (n69717 & n55574) | (n55573 & n55574);
  assign n55576 = n30037 | n55471;
  assign n55577 = n29598 | n30037;
  assign n55578 = (n69717 & n55576) | (n69717 & n55577) | (n55576 & n55577);
  assign n30040 = ~n55575 & n55578;
  assign n30041 = x149 & x195;
  assign n30042 = n30040 & n30041;
  assign n30043 = n30040 | n30041;
  assign n30044 = ~n30042 & n30043;
  assign n55579 = n29605 & n30044;
  assign n69934 = (n30044 & n55364) | (n30044 & n55579) | (n55364 & n55579);
  assign n69935 = (n30044 & n55363) | (n30044 & n55579) | (n55363 & n55579);
  assign n69936 = (n69561 & n69934) | (n69561 & n69935) | (n69934 & n69935);
  assign n55581 = n29605 | n30044;
  assign n69937 = n55364 | n55581;
  assign n69938 = n55363 | n55581;
  assign n69939 = (n69561 & n69937) | (n69561 & n69938) | (n69937 & n69938);
  assign n30047 = ~n69936 & n69939;
  assign n30048 = x148 & x196;
  assign n30049 = n30047 & n30048;
  assign n30050 = n30047 | n30048;
  assign n30051 = ~n30049 & n30050;
  assign n30052 = n69860 & n30051;
  assign n30053 = n69860 | n30051;
  assign n30054 = ~n30052 & n30053;
  assign n30055 = x147 & x197;
  assign n30056 = n30054 & n30055;
  assign n30057 = n30054 | n30055;
  assign n30058 = ~n30056 & n30057;
  assign n55466 = n29619 | n29621;
  assign n55583 = n30058 & n55466;
  assign n55584 = n29619 & n30058;
  assign n55585 = (n69712 & n55583) | (n69712 & n55584) | (n55583 & n55584);
  assign n55586 = n30058 | n55466;
  assign n55587 = n29619 | n30058;
  assign n55588 = (n69712 & n55586) | (n69712 & n55587) | (n55586 & n55587);
  assign n30061 = ~n55585 & n55588;
  assign n30062 = x146 & x198;
  assign n30063 = n30061 & n30062;
  assign n30064 = n30061 | n30062;
  assign n30065 = ~n30063 & n30064;
  assign n55589 = n29626 & n30065;
  assign n69940 = (n30065 & n55374) | (n30065 & n55589) | (n55374 & n55589);
  assign n69941 = (n30065 & n55373) | (n30065 & n55589) | (n55373 & n55589);
  assign n69942 = (n55063 & n69940) | (n55063 & n69941) | (n69940 & n69941);
  assign n55591 = n29626 | n30065;
  assign n69943 = n55374 | n55591;
  assign n69944 = n55373 | n55591;
  assign n69945 = (n55063 & n69943) | (n55063 & n69944) | (n69943 & n69944);
  assign n30068 = ~n69942 & n69945;
  assign n30069 = x145 & x199;
  assign n30070 = n30068 & n30069;
  assign n30071 = n30068 | n30069;
  assign n30072 = ~n30070 & n30071;
  assign n55464 = n29633 | n29635;
  assign n69946 = n30072 & n55464;
  assign n69854 = n29204 | n29633;
  assign n69855 = (n29633 & n29635) | (n29633 & n69854) | (n29635 & n69854);
  assign n69947 = n30072 & n69855;
  assign n69948 = (n69688 & n69946) | (n69688 & n69947) | (n69946 & n69947);
  assign n69949 = n30072 | n55464;
  assign n69950 = n30072 | n69855;
  assign n69951 = (n69688 & n69949) | (n69688 & n69950) | (n69949 & n69950);
  assign n30075 = ~n69948 & n69951;
  assign n30076 = x144 & x200;
  assign n30077 = n30075 & n30076;
  assign n30078 = n30075 | n30076;
  assign n30079 = ~n30077 & n30078;
  assign n55593 = n29640 & n30079;
  assign n69952 = (n30079 & n55383) | (n30079 & n55593) | (n55383 & n55593);
  assign n69953 = (n29642 & n30079) | (n29642 & n55593) | (n30079 & n55593);
  assign n69954 = (n55190 & n69952) | (n55190 & n69953) | (n69952 & n69953);
  assign n55595 = n29640 | n30079;
  assign n69955 = n55383 | n55595;
  assign n69956 = n29642 | n55595;
  assign n69957 = (n55190 & n69955) | (n55190 & n69956) | (n69955 & n69956);
  assign n30082 = ~n69954 & n69957;
  assign n30083 = x143 & x201;
  assign n30084 = n30082 & n30083;
  assign n30085 = n30082 | n30083;
  assign n30086 = ~n30084 & n30085;
  assign n55597 = n29647 & n30086;
  assign n55598 = (n30086 & n55388) | (n30086 & n55597) | (n55388 & n55597);
  assign n55599 = n29647 | n30086;
  assign n55600 = n55388 | n55599;
  assign n30089 = ~n55598 & n55600;
  assign n30090 = x142 & x202;
  assign n30091 = n30089 & n30090;
  assign n30092 = n30089 | n30090;
  assign n30093 = ~n30091 & n30092;
  assign n55601 = n29654 & n30093;
  assign n55602 = (n30093 & n55392) | (n30093 & n55601) | (n55392 & n55601);
  assign n55603 = n29654 | n30093;
  assign n55604 = n55392 | n55603;
  assign n30096 = ~n55602 & n55604;
  assign n30097 = x141 & x203;
  assign n30098 = n30096 & n30097;
  assign n30099 = n30096 | n30097;
  assign n30100 = ~n30098 & n30099;
  assign n55605 = n29661 & n30100;
  assign n55606 = (n30100 & n55396) | (n30100 & n55605) | (n55396 & n55605);
  assign n55607 = n29661 | n30100;
  assign n55608 = n55396 | n55607;
  assign n30103 = ~n55606 & n55608;
  assign n30104 = x140 & x204;
  assign n30105 = n30103 & n30104;
  assign n30106 = n30103 | n30104;
  assign n30107 = ~n30105 & n30106;
  assign n55609 = n29668 & n30107;
  assign n55610 = (n30107 & n55400) | (n30107 & n55609) | (n55400 & n55609);
  assign n55611 = n29668 | n30107;
  assign n55612 = n55400 | n55611;
  assign n30110 = ~n55610 & n55612;
  assign n30111 = x139 & x205;
  assign n30112 = n30110 & n30111;
  assign n30113 = n30110 | n30111;
  assign n30114 = ~n30112 & n30113;
  assign n55613 = n29675 & n30114;
  assign n55614 = (n30114 & n55404) | (n30114 & n55613) | (n55404 & n55613);
  assign n55615 = n29675 | n30114;
  assign n55616 = n55404 | n55615;
  assign n30117 = ~n55614 & n55616;
  assign n30118 = x138 & x206;
  assign n30119 = n30117 & n30118;
  assign n30120 = n30117 | n30118;
  assign n30121 = ~n30119 & n30120;
  assign n55617 = n29682 & n30121;
  assign n55618 = (n30121 & n55408) | (n30121 & n55617) | (n55408 & n55617);
  assign n55619 = n29682 | n30121;
  assign n55620 = n55408 | n55619;
  assign n30124 = ~n55618 & n55620;
  assign n30125 = x137 & x207;
  assign n30126 = n30124 & n30125;
  assign n30127 = n30124 | n30125;
  assign n30128 = ~n30126 & n30127;
  assign n55621 = n29689 & n30128;
  assign n55622 = (n30128 & n55412) | (n30128 & n55621) | (n55412 & n55621);
  assign n55623 = n29689 | n30128;
  assign n55624 = n55412 | n55623;
  assign n30131 = ~n55622 & n55624;
  assign n30132 = x136 & x208;
  assign n30133 = n30131 & n30132;
  assign n30134 = n30131 | n30132;
  assign n30135 = ~n30133 & n30134;
  assign n55625 = n29696 & n30135;
  assign n55626 = (n30135 & n55416) | (n30135 & n55625) | (n55416 & n55625);
  assign n55627 = n29696 | n30135;
  assign n55628 = n55416 | n55627;
  assign n30138 = ~n55626 & n55628;
  assign n30139 = x135 & x209;
  assign n30140 = n30138 & n30139;
  assign n30141 = n30138 | n30139;
  assign n30142 = ~n30140 & n30141;
  assign n55629 = n29703 & n30142;
  assign n55630 = (n30142 & n55420) | (n30142 & n55629) | (n55420 & n55629);
  assign n55631 = n29703 | n30142;
  assign n55632 = n55420 | n55631;
  assign n30145 = ~n55630 & n55632;
  assign n30146 = x134 & x210;
  assign n30147 = n30145 & n30146;
  assign n30148 = n30145 | n30146;
  assign n30149 = ~n30147 & n30148;
  assign n55633 = n29710 & n30149;
  assign n55634 = (n30149 & n55424) | (n30149 & n55633) | (n55424 & n55633);
  assign n55635 = n29710 | n30149;
  assign n55636 = n55424 | n55635;
  assign n30152 = ~n55634 & n55636;
  assign n30153 = x133 & x211;
  assign n30154 = n30152 & n30153;
  assign n30155 = n30152 | n30153;
  assign n30156 = ~n30154 & n30155;
  assign n55637 = n29717 & n30156;
  assign n55638 = (n30156 & n55428) | (n30156 & n55637) | (n55428 & n55637);
  assign n55639 = n29717 | n30156;
  assign n55640 = n55428 | n55639;
  assign n30159 = ~n55638 & n55640;
  assign n30160 = x132 & x212;
  assign n30161 = n30159 & n30160;
  assign n30162 = n30159 | n30160;
  assign n30163 = ~n30161 & n30162;
  assign n55641 = n29724 & n30163;
  assign n55642 = (n30163 & n55432) | (n30163 & n55641) | (n55432 & n55641);
  assign n55643 = n29724 | n30163;
  assign n55644 = n55432 | n55643;
  assign n30166 = ~n55642 & n55644;
  assign n30167 = x131 & x213;
  assign n30168 = n30166 & n30167;
  assign n30169 = n30166 | n30167;
  assign n30170 = ~n30168 & n30169;
  assign n55645 = n29731 & n30170;
  assign n55646 = (n30170 & n55436) | (n30170 & n55645) | (n55436 & n55645);
  assign n55647 = n29731 | n30170;
  assign n55648 = n55436 | n55647;
  assign n30173 = ~n55646 & n55648;
  assign n30174 = x130 & x214;
  assign n30175 = n30173 & n30174;
  assign n30176 = n30173 | n30174;
  assign n30177 = ~n30175 & n30176;
  assign n55649 = n29738 & n30177;
  assign n55650 = (n30177 & n55441) | (n30177 & n55649) | (n55441 & n55649);
  assign n55651 = n29738 | n30177;
  assign n55652 = n55441 | n55651;
  assign n30180 = ~n55650 & n55652;
  assign n30181 = x129 & x215;
  assign n30182 = n30180 & n30181;
  assign n30183 = n30180 | n30181;
  assign n30184 = ~n30182 & n30183;
  assign n55461 = n29745 | n29747;
  assign n55653 = n30184 & n55461;
  assign n55654 = n29745 & n30184;
  assign n55655 = (n55260 & n55653) | (n55260 & n55654) | (n55653 & n55654);
  assign n55656 = n30184 | n55461;
  assign n55657 = n29745 | n30184;
  assign n55658 = (n55260 & n55656) | (n55260 & n55657) | (n55656 & n55657);
  assign n30187 = ~n55655 & n55658;
  assign n30188 = x128 & x216;
  assign n30189 = n30187 & n30188;
  assign n30190 = n30187 | n30188;
  assign n30191 = ~n30189 & n30190;
  assign n55459 = n29752 | n29754;
  assign n69958 = n30191 & n55459;
  assign n69959 = n29752 & n30191;
  assign n69960 = (n55258 & n69958) | (n55258 & n69959) | (n69958 & n69959);
  assign n69961 = n30191 | n55459;
  assign n69962 = n29752 | n30191;
  assign n69963 = (n55258 & n69961) | (n55258 & n69962) | (n69961 & n69962);
  assign n30194 = ~n69960 & n69963;
  assign n30195 = x127 & x217;
  assign n30196 = n30194 & n30195;
  assign n30197 = n30194 | n30195;
  assign n30198 = ~n30196 & n30197;
  assign n55457 = n29759 | n29761;
  assign n69964 = n30198 & n55457;
  assign n69965 = n29759 & n30198;
  assign n69966 = (n55256 & n69964) | (n55256 & n69965) | (n69964 & n69965);
  assign n69967 = n30198 | n55457;
  assign n69968 = n29759 | n30198;
  assign n69969 = (n55256 & n69967) | (n55256 & n69968) | (n69967 & n69968);
  assign n30201 = ~n69966 & n69969;
  assign n30202 = x126 & x218;
  assign n30203 = n30201 & n30202;
  assign n30204 = n30201 | n30202;
  assign n30205 = ~n30203 & n30204;
  assign n30206 = n55456 & n30205;
  assign n30207 = n55456 | n30205;
  assign n30208 = ~n30206 & n30207;
  assign n30209 = x125 & x219;
  assign n30210 = n30208 & n30209;
  assign n30211 = n30208 | n30209;
  assign n30212 = ~n30210 & n30211;
  assign n30213 = n55454 & n30212;
  assign n30214 = n55454 | n30212;
  assign n30215 = ~n30213 & n30214;
  assign n30216 = x124 & x220;
  assign n30217 = n30215 & n30216;
  assign n30218 = n30215 | n30216;
  assign n30219 = ~n30217 & n30218;
  assign n30220 = n55452 & n30219;
  assign n30221 = n55452 | n30219;
  assign n30222 = ~n30220 & n30221;
  assign n30223 = x123 & x221;
  assign n30224 = n30222 & n30223;
  assign n30225 = n30222 | n30223;
  assign n30226 = ~n30224 & n30225;
  assign n30227 = n29869 & n30226;
  assign n30228 = n29869 | n30226;
  assign n30229 = ~n30227 & n30228;
  assign n30230 = x122 & x222;
  assign n30231 = n30229 & n30230;
  assign n30232 = n30229 | n30230;
  assign n30233 = ~n30231 & n30232;
  assign n30234 = n29868 & n30233;
  assign n30235 = n29868 | n30233;
  assign n30236 = ~n30234 & n30235;
  assign n30237 = x121 & x223;
  assign n30238 = n30236 & n30237;
  assign n30239 = n30236 | n30237;
  assign n30240 = ~n30238 & n30239;
  assign n30241 = n29867 & n30240;
  assign n30242 = n29867 | n30240;
  assign n30243 = ~n30241 & n30242;
  assign n30244 = x120 & x224;
  assign n30245 = n30243 & n30244;
  assign n30246 = n30243 | n30244;
  assign n30247 = ~n30245 & n30246;
  assign n30248 = n29866 & n30247;
  assign n30249 = n29866 | n30247;
  assign n30250 = ~n30248 & n30249;
  assign n30251 = x119 & x225;
  assign n30252 = n30250 & n30251;
  assign n30253 = n30250 | n30251;
  assign n30254 = ~n30252 & n30253;
  assign n30255 = n29865 & n30254;
  assign n30256 = n29865 | n30254;
  assign n30257 = ~n30255 & n30256;
  assign n30258 = x118 & x226;
  assign n30259 = n30257 & n30258;
  assign n30260 = n30257 | n30258;
  assign n30261 = ~n30259 & n30260;
  assign n30262 = n29864 & n30261;
  assign n30263 = n29864 | n30261;
  assign n30264 = ~n30262 & n30263;
  assign n30265 = x117 & x227;
  assign n30266 = n30264 & n30265;
  assign n30267 = n30264 | n30265;
  assign n30268 = ~n30266 & n30267;
  assign n30269 = n69853 & n30268;
  assign n30270 = n69853 | n30268;
  assign n30271 = ~n30269 & n30270;
  assign n30272 = x116 & x228;
  assign n30273 = n30271 & n30272;
  assign n30274 = n30271 | n30272;
  assign n30275 = ~n30273 & n30274;
  assign n30276 = n55450 & n30275;
  assign n30277 = n55450 | n30275;
  assign n30278 = ~n30276 & n30277;
  assign n30279 = x115 & x229;
  assign n30280 = n30278 & n30279;
  assign n30281 = n30278 | n30279;
  assign n30282 = ~n30280 & n30281;
  assign n30283 = n55448 & n30282;
  assign n30284 = n55448 | n30282;
  assign n30285 = ~n30283 & n30284;
  assign n30286 = x114 & x230;
  assign n30287 = n30285 & n30286;
  assign n30288 = n30285 | n30286;
  assign n30289 = ~n30287 & n30288;
  assign n30290 = n55446 & n30289;
  assign n30291 = n55446 | n30289;
  assign n30292 = ~n30290 & n30291;
  assign n30293 = x113 & x231;
  assign n30294 = n30292 & n30293;
  assign n30295 = n30292 | n30293;
  assign n30296 = ~n30294 & n30295;
  assign n30297 = n29857 & n30296;
  assign n30298 = n29857 | n30296;
  assign n30299 = ~n30297 & n30298;
  assign n30300 = x112 & x232;
  assign n30301 = n30299 & n30300;
  assign n30302 = n30299 | n30300;
  assign n30303 = ~n30301 & n30302;
  assign n69970 = n29857 | n30293;
  assign n69971 = (n29857 & n30292) | (n29857 & n69970) | (n30292 & n69970);
  assign n55660 = (n30294 & n30296) | (n30294 & n69971) | (n30296 & n69971);
  assign n55661 = n30287 | n55446;
  assign n55662 = (n30287 & n30289) | (n30287 & n55661) | (n30289 & n55661);
  assign n55663 = n30280 | n55448;
  assign n55664 = (n30280 & n30282) | (n30280 & n55663) | (n30282 & n55663);
  assign n55665 = n30273 | n55450;
  assign n55666 = (n30273 & n30275) | (n30273 & n55665) | (n30275 & n55665);
  assign n69972 = n30266 | n69853;
  assign n69973 = (n30266 & n30268) | (n30266 & n69972) | (n30268 & n69972);
  assign n30309 = n30259 | n30262;
  assign n30310 = n30252 | n30255;
  assign n30311 = n30245 | n30248;
  assign n30312 = n30238 | n30241;
  assign n30313 = n30231 | n30234;
  assign n55667 = n30224 | n30226;
  assign n55668 = (n29869 & n30224) | (n29869 & n55667) | (n30224 & n55667);
  assign n55669 = n30217 | n30219;
  assign n55670 = (n30217 & n55452) | (n30217 & n55669) | (n55452 & n55669);
  assign n55671 = n30210 | n30212;
  assign n55672 = (n30210 & n55454) | (n30210 & n55671) | (n55454 & n55671);
  assign n55458 = (n29759 & n55256) | (n29759 & n55457) | (n55256 & n55457);
  assign n55460 = (n29752 & n55258) | (n29752 & n55459) | (n55258 & n55459);
  assign n55465 = (n69688 & n69855) | (n69688 & n55464) | (n69855 & n55464);
  assign n55682 = n30063 | n30065;
  assign n69974 = n29626 | n30063;
  assign n69975 = (n30063 & n30065) | (n30063 & n69974) | (n30065 & n69974);
  assign n69976 = (n55374 & n55682) | (n55374 & n69975) | (n55682 & n69975);
  assign n69977 = (n55373 & n55682) | (n55373 & n69975) | (n55682 & n69975);
  assign n69978 = (n55063 & n69976) | (n55063 & n69977) | (n69976 & n69977);
  assign n55687 = n30042 | n30044;
  assign n69979 = n29605 | n30042;
  assign n69980 = (n30042 & n30044) | (n30042 & n69979) | (n30044 & n69979);
  assign n69981 = (n55364 & n55687) | (n55364 & n69980) | (n55687 & n69980);
  assign n69982 = (n55363 & n55687) | (n55363 & n69980) | (n55687 & n69980);
  assign n69983 = (n69561 & n69981) | (n69561 & n69982) | (n69981 & n69982);
  assign n69988 = n29542 | n29979;
  assign n69989 = (n29979 & n29981) | (n29979 & n69988) | (n29981 & n69988);
  assign n69990 = n29979 | n29981;
  assign n69991 = (n29979 & n55486) | (n29979 & n69990) | (n55486 & n69990);
  assign n69992 = (n55284 & n69989) | (n55284 & n69991) | (n69989 & n69991);
  assign n69993 = (n69723 & n69989) | (n69723 & n69991) | (n69989 & n69991);
  assign n69994 = (n54881 & n69992) | (n54881 & n69993) | (n69992 & n69993);
  assign n30359 = x169 & x176;
  assign n30360 = x168 & x177;
  assign n30361 = n30359 & n30360;
  assign n30362 = n30359 | n30360;
  assign n30363 = ~n30361 & n30362;
  assign n69997 = n29916 | n29918;
  assign n69998 = (n29916 & n55509) | (n29916 & n69997) | (n55509 & n69997);
  assign n55725 = n30363 & n69998;
  assign n69999 = n29479 | n29916;
  assign n70000 = (n29916 & n29918) | (n29916 & n69999) | (n29918 & n69999);
  assign n55726 = n30363 & n70000;
  assign n70001 = (n55725 & n55726) | (n55725 & n69747) | (n55726 & n69747);
  assign n70002 = (n55725 & n55726) | (n55725 & n69746) | (n55726 & n69746);
  assign n70003 = (n68195 & n70001) | (n68195 & n70002) | (n70001 & n70002);
  assign n55728 = n30363 | n69998;
  assign n55729 = n30363 | n70000;
  assign n70004 = (n55728 & n55729) | (n55728 & n69747) | (n55729 & n69747);
  assign n70005 = (n55728 & n55729) | (n55728 & n69746) | (n55729 & n69746);
  assign n70006 = (n68195 & n70004) | (n68195 & n70005) | (n70004 & n70005);
  assign n30366 = ~n70003 & n70006;
  assign n30367 = x167 & x178;
  assign n30368 = n30366 & n30367;
  assign n30369 = n30366 | n30367;
  assign n30370 = ~n30368 & n30369;
  assign n55720 = n29923 | n29925;
  assign n55731 = n30370 & n55720;
  assign n55732 = n29923 & n30370;
  assign n55733 = (n69887 & n55731) | (n69887 & n55732) | (n55731 & n55732);
  assign n55734 = n30370 | n55720;
  assign n55735 = n29923 | n30370;
  assign n55736 = (n69887 & n55734) | (n69887 & n55735) | (n55734 & n55735);
  assign n30373 = ~n55733 & n55736;
  assign n30374 = x166 & x179;
  assign n30375 = n30373 & n30374;
  assign n30376 = n30373 | n30374;
  assign n30377 = ~n30375 & n30376;
  assign n70007 = n29930 | n29932;
  assign n70008 = (n29930 & n69895) | (n29930 & n70007) | (n69895 & n70007);
  assign n55737 = n30377 & n70008;
  assign n70009 = n29930 & n30377;
  assign n70010 = (n30377 & n55518) | (n30377 & n70009) | (n55518 & n70009);
  assign n70011 = (n55737 & n69590) | (n55737 & n70010) | (n69590 & n70010);
  assign n70012 = (n55737 & n69589) | (n55737 & n70010) | (n69589 & n70010);
  assign n70013 = (n68776 & n70011) | (n68776 & n70012) | (n70011 & n70012);
  assign n55740 = n30377 | n70008;
  assign n70014 = n29930 | n30377;
  assign n70015 = n55518 | n70014;
  assign n70016 = (n55740 & n69590) | (n55740 & n70015) | (n69590 & n70015);
  assign n70017 = (n55740 & n69589) | (n55740 & n70015) | (n69589 & n70015);
  assign n70018 = (n68776 & n70016) | (n68776 & n70017) | (n70016 & n70017);
  assign n30380 = ~n70013 & n70018;
  assign n30381 = x165 & x180;
  assign n30382 = n30380 & n30381;
  assign n30383 = n30380 | n30381;
  assign n30384 = ~n30382 & n30383;
  assign n70019 = n29937 | n29939;
  assign n70020 = (n29937 & n55501) | (n29937 & n70019) | (n55501 & n70019);
  assign n55743 = n30384 & n70020;
  assign n70021 = n29500 | n29937;
  assign n70022 = (n29937 & n29939) | (n29937 & n70021) | (n29939 & n70021);
  assign n55744 = n30384 & n70022;
  assign n70023 = (n55743 & n55744) | (n55743 & n69741) | (n55744 & n69741);
  assign n70024 = (n55743 & n55744) | (n55743 & n69740) | (n55744 & n69740);
  assign n70025 = (n68982 & n70023) | (n68982 & n70024) | (n70023 & n70024);
  assign n55746 = n30384 | n70020;
  assign n55747 = n30384 | n70022;
  assign n70026 = (n55746 & n55747) | (n55746 & n69741) | (n55747 & n69741);
  assign n70027 = (n55746 & n55747) | (n55746 & n69740) | (n55747 & n69740);
  assign n70028 = (n68982 & n70026) | (n68982 & n70027) | (n70026 & n70027);
  assign n30387 = ~n70025 & n70028;
  assign n30388 = x164 & x181;
  assign n30389 = n30387 & n30388;
  assign n30390 = n30387 | n30388;
  assign n30391 = ~n30389 & n30390;
  assign n70029 = n29944 | n29946;
  assign n70030 = (n29944 & n55499) | (n29944 & n70029) | (n55499 & n70029);
  assign n55749 = n30391 & n70030;
  assign n70031 = n29507 | n29944;
  assign n70032 = (n29944 & n29946) | (n29944 & n70031) | (n29946 & n70031);
  assign n55750 = n30391 & n70032;
  assign n55751 = (n69736 & n55749) | (n69736 & n55750) | (n55749 & n55750);
  assign n55752 = n30391 | n70030;
  assign n55753 = n30391 | n70032;
  assign n55754 = (n69736 & n55752) | (n69736 & n55753) | (n55752 & n55753);
  assign n30394 = ~n55751 & n55754;
  assign n30395 = x163 & x182;
  assign n30396 = n30394 & n30395;
  assign n30397 = n30394 | n30395;
  assign n30398 = ~n30396 & n30397;
  assign n55755 = n29951 & n30398;
  assign n55756 = (n30398 & n69916) | (n30398 & n55755) | (n69916 & n55755);
  assign n55757 = n29951 | n30398;
  assign n55758 = n69916 | n55757;
  assign n30401 = ~n55756 & n55758;
  assign n30402 = x162 & x183;
  assign n30403 = n30401 & n30402;
  assign n30404 = n30401 | n30402;
  assign n30405 = ~n30403 & n30404;
  assign n55709 = n29958 | n29960;
  assign n55759 = n30405 & n55709;
  assign n55760 = n29958 & n30405;
  assign n55761 = (n69884 & n55759) | (n69884 & n55760) | (n55759 & n55760);
  assign n55762 = n30405 | n55709;
  assign n55763 = n29958 | n30405;
  assign n55764 = (n69884 & n55762) | (n69884 & n55763) | (n55762 & n55763);
  assign n30408 = ~n55761 & n55764;
  assign n30409 = x161 & x184;
  assign n30410 = n30408 & n30409;
  assign n30411 = n30408 | n30409;
  assign n30412 = ~n30410 & n30411;
  assign n55707 = n29965 | n55541;
  assign n70033 = n30412 & n55707;
  assign n69995 = n29528 | n29965;
  assign n69996 = (n29965 & n29967) | (n29965 & n69995) | (n29967 & n69995);
  assign n70034 = n30412 & n69996;
  assign n70035 = (n69730 & n70033) | (n69730 & n70034) | (n70033 & n70034);
  assign n70036 = n30412 | n55707;
  assign n70037 = n30412 | n69996;
  assign n70038 = (n69730 & n70036) | (n69730 & n70037) | (n70036 & n70037);
  assign n30415 = ~n70035 & n70038;
  assign n30416 = x160 & x185;
  assign n30417 = n30415 & n30416;
  assign n30418 = n30415 | n30416;
  assign n30419 = ~n30417 & n30418;
  assign n55704 = n29972 | n29974;
  assign n55765 = n30419 & n55704;
  assign n55766 = n29972 & n30419;
  assign n70039 = (n55489 & n55765) | (n55489 & n55766) | (n55765 & n55766);
  assign n70040 = (n55765 & n55766) | (n55765 & n69877) | (n55766 & n69877);
  assign n70041 = (n69578 & n70039) | (n69578 & n70040) | (n70039 & n70040);
  assign n55768 = n30419 | n55704;
  assign n55769 = n29972 | n30419;
  assign n70042 = (n55489 & n55768) | (n55489 & n55769) | (n55768 & n55769);
  assign n70043 = (n55768 & n55769) | (n55768 & n69877) | (n55769 & n69877);
  assign n70044 = (n69578 & n70042) | (n69578 & n70043) | (n70042 & n70043);
  assign n30422 = ~n70041 & n70044;
  assign n30423 = x159 & x186;
  assign n30424 = n30422 & n30423;
  assign n30425 = n30422 | n30423;
  assign n30426 = ~n30424 & n30425;
  assign n30427 = n69994 & n30426;
  assign n30428 = n69994 | n30426;
  assign n30429 = ~n30427 & n30428;
  assign n30430 = x158 & x187;
  assign n30431 = n30429 & n30430;
  assign n30432 = n30429 | n30430;
  assign n30433 = ~n30431 & n30432;
  assign n55699 = n29986 | n29988;
  assign n55771 = n30433 & n55699;
  assign n55772 = n29986 & n30433;
  assign n55773 = (n69875 & n55771) | (n69875 & n55772) | (n55771 & n55772);
  assign n55774 = n30433 | n55699;
  assign n55775 = n29986 | n30433;
  assign n55776 = (n69875 & n55774) | (n69875 & n55775) | (n55774 & n55775);
  assign n30436 = ~n55773 & n55776;
  assign n30437 = x157 & x188;
  assign n30438 = n30436 & n30437;
  assign n30439 = n30436 | n30437;
  assign n30440 = ~n30438 & n30439;
  assign n55777 = n29993 & n30440;
  assign n70045 = (n30440 & n55554) | (n30440 & n55777) | (n55554 & n55777);
  assign n70046 = (n30440 & n55553) | (n30440 & n55777) | (n55553 & n55777);
  assign n70047 = (n55282 & n70045) | (n55282 & n70046) | (n70045 & n70046);
  assign n55779 = n29993 | n30440;
  assign n70048 = n55554 | n55779;
  assign n70049 = n55553 | n55779;
  assign n70050 = (n55282 & n70048) | (n55282 & n70049) | (n70048 & n70049);
  assign n30443 = ~n70047 & n70050;
  assign n30444 = x156 & x189;
  assign n30445 = n30443 & n30444;
  assign n30446 = n30443 | n30444;
  assign n30447 = ~n30445 & n30446;
  assign n55697 = n30000 | n30002;
  assign n70051 = n30447 & n55697;
  assign n69986 = n29563 | n30000;
  assign n69987 = (n30000 & n30002) | (n30000 & n69986) | (n30002 & n69986);
  assign n70052 = n30447 & n69987;
  assign n70053 = (n55345 & n70051) | (n55345 & n70052) | (n70051 & n70052);
  assign n70054 = n30447 | n55697;
  assign n70055 = n30447 | n69987;
  assign n70056 = (n55345 & n70054) | (n55345 & n70055) | (n70054 & n70055);
  assign n30450 = ~n70053 & n70056;
  assign n30451 = x155 & x190;
  assign n30452 = n30450 & n30451;
  assign n30453 = n30450 | n30451;
  assign n30454 = ~n30452 & n30453;
  assign n55694 = n30007 | n30009;
  assign n55781 = n30454 & n55694;
  assign n55782 = n30007 & n30454;
  assign n55783 = (n69870 & n55781) | (n69870 & n55782) | (n55781 & n55782);
  assign n55784 = n30454 | n55694;
  assign n55785 = n30007 | n30454;
  assign n55786 = (n69870 & n55784) | (n69870 & n55785) | (n55784 & n55785);
  assign n30457 = ~n55783 & n55786;
  assign n30458 = x154 & x191;
  assign n30459 = n30457 & n30458;
  assign n30460 = n30457 | n30458;
  assign n30461 = ~n30459 & n30460;
  assign n55787 = n30014 & n30461;
  assign n70057 = (n30461 & n55564) | (n30461 & n55787) | (n55564 & n55787);
  assign n70058 = (n30461 & n55563) | (n30461 & n55787) | (n55563 & n55787);
  assign n70059 = (n55277 & n70057) | (n55277 & n70058) | (n70057 & n70058);
  assign n55789 = n30014 | n30461;
  assign n70060 = n55564 | n55789;
  assign n70061 = n55563 | n55789;
  assign n70062 = (n55277 & n70060) | (n55277 & n70061) | (n70060 & n70061);
  assign n30464 = ~n70059 & n70062;
  assign n30465 = x153 & x192;
  assign n30466 = n30464 & n30465;
  assign n30467 = n30464 | n30465;
  assign n30468 = ~n30466 & n30467;
  assign n55692 = n30021 | n30023;
  assign n70063 = n30468 & n55692;
  assign n69984 = n29584 | n30021;
  assign n69985 = (n30021 & n30023) | (n30021 & n69984) | (n30023 & n69984);
  assign n70064 = n30468 & n69985;
  assign n70065 = (n55355 & n70063) | (n55355 & n70064) | (n70063 & n70064);
  assign n70066 = n30468 | n55692;
  assign n70067 = n30468 | n69985;
  assign n70068 = (n55355 & n70066) | (n55355 & n70067) | (n70066 & n70067);
  assign n30471 = ~n70065 & n70068;
  assign n30472 = x152 & x193;
  assign n30473 = n30471 & n30472;
  assign n30474 = n30471 | n30472;
  assign n30475 = ~n30473 & n30474;
  assign n55689 = n30028 | n30030;
  assign n55791 = n30475 & n55689;
  assign n55792 = n30028 & n30475;
  assign n55793 = (n69865 & n55791) | (n69865 & n55792) | (n55791 & n55792);
  assign n55794 = n30475 | n55689;
  assign n55795 = n30028 | n30475;
  assign n55796 = (n69865 & n55794) | (n69865 & n55795) | (n55794 & n55795);
  assign n30478 = ~n55793 & n55796;
  assign n30479 = x151 & x194;
  assign n30480 = n30478 & n30479;
  assign n30481 = n30478 | n30479;
  assign n30482 = ~n30480 & n30481;
  assign n55797 = n30035 & n30482;
  assign n70069 = (n30482 & n55574) | (n30482 & n55797) | (n55574 & n55797);
  assign n70070 = (n30482 & n55573) | (n30482 & n55797) | (n55573 & n55797);
  assign n70071 = (n69717 & n70069) | (n69717 & n70070) | (n70069 & n70070);
  assign n55799 = n30035 | n30482;
  assign n70072 = n55574 | n55799;
  assign n70073 = n55573 | n55799;
  assign n70074 = (n69717 & n70072) | (n69717 & n70073) | (n70072 & n70073);
  assign n30485 = ~n70071 & n70074;
  assign n30486 = x150 & x195;
  assign n30487 = n30485 & n30486;
  assign n30488 = n30485 | n30486;
  assign n30489 = ~n30487 & n30488;
  assign n30490 = n69983 & n30489;
  assign n30491 = n69983 | n30489;
  assign n30492 = ~n30490 & n30491;
  assign n30493 = x149 & x196;
  assign n30494 = n30492 & n30493;
  assign n30495 = n30492 | n30493;
  assign n30496 = ~n30494 & n30495;
  assign n55684 = n30049 | n30051;
  assign n55801 = n30496 & n55684;
  assign n55802 = n30049 & n30496;
  assign n55803 = (n69860 & n55801) | (n69860 & n55802) | (n55801 & n55802);
  assign n55804 = n30496 | n55684;
  assign n55805 = n30049 | n30496;
  assign n55806 = (n69860 & n55804) | (n69860 & n55805) | (n55804 & n55805);
  assign n30499 = ~n55803 & n55806;
  assign n30500 = x148 & x197;
  assign n30501 = n30499 & n30500;
  assign n30502 = n30499 | n30500;
  assign n30503 = ~n30501 & n30502;
  assign n55807 = n30056 & n30503;
  assign n70075 = (n30503 & n55584) | (n30503 & n55807) | (n55584 & n55807);
  assign n70076 = (n30503 & n55583) | (n30503 & n55807) | (n55583 & n55807);
  assign n70077 = (n69712 & n70075) | (n69712 & n70076) | (n70075 & n70076);
  assign n55809 = n30056 | n30503;
  assign n70078 = n55584 | n55809;
  assign n70079 = n55583 | n55809;
  assign n70080 = (n69712 & n70078) | (n69712 & n70079) | (n70078 & n70079);
  assign n30506 = ~n70077 & n70080;
  assign n30507 = x147 & x198;
  assign n30508 = n30506 & n30507;
  assign n30509 = n30506 | n30507;
  assign n30510 = ~n30508 & n30509;
  assign n30511 = n69978 & n30510;
  assign n30512 = n69978 | n30510;
  assign n30513 = ~n30511 & n30512;
  assign n30514 = x146 & x199;
  assign n30515 = n30513 & n30514;
  assign n30516 = n30513 | n30514;
  assign n30517 = ~n30515 & n30516;
  assign n55679 = n30070 | n30072;
  assign n55811 = n30517 & n55679;
  assign n55812 = n30070 & n30517;
  assign n55813 = (n55465 & n55811) | (n55465 & n55812) | (n55811 & n55812);
  assign n55814 = n30517 | n55679;
  assign n55815 = n30070 | n30517;
  assign n55816 = (n55465 & n55814) | (n55465 & n55815) | (n55814 & n55815);
  assign n30520 = ~n55813 & n55816;
  assign n30521 = x145 & x200;
  assign n30522 = n30520 & n30521;
  assign n30523 = n30520 | n30521;
  assign n30524 = ~n30522 & n30523;
  assign n55817 = n30077 & n30524;
  assign n55818 = (n30524 & n69954) | (n30524 & n55817) | (n69954 & n55817);
  assign n55819 = n30077 | n30524;
  assign n55820 = n69954 | n55819;
  assign n30527 = ~n55818 & n55820;
  assign n30528 = x144 & x201;
  assign n30529 = n30527 & n30528;
  assign n30530 = n30527 | n30528;
  assign n30531 = ~n30529 & n30530;
  assign n55821 = n30084 & n30531;
  assign n55822 = (n30531 & n55598) | (n30531 & n55821) | (n55598 & n55821);
  assign n55823 = n30084 | n30531;
  assign n55824 = n55598 | n55823;
  assign n30534 = ~n55822 & n55824;
  assign n30535 = x143 & x202;
  assign n30536 = n30534 & n30535;
  assign n30537 = n30534 | n30535;
  assign n30538 = ~n30536 & n30537;
  assign n55825 = n30091 & n30538;
  assign n55826 = (n30538 & n55602) | (n30538 & n55825) | (n55602 & n55825);
  assign n55827 = n30091 | n30538;
  assign n55828 = n55602 | n55827;
  assign n30541 = ~n55826 & n55828;
  assign n30542 = x142 & x203;
  assign n30543 = n30541 & n30542;
  assign n30544 = n30541 | n30542;
  assign n30545 = ~n30543 & n30544;
  assign n55829 = n30098 & n30545;
  assign n55830 = (n30545 & n55606) | (n30545 & n55829) | (n55606 & n55829);
  assign n55831 = n30098 | n30545;
  assign n55832 = n55606 | n55831;
  assign n30548 = ~n55830 & n55832;
  assign n30549 = x141 & x204;
  assign n30550 = n30548 & n30549;
  assign n30551 = n30548 | n30549;
  assign n30552 = ~n30550 & n30551;
  assign n55833 = n30105 & n30552;
  assign n55834 = (n30552 & n55610) | (n30552 & n55833) | (n55610 & n55833);
  assign n55835 = n30105 | n30552;
  assign n55836 = n55610 | n55835;
  assign n30555 = ~n55834 & n55836;
  assign n30556 = x140 & x205;
  assign n30557 = n30555 & n30556;
  assign n30558 = n30555 | n30556;
  assign n30559 = ~n30557 & n30558;
  assign n55837 = n30112 & n30559;
  assign n55838 = (n30559 & n55614) | (n30559 & n55837) | (n55614 & n55837);
  assign n55839 = n30112 | n30559;
  assign n55840 = n55614 | n55839;
  assign n30562 = ~n55838 & n55840;
  assign n30563 = x139 & x206;
  assign n30564 = n30562 & n30563;
  assign n30565 = n30562 | n30563;
  assign n30566 = ~n30564 & n30565;
  assign n55841 = n30119 & n30566;
  assign n55842 = (n30566 & n55618) | (n30566 & n55841) | (n55618 & n55841);
  assign n55843 = n30119 | n30566;
  assign n55844 = n55618 | n55843;
  assign n30569 = ~n55842 & n55844;
  assign n30570 = x138 & x207;
  assign n30571 = n30569 & n30570;
  assign n30572 = n30569 | n30570;
  assign n30573 = ~n30571 & n30572;
  assign n55845 = n30126 & n30573;
  assign n55846 = (n30573 & n55622) | (n30573 & n55845) | (n55622 & n55845);
  assign n55847 = n30126 | n30573;
  assign n55848 = n55622 | n55847;
  assign n30576 = ~n55846 & n55848;
  assign n30577 = x137 & x208;
  assign n30578 = n30576 & n30577;
  assign n30579 = n30576 | n30577;
  assign n30580 = ~n30578 & n30579;
  assign n55849 = n30133 & n30580;
  assign n55850 = (n30580 & n55626) | (n30580 & n55849) | (n55626 & n55849);
  assign n55851 = n30133 | n30580;
  assign n55852 = n55626 | n55851;
  assign n30583 = ~n55850 & n55852;
  assign n30584 = x136 & x209;
  assign n30585 = n30583 & n30584;
  assign n30586 = n30583 | n30584;
  assign n30587 = ~n30585 & n30586;
  assign n55853 = n30140 & n30587;
  assign n55854 = (n30587 & n55630) | (n30587 & n55853) | (n55630 & n55853);
  assign n55855 = n30140 | n30587;
  assign n55856 = n55630 | n55855;
  assign n30590 = ~n55854 & n55856;
  assign n30591 = x135 & x210;
  assign n30592 = n30590 & n30591;
  assign n30593 = n30590 | n30591;
  assign n30594 = ~n30592 & n30593;
  assign n55857 = n30147 & n30594;
  assign n55858 = (n30594 & n55634) | (n30594 & n55857) | (n55634 & n55857);
  assign n55859 = n30147 | n30594;
  assign n55860 = n55634 | n55859;
  assign n30597 = ~n55858 & n55860;
  assign n30598 = x134 & x211;
  assign n30599 = n30597 & n30598;
  assign n30600 = n30597 | n30598;
  assign n30601 = ~n30599 & n30600;
  assign n55861 = n30154 & n30601;
  assign n55862 = (n30601 & n55638) | (n30601 & n55861) | (n55638 & n55861);
  assign n55863 = n30154 | n30601;
  assign n55864 = n55638 | n55863;
  assign n30604 = ~n55862 & n55864;
  assign n30605 = x133 & x212;
  assign n30606 = n30604 & n30605;
  assign n30607 = n30604 | n30605;
  assign n30608 = ~n30606 & n30607;
  assign n55865 = n30161 & n30608;
  assign n55866 = (n30608 & n55642) | (n30608 & n55865) | (n55642 & n55865);
  assign n55867 = n30161 | n30608;
  assign n55868 = n55642 | n55867;
  assign n30611 = ~n55866 & n55868;
  assign n30612 = x132 & x213;
  assign n30613 = n30611 & n30612;
  assign n30614 = n30611 | n30612;
  assign n30615 = ~n30613 & n30614;
  assign n55869 = n30168 & n30615;
  assign n55870 = (n30615 & n55646) | (n30615 & n55869) | (n55646 & n55869);
  assign n55871 = n30168 | n30615;
  assign n55872 = n55646 | n55871;
  assign n30618 = ~n55870 & n55872;
  assign n30619 = x131 & x214;
  assign n30620 = n30618 & n30619;
  assign n30621 = n30618 | n30619;
  assign n30622 = ~n30620 & n30621;
  assign n55873 = n30175 & n30622;
  assign n55874 = (n30622 & n55650) | (n30622 & n55873) | (n55650 & n55873);
  assign n55875 = n30175 | n30622;
  assign n55876 = n55650 | n55875;
  assign n30625 = ~n55874 & n55876;
  assign n30626 = x130 & x215;
  assign n30627 = n30625 & n30626;
  assign n30628 = n30625 | n30626;
  assign n30629 = ~n30627 & n30628;
  assign n55877 = n30182 & n30629;
  assign n55878 = (n30629 & n55655) | (n30629 & n55877) | (n55655 & n55877);
  assign n55879 = n30182 | n30629;
  assign n55880 = n55655 | n55879;
  assign n30632 = ~n55878 & n55880;
  assign n30633 = x129 & x216;
  assign n30634 = n30632 & n30633;
  assign n30635 = n30632 | n30633;
  assign n30636 = ~n30634 & n30635;
  assign n55677 = n30189 | n30191;
  assign n55881 = n30636 & n55677;
  assign n55882 = n30189 & n30636;
  assign n55883 = (n55460 & n55881) | (n55460 & n55882) | (n55881 & n55882);
  assign n55884 = n30636 | n55677;
  assign n55885 = n30189 | n30636;
  assign n55886 = (n55460 & n55884) | (n55460 & n55885) | (n55884 & n55885);
  assign n30639 = ~n55883 & n55886;
  assign n30640 = x128 & x217;
  assign n30641 = n30639 & n30640;
  assign n30642 = n30639 | n30640;
  assign n30643 = ~n30641 & n30642;
  assign n55675 = n30196 | n30198;
  assign n70081 = n30643 & n55675;
  assign n70082 = n30196 & n30643;
  assign n70083 = (n55458 & n70081) | (n55458 & n70082) | (n70081 & n70082);
  assign n70084 = n30643 | n55675;
  assign n70085 = n30196 | n30643;
  assign n70086 = (n55458 & n70084) | (n55458 & n70085) | (n70084 & n70085);
  assign n30646 = ~n70083 & n70086;
  assign n30647 = x127 & x218;
  assign n30648 = n30646 & n30647;
  assign n30649 = n30646 | n30647;
  assign n30650 = ~n30648 & n30649;
  assign n55673 = n30203 | n30205;
  assign n70087 = n30650 & n55673;
  assign n70088 = n30203 & n30650;
  assign n70089 = (n55456 & n70087) | (n55456 & n70088) | (n70087 & n70088);
  assign n70090 = n30650 | n55673;
  assign n70091 = n30203 | n30650;
  assign n70092 = (n55456 & n70090) | (n55456 & n70091) | (n70090 & n70091);
  assign n30653 = ~n70089 & n70092;
  assign n30654 = x126 & x219;
  assign n30655 = n30653 & n30654;
  assign n30656 = n30653 | n30654;
  assign n30657 = ~n30655 & n30656;
  assign n30658 = n55672 & n30657;
  assign n30659 = n55672 | n30657;
  assign n30660 = ~n30658 & n30659;
  assign n30661 = x125 & x220;
  assign n30662 = n30660 & n30661;
  assign n30663 = n30660 | n30661;
  assign n30664 = ~n30662 & n30663;
  assign n30665 = n55670 & n30664;
  assign n30666 = n55670 | n30664;
  assign n30667 = ~n30665 & n30666;
  assign n30668 = x124 & x221;
  assign n30669 = n30667 & n30668;
  assign n30670 = n30667 | n30668;
  assign n30671 = ~n30669 & n30670;
  assign n30672 = n55668 & n30671;
  assign n30673 = n55668 | n30671;
  assign n30674 = ~n30672 & n30673;
  assign n30675 = x123 & x222;
  assign n30676 = n30674 & n30675;
  assign n30677 = n30674 | n30675;
  assign n30678 = ~n30676 & n30677;
  assign n30679 = n30313 & n30678;
  assign n30680 = n30313 | n30678;
  assign n30681 = ~n30679 & n30680;
  assign n30682 = x122 & x223;
  assign n30683 = n30681 & n30682;
  assign n30684 = n30681 | n30682;
  assign n30685 = ~n30683 & n30684;
  assign n30686 = n30312 & n30685;
  assign n30687 = n30312 | n30685;
  assign n30688 = ~n30686 & n30687;
  assign n30689 = x121 & x224;
  assign n30690 = n30688 & n30689;
  assign n30691 = n30688 | n30689;
  assign n30692 = ~n30690 & n30691;
  assign n30693 = n30311 & n30692;
  assign n30694 = n30311 | n30692;
  assign n30695 = ~n30693 & n30694;
  assign n30696 = x120 & x225;
  assign n30697 = n30695 & n30696;
  assign n30698 = n30695 | n30696;
  assign n30699 = ~n30697 & n30698;
  assign n30700 = n30310 & n30699;
  assign n30701 = n30310 | n30699;
  assign n30702 = ~n30700 & n30701;
  assign n30703 = x119 & x226;
  assign n30704 = n30702 & n30703;
  assign n30705 = n30702 | n30703;
  assign n30706 = ~n30704 & n30705;
  assign n30707 = n30309 & n30706;
  assign n30708 = n30309 | n30706;
  assign n30709 = ~n30707 & n30708;
  assign n30710 = x118 & x227;
  assign n30711 = n30709 & n30710;
  assign n30712 = n30709 | n30710;
  assign n30713 = ~n30711 & n30712;
  assign n30714 = n69973 & n30713;
  assign n30715 = n69973 | n30713;
  assign n30716 = ~n30714 & n30715;
  assign n30717 = x117 & x228;
  assign n30718 = n30716 & n30717;
  assign n30719 = n30716 | n30717;
  assign n30720 = ~n30718 & n30719;
  assign n30721 = n55666 & n30720;
  assign n30722 = n55666 | n30720;
  assign n30723 = ~n30721 & n30722;
  assign n30724 = x116 & x229;
  assign n30725 = n30723 & n30724;
  assign n30726 = n30723 | n30724;
  assign n30727 = ~n30725 & n30726;
  assign n30728 = n55664 & n30727;
  assign n30729 = n55664 | n30727;
  assign n30730 = ~n30728 & n30729;
  assign n30731 = x115 & x230;
  assign n30732 = n30730 & n30731;
  assign n30733 = n30730 | n30731;
  assign n30734 = ~n30732 & n30733;
  assign n30735 = n55662 & n30734;
  assign n30736 = n55662 | n30734;
  assign n30737 = ~n30735 & n30736;
  assign n30738 = x114 & x231;
  assign n30739 = n30737 & n30738;
  assign n30740 = n30737 | n30738;
  assign n30741 = ~n30739 & n30740;
  assign n30742 = n55660 & n30741;
  assign n30743 = n55660 | n30741;
  assign n30744 = ~n30742 & n30743;
  assign n30745 = x113 & x232;
  assign n30746 = n30744 & n30745;
  assign n30747 = n30744 | n30745;
  assign n30748 = ~n30746 & n30747;
  assign n30749 = n30301 & n30748;
  assign n30750 = n30301 | n30748;
  assign n30751 = ~n30749 & n30750;
  assign n30752 = x112 & x233;
  assign n30753 = n30751 & n30752;
  assign n30754 = n30751 | n30752;
  assign n30755 = ~n30753 & n30754;
  assign n70093 = n30301 | n30745;
  assign n70094 = (n30301 & n30744) | (n30301 & n70093) | (n30744 & n70093);
  assign n55888 = (n30746 & n30748) | (n30746 & n70094) | (n30748 & n70094);
  assign n55889 = n30739 | n55660;
  assign n55890 = (n30739 & n30741) | (n30739 & n55889) | (n30741 & n55889);
  assign n55891 = n30732 | n55662;
  assign n55892 = (n30732 & n30734) | (n30732 & n55891) | (n30734 & n55891);
  assign n55893 = n30725 | n55664;
  assign n55894 = (n30725 & n30727) | (n30725 & n55893) | (n30727 & n55893);
  assign n55895 = n30718 | n55666;
  assign n55896 = (n30718 & n30720) | (n30718 & n55895) | (n30720 & n55895);
  assign n70095 = n30711 | n69973;
  assign n70096 = (n30711 & n30713) | (n30711 & n70095) | (n30713 & n70095);
  assign n30762 = n30704 | n30707;
  assign n30763 = n30697 | n30700;
  assign n30764 = n30690 | n30693;
  assign n30765 = n30683 | n30686;
  assign n55897 = n30676 | n30678;
  assign n55898 = (n30313 & n30676) | (n30313 & n55897) | (n30676 & n55897);
  assign n55899 = n30669 | n30671;
  assign n55900 = (n30669 & n55668) | (n30669 & n55899) | (n55668 & n55899);
  assign n55901 = n30662 | n30664;
  assign n55902 = (n30662 & n55670) | (n30662 & n55901) | (n55670 & n55901);
  assign n55674 = (n30203 & n55456) | (n30203 & n55673) | (n55456 & n55673);
  assign n55676 = (n30196 & n55458) | (n30196 & n55675) | (n55458 & n55675);
  assign n55915 = n30501 | n30503;
  assign n70099 = n30056 | n30501;
  assign n70100 = (n30501 & n30503) | (n30501 & n70099) | (n30503 & n70099);
  assign n70101 = (n55584 & n55915) | (n55584 & n70100) | (n55915 & n70100);
  assign n70102 = (n55583 & n55915) | (n55583 & n70100) | (n55915 & n70100);
  assign n70103 = (n69712 & n70101) | (n69712 & n70102) | (n70101 & n70102);
  assign n55920 = n30480 | n30482;
  assign n70104 = n30035 | n30480;
  assign n70105 = (n30480 & n30482) | (n30480 & n70104) | (n30482 & n70104);
  assign n70106 = (n55574 & n55920) | (n55574 & n70105) | (n55920 & n70105);
  assign n70107 = (n55573 & n55920) | (n55573 & n70105) | (n55920 & n70105);
  assign n70108 = (n69717 & n70106) | (n69717 & n70107) | (n70106 & n70107);
  assign n55693 = (n55355 & n69985) | (n55355 & n55692) | (n69985 & n55692);
  assign n55925 = n30459 | n30461;
  assign n70109 = n30014 | n30459;
  assign n70110 = (n30459 & n30461) | (n30459 & n70109) | (n30461 & n70109);
  assign n70111 = (n55564 & n55925) | (n55564 & n70110) | (n55925 & n70110);
  assign n70112 = (n55563 & n55925) | (n55563 & n70110) | (n55925 & n70110);
  assign n70113 = (n55277 & n70111) | (n55277 & n70112) | (n70111 & n70112);
  assign n55698 = (n55345 & n69987) | (n55345 & n55697) | (n69987 & n55697);
  assign n55930 = n30438 | n30440;
  assign n70114 = n29993 | n30438;
  assign n70115 = (n30438 & n30440) | (n30438 & n70114) | (n30440 & n70114);
  assign n70116 = (n55554 & n55930) | (n55554 & n70115) | (n55930 & n70115);
  assign n70117 = (n55553 & n55930) | (n55553 & n70115) | (n55930 & n70115);
  assign n70118 = (n55282 & n70116) | (n55282 & n70117) | (n70116 & n70117);
  assign n70119 = n29986 | n30431;
  assign n70120 = (n30431 & n30433) | (n30431 & n70119) | (n30433 & n70119);
  assign n55933 = n30431 | n55771;
  assign n55934 = (n69875 & n70120) | (n69875 & n55933) | (n70120 & n55933);
  assign n70121 = n29972 | n30417;
  assign n70122 = (n30417 & n30419) | (n30417 & n70121) | (n30419 & n70121);
  assign n70123 = n30417 | n30419;
  assign n70124 = (n30417 & n55704) | (n30417 & n70123) | (n55704 & n70123);
  assign n70125 = (n55489 & n70122) | (n55489 & n70124) | (n70122 & n70124);
  assign n70126 = (n69877 & n70122) | (n69877 & n70124) | (n70122 & n70124);
  assign n70127 = (n69578 & n70125) | (n69578 & n70126) | (n70125 & n70126);
  assign n70128 = n30382 | n30384;
  assign n70129 = (n30382 & n70020) | (n30382 & n70128) | (n70020 & n70128);
  assign n70130 = (n30382 & n70022) | (n30382 & n70128) | (n70022 & n70128);
  assign n70131 = (n69741 & n70129) | (n69741 & n70130) | (n70129 & n70130);
  assign n70132 = (n69740 & n70129) | (n69740 & n70130) | (n70129 & n70130);
  assign n70133 = (n68982 & n70131) | (n68982 & n70132) | (n70131 & n70132);
  assign n30812 = x170 & x176;
  assign n30813 = x169 & x177;
  assign n30814 = n30812 & n30813;
  assign n30815 = n30812 | n30813;
  assign n30816 = ~n30814 & n30815;
  assign n70134 = n30361 | n30363;
  assign n70139 = (n30361 & n70000) | (n30361 & n70134) | (n70000 & n70134);
  assign n55958 = n30816 & n70139;
  assign n70136 = n30816 & n70134;
  assign n70137 = n30361 & n30816;
  assign n70138 = (n69998 & n70136) | (n69998 & n70137) | (n70136 & n70137);
  assign n70140 = (n55958 & n69747) | (n55958 & n70138) | (n69747 & n70138);
  assign n70141 = (n55958 & n69746) | (n55958 & n70138) | (n69746 & n70138);
  assign n70142 = (n68195 & n70140) | (n68195 & n70141) | (n70140 & n70141);
  assign n55961 = n30816 | n70139;
  assign n70143 = n30816 | n70134;
  assign n70144 = n30361 | n30816;
  assign n70145 = (n69998 & n70143) | (n69998 & n70144) | (n70143 & n70144);
  assign n70146 = (n55961 & n69747) | (n55961 & n70145) | (n69747 & n70145);
  assign n70147 = (n55961 & n69746) | (n55961 & n70145) | (n69746 & n70145);
  assign n70148 = (n68195 & n70146) | (n68195 & n70147) | (n70146 & n70147);
  assign n30819 = ~n70142 & n70148;
  assign n30820 = x168 & x178;
  assign n30821 = n30819 & n30820;
  assign n30822 = n30819 | n30820;
  assign n30823 = ~n30821 & n30822;
  assign n70149 = n30368 | n30370;
  assign n70150 = (n30368 & n55720) | (n30368 & n70149) | (n55720 & n70149);
  assign n55963 = n30823 & n70150;
  assign n70151 = n29923 | n30368;
  assign n70152 = (n30368 & n30370) | (n30368 & n70151) | (n30370 & n70151);
  assign n55964 = n30823 & n70152;
  assign n55965 = (n69887 & n55963) | (n69887 & n55964) | (n55963 & n55964);
  assign n55966 = n30823 | n70150;
  assign n55967 = n30823 | n70152;
  assign n55968 = (n69887 & n55966) | (n69887 & n55967) | (n55966 & n55967);
  assign n30826 = ~n55965 & n55968;
  assign n30827 = x167 & x179;
  assign n30828 = n30826 & n30827;
  assign n30829 = n30826 | n30827;
  assign n30830 = ~n30828 & n30829;
  assign n55969 = n30375 & n30830;
  assign n55970 = (n30830 & n70013) | (n30830 & n55969) | (n70013 & n55969);
  assign n55971 = n30375 | n30830;
  assign n55972 = n70013 | n55971;
  assign n30833 = ~n55970 & n55972;
  assign n30834 = x166 & x180;
  assign n30835 = n30833 & n30834;
  assign n30836 = n30833 | n30834;
  assign n30837 = ~n30835 & n30836;
  assign n30838 = n70133 & n30837;
  assign n30839 = n70133 | n30837;
  assign n30840 = ~n30838 & n30839;
  assign n30841 = x165 & x181;
  assign n30842 = n30840 & n30841;
  assign n30843 = n30840 | n30841;
  assign n30844 = ~n30842 & n30843;
  assign n55973 = n30389 & n30844;
  assign n70153 = (n30844 & n55749) | (n30844 & n55973) | (n55749 & n55973);
  assign n70154 = (n30844 & n55750) | (n30844 & n55973) | (n55750 & n55973);
  assign n70155 = (n69736 & n70153) | (n69736 & n70154) | (n70153 & n70154);
  assign n55975 = n30389 | n30844;
  assign n70156 = n55749 | n55975;
  assign n70157 = n55750 | n55975;
  assign n70158 = (n69736 & n70156) | (n69736 & n70157) | (n70156 & n70157);
  assign n30847 = ~n70155 & n70158;
  assign n30848 = x164 & x182;
  assign n30849 = n30847 & n30848;
  assign n30850 = n30847 | n30848;
  assign n30851 = ~n30849 & n30850;
  assign n70159 = n29951 | n30396;
  assign n70160 = (n30396 & n30398) | (n30396 & n70159) | (n30398 & n70159);
  assign n55977 = n30851 & n70160;
  assign n55946 = n30396 | n30398;
  assign n55978 = n30851 & n55946;
  assign n55979 = (n69916 & n55977) | (n69916 & n55978) | (n55977 & n55978);
  assign n55980 = n30851 | n70160;
  assign n55981 = n30851 | n55946;
  assign n55982 = (n69916 & n55980) | (n69916 & n55981) | (n55980 & n55981);
  assign n30854 = ~n55979 & n55982;
  assign n30855 = x163 & x183;
  assign n30856 = n30854 & n30855;
  assign n30857 = n30854 | n30855;
  assign n30858 = ~n30856 & n30857;
  assign n70161 = n30403 & n30858;
  assign n70162 = (n30858 & n55759) | (n30858 & n70161) | (n55759 & n70161);
  assign n70163 = n29958 | n30403;
  assign n70164 = (n30403 & n30405) | (n30403 & n70163) | (n30405 & n70163);
  assign n55984 = n30858 & n70164;
  assign n55985 = (n69884 & n70162) | (n69884 & n55984) | (n70162 & n55984);
  assign n70165 = n30403 | n30858;
  assign n70166 = n55759 | n70165;
  assign n55987 = n30858 | n70164;
  assign n55988 = (n69884 & n70166) | (n69884 & n55987) | (n70166 & n55987);
  assign n30861 = ~n55985 & n55988;
  assign n30862 = x162 & x184;
  assign n30863 = n30861 & n30862;
  assign n30864 = n30861 | n30862;
  assign n30865 = ~n30863 & n30864;
  assign n55940 = n30410 | n30412;
  assign n55989 = n30865 & n55940;
  assign n55990 = n30410 & n30865;
  assign n70167 = (n55707 & n55989) | (n55707 & n55990) | (n55989 & n55990);
  assign n70168 = (n55989 & n55990) | (n55989 & n69996) | (n55990 & n69996);
  assign n70169 = (n69730 & n70167) | (n69730 & n70168) | (n70167 & n70168);
  assign n55992 = n30865 | n55940;
  assign n55993 = n30410 | n30865;
  assign n70170 = (n55707 & n55992) | (n55707 & n55993) | (n55992 & n55993);
  assign n70171 = (n55992 & n55993) | (n55992 & n69996) | (n55993 & n69996);
  assign n70172 = (n69730 & n70170) | (n69730 & n70171) | (n70170 & n70171);
  assign n30868 = ~n70169 & n70172;
  assign n30869 = x161 & x185;
  assign n30870 = n30868 & n30869;
  assign n30871 = n30868 | n30869;
  assign n30872 = ~n30870 & n30871;
  assign n30873 = n70127 & n30872;
  assign n30874 = n70127 | n30872;
  assign n30875 = ~n30873 & n30874;
  assign n30876 = x160 & x186;
  assign n30877 = n30875 & n30876;
  assign n30878 = n30875 | n30876;
  assign n30879 = ~n30877 & n30878;
  assign n55935 = n30424 | n30426;
  assign n55995 = n30879 & n55935;
  assign n55996 = n30424 & n30879;
  assign n55997 = (n69994 & n55995) | (n69994 & n55996) | (n55995 & n55996);
  assign n55998 = n30879 | n55935;
  assign n55999 = n30424 | n30879;
  assign n56000 = (n69994 & n55998) | (n69994 & n55999) | (n55998 & n55999);
  assign n30882 = ~n55997 & n56000;
  assign n30883 = x159 & x187;
  assign n30884 = n30882 & n30883;
  assign n30885 = n30882 | n30883;
  assign n30886 = ~n30884 & n30885;
  assign n30887 = n55934 & n30886;
  assign n30888 = n55934 | n30886;
  assign n30889 = ~n30887 & n30888;
  assign n30890 = x158 & x188;
  assign n30891 = n30889 & n30890;
  assign n30892 = n30889 | n30890;
  assign n30893 = ~n30891 & n30892;
  assign n30894 = n70118 & n30893;
  assign n30895 = n70118 | n30893;
  assign n30896 = ~n30894 & n30895;
  assign n30897 = x157 & x189;
  assign n30898 = n30896 & n30897;
  assign n30899 = n30896 | n30897;
  assign n30900 = ~n30898 & n30899;
  assign n55927 = n30445 | n30447;
  assign n56001 = n30900 & n55927;
  assign n56002 = n30445 & n30900;
  assign n56003 = (n55698 & n56001) | (n55698 & n56002) | (n56001 & n56002);
  assign n56004 = n30900 | n55927;
  assign n56005 = n30445 | n30900;
  assign n56006 = (n55698 & n56004) | (n55698 & n56005) | (n56004 & n56005);
  assign n30903 = ~n56003 & n56006;
  assign n30904 = x156 & x190;
  assign n30905 = n30903 & n30904;
  assign n30906 = n30903 | n30904;
  assign n30907 = ~n30905 & n30906;
  assign n56007 = n30452 & n30907;
  assign n56008 = (n30907 & n55783) | (n30907 & n56007) | (n55783 & n56007);
  assign n56009 = n30452 | n30907;
  assign n56010 = n55783 | n56009;
  assign n30910 = ~n56008 & n56010;
  assign n30911 = x155 & x191;
  assign n30912 = n30910 & n30911;
  assign n30913 = n30910 | n30911;
  assign n30914 = ~n30912 & n30913;
  assign n30915 = n70113 & n30914;
  assign n30916 = n70113 | n30914;
  assign n30917 = ~n30915 & n30916;
  assign n30918 = x154 & x192;
  assign n30919 = n30917 & n30918;
  assign n30920 = n30917 | n30918;
  assign n30921 = ~n30919 & n30920;
  assign n55922 = n30466 | n30468;
  assign n56011 = n30921 & n55922;
  assign n56012 = n30466 & n30921;
  assign n56013 = (n55693 & n56011) | (n55693 & n56012) | (n56011 & n56012);
  assign n56014 = n30921 | n55922;
  assign n56015 = n30466 | n30921;
  assign n56016 = (n55693 & n56014) | (n55693 & n56015) | (n56014 & n56015);
  assign n30924 = ~n56013 & n56016;
  assign n30925 = x153 & x193;
  assign n30926 = n30924 & n30925;
  assign n30927 = n30924 | n30925;
  assign n30928 = ~n30926 & n30927;
  assign n56017 = n30473 & n30928;
  assign n56018 = (n30928 & n55793) | (n30928 & n56017) | (n55793 & n56017);
  assign n56019 = n30473 | n30928;
  assign n56020 = n55793 | n56019;
  assign n30931 = ~n56018 & n56020;
  assign n30932 = x152 & x194;
  assign n30933 = n30931 & n30932;
  assign n30934 = n30931 | n30932;
  assign n30935 = ~n30933 & n30934;
  assign n30936 = n70108 & n30935;
  assign n30937 = n70108 | n30935;
  assign n30938 = ~n30936 & n30937;
  assign n30939 = x151 & x195;
  assign n30940 = n30938 & n30939;
  assign n30941 = n30938 | n30939;
  assign n30942 = ~n30940 & n30941;
  assign n55917 = n30487 | n30489;
  assign n56021 = n30942 & n55917;
  assign n56022 = n30487 & n30942;
  assign n56023 = (n69983 & n56021) | (n69983 & n56022) | (n56021 & n56022);
  assign n56024 = n30942 | n55917;
  assign n56025 = n30487 | n30942;
  assign n56026 = (n69983 & n56024) | (n69983 & n56025) | (n56024 & n56025);
  assign n30945 = ~n56023 & n56026;
  assign n30946 = x150 & x196;
  assign n30947 = n30945 & n30946;
  assign n30948 = n30945 | n30946;
  assign n30949 = ~n30947 & n30948;
  assign n56027 = n30494 & n30949;
  assign n70173 = (n30949 & n55802) | (n30949 & n56027) | (n55802 & n56027);
  assign n70174 = (n30949 & n55801) | (n30949 & n56027) | (n55801 & n56027);
  assign n70175 = (n69860 & n70173) | (n69860 & n70174) | (n70173 & n70174);
  assign n56029 = n30494 | n30949;
  assign n70176 = n55802 | n56029;
  assign n70177 = n55801 | n56029;
  assign n70178 = (n69860 & n70176) | (n69860 & n70177) | (n70176 & n70177);
  assign n30952 = ~n70175 & n70178;
  assign n30953 = x149 & x197;
  assign n30954 = n30952 & n30953;
  assign n30955 = n30952 | n30953;
  assign n30956 = ~n30954 & n30955;
  assign n30957 = n70103 & n30956;
  assign n30958 = n70103 | n30956;
  assign n30959 = ~n30957 & n30958;
  assign n30960 = x148 & x198;
  assign n30961 = n30959 & n30960;
  assign n30962 = n30959 | n30960;
  assign n30963 = ~n30961 & n30962;
  assign n55912 = n30508 | n30510;
  assign n56031 = n30963 & n55912;
  assign n56032 = n30508 & n30963;
  assign n56033 = (n69978 & n56031) | (n69978 & n56032) | (n56031 & n56032);
  assign n56034 = n30963 | n55912;
  assign n56035 = n30508 | n30963;
  assign n56036 = (n69978 & n56034) | (n69978 & n56035) | (n56034 & n56035);
  assign n30966 = ~n56033 & n56036;
  assign n30967 = x147 & x199;
  assign n30968 = n30966 & n30967;
  assign n30969 = n30966 | n30967;
  assign n30970 = ~n30968 & n30969;
  assign n56037 = n30515 & n30970;
  assign n70179 = (n30970 & n55812) | (n30970 & n56037) | (n55812 & n56037);
  assign n70180 = (n30970 & n55811) | (n30970 & n56037) | (n55811 & n56037);
  assign n70181 = (n55465 & n70179) | (n55465 & n70180) | (n70179 & n70180);
  assign n56039 = n30515 | n30970;
  assign n70182 = n55812 | n56039;
  assign n70183 = n55811 | n56039;
  assign n70184 = (n55465 & n70182) | (n55465 & n70183) | (n70182 & n70183);
  assign n30973 = ~n70181 & n70184;
  assign n30974 = x146 & x200;
  assign n30975 = n30973 & n30974;
  assign n30976 = n30973 | n30974;
  assign n30977 = ~n30975 & n30976;
  assign n55910 = n30522 | n30524;
  assign n70185 = n30977 & n55910;
  assign n70097 = n30077 | n30522;
  assign n70098 = (n30522 & n30524) | (n30522 & n70097) | (n30524 & n70097);
  assign n70186 = n30977 & n70098;
  assign n70187 = (n69954 & n70185) | (n69954 & n70186) | (n70185 & n70186);
  assign n70188 = n30977 | n55910;
  assign n70189 = n30977 | n70098;
  assign n70190 = (n69954 & n70188) | (n69954 & n70189) | (n70188 & n70189);
  assign n30980 = ~n70187 & n70190;
  assign n30981 = x145 & x201;
  assign n30982 = n30980 & n30981;
  assign n30983 = n30980 | n30981;
  assign n30984 = ~n30982 & n30983;
  assign n56041 = n30529 & n30984;
  assign n70191 = (n30984 & n55821) | (n30984 & n56041) | (n55821 & n56041);
  assign n70192 = (n30531 & n30984) | (n30531 & n56041) | (n30984 & n56041);
  assign n70193 = (n55598 & n70191) | (n55598 & n70192) | (n70191 & n70192);
  assign n56043 = n30529 | n30984;
  assign n70194 = n55821 | n56043;
  assign n70195 = n30531 | n56043;
  assign n70196 = (n55598 & n70194) | (n55598 & n70195) | (n70194 & n70195);
  assign n30987 = ~n70193 & n70196;
  assign n30988 = x144 & x202;
  assign n30989 = n30987 & n30988;
  assign n30990 = n30987 | n30988;
  assign n30991 = ~n30989 & n30990;
  assign n56045 = n30536 & n30991;
  assign n56046 = (n30991 & n55826) | (n30991 & n56045) | (n55826 & n56045);
  assign n56047 = n30536 | n30991;
  assign n56048 = n55826 | n56047;
  assign n30994 = ~n56046 & n56048;
  assign n30995 = x143 & x203;
  assign n30996 = n30994 & n30995;
  assign n30997 = n30994 | n30995;
  assign n30998 = ~n30996 & n30997;
  assign n56049 = n30543 & n30998;
  assign n56050 = (n30998 & n55830) | (n30998 & n56049) | (n55830 & n56049);
  assign n56051 = n30543 | n30998;
  assign n56052 = n55830 | n56051;
  assign n31001 = ~n56050 & n56052;
  assign n31002 = x142 & x204;
  assign n31003 = n31001 & n31002;
  assign n31004 = n31001 | n31002;
  assign n31005 = ~n31003 & n31004;
  assign n56053 = n30550 & n31005;
  assign n56054 = (n31005 & n55834) | (n31005 & n56053) | (n55834 & n56053);
  assign n56055 = n30550 | n31005;
  assign n56056 = n55834 | n56055;
  assign n31008 = ~n56054 & n56056;
  assign n31009 = x141 & x205;
  assign n31010 = n31008 & n31009;
  assign n31011 = n31008 | n31009;
  assign n31012 = ~n31010 & n31011;
  assign n56057 = n30557 & n31012;
  assign n56058 = (n31012 & n55838) | (n31012 & n56057) | (n55838 & n56057);
  assign n56059 = n30557 | n31012;
  assign n56060 = n55838 | n56059;
  assign n31015 = ~n56058 & n56060;
  assign n31016 = x140 & x206;
  assign n31017 = n31015 & n31016;
  assign n31018 = n31015 | n31016;
  assign n31019 = ~n31017 & n31018;
  assign n56061 = n30564 & n31019;
  assign n56062 = (n31019 & n55842) | (n31019 & n56061) | (n55842 & n56061);
  assign n56063 = n30564 | n31019;
  assign n56064 = n55842 | n56063;
  assign n31022 = ~n56062 & n56064;
  assign n31023 = x139 & x207;
  assign n31024 = n31022 & n31023;
  assign n31025 = n31022 | n31023;
  assign n31026 = ~n31024 & n31025;
  assign n56065 = n30571 & n31026;
  assign n56066 = (n31026 & n55846) | (n31026 & n56065) | (n55846 & n56065);
  assign n56067 = n30571 | n31026;
  assign n56068 = n55846 | n56067;
  assign n31029 = ~n56066 & n56068;
  assign n31030 = x138 & x208;
  assign n31031 = n31029 & n31030;
  assign n31032 = n31029 | n31030;
  assign n31033 = ~n31031 & n31032;
  assign n56069 = n30578 & n31033;
  assign n56070 = (n31033 & n55850) | (n31033 & n56069) | (n55850 & n56069);
  assign n56071 = n30578 | n31033;
  assign n56072 = n55850 | n56071;
  assign n31036 = ~n56070 & n56072;
  assign n31037 = x137 & x209;
  assign n31038 = n31036 & n31037;
  assign n31039 = n31036 | n31037;
  assign n31040 = ~n31038 & n31039;
  assign n56073 = n30585 & n31040;
  assign n56074 = (n31040 & n55854) | (n31040 & n56073) | (n55854 & n56073);
  assign n56075 = n30585 | n31040;
  assign n56076 = n55854 | n56075;
  assign n31043 = ~n56074 & n56076;
  assign n31044 = x136 & x210;
  assign n31045 = n31043 & n31044;
  assign n31046 = n31043 | n31044;
  assign n31047 = ~n31045 & n31046;
  assign n56077 = n30592 & n31047;
  assign n56078 = (n31047 & n55858) | (n31047 & n56077) | (n55858 & n56077);
  assign n56079 = n30592 | n31047;
  assign n56080 = n55858 | n56079;
  assign n31050 = ~n56078 & n56080;
  assign n31051 = x135 & x211;
  assign n31052 = n31050 & n31051;
  assign n31053 = n31050 | n31051;
  assign n31054 = ~n31052 & n31053;
  assign n56081 = n30599 & n31054;
  assign n56082 = (n31054 & n55862) | (n31054 & n56081) | (n55862 & n56081);
  assign n56083 = n30599 | n31054;
  assign n56084 = n55862 | n56083;
  assign n31057 = ~n56082 & n56084;
  assign n31058 = x134 & x212;
  assign n31059 = n31057 & n31058;
  assign n31060 = n31057 | n31058;
  assign n31061 = ~n31059 & n31060;
  assign n56085 = n30606 & n31061;
  assign n56086 = (n31061 & n55866) | (n31061 & n56085) | (n55866 & n56085);
  assign n56087 = n30606 | n31061;
  assign n56088 = n55866 | n56087;
  assign n31064 = ~n56086 & n56088;
  assign n31065 = x133 & x213;
  assign n31066 = n31064 & n31065;
  assign n31067 = n31064 | n31065;
  assign n31068 = ~n31066 & n31067;
  assign n56089 = n30613 & n31068;
  assign n56090 = (n31068 & n55870) | (n31068 & n56089) | (n55870 & n56089);
  assign n56091 = n30613 | n31068;
  assign n56092 = n55870 | n56091;
  assign n31071 = ~n56090 & n56092;
  assign n31072 = x132 & x214;
  assign n31073 = n31071 & n31072;
  assign n31074 = n31071 | n31072;
  assign n31075 = ~n31073 & n31074;
  assign n56093 = n30620 & n31075;
  assign n56094 = (n31075 & n55874) | (n31075 & n56093) | (n55874 & n56093);
  assign n56095 = n30620 | n31075;
  assign n56096 = n55874 | n56095;
  assign n31078 = ~n56094 & n56096;
  assign n31079 = x131 & x215;
  assign n31080 = n31078 & n31079;
  assign n31081 = n31078 | n31079;
  assign n31082 = ~n31080 & n31081;
  assign n56097 = n30627 & n31082;
  assign n56098 = (n31082 & n55878) | (n31082 & n56097) | (n55878 & n56097);
  assign n56099 = n30627 | n31082;
  assign n56100 = n55878 | n56099;
  assign n31085 = ~n56098 & n56100;
  assign n31086 = x130 & x216;
  assign n31087 = n31085 & n31086;
  assign n31088 = n31085 | n31086;
  assign n31089 = ~n31087 & n31088;
  assign n56101 = n30634 & n31089;
  assign n56102 = (n31089 & n55883) | (n31089 & n56101) | (n55883 & n56101);
  assign n56103 = n30634 | n31089;
  assign n56104 = n55883 | n56103;
  assign n31092 = ~n56102 & n56104;
  assign n31093 = x129 & x217;
  assign n31094 = n31092 & n31093;
  assign n31095 = n31092 | n31093;
  assign n31096 = ~n31094 & n31095;
  assign n55907 = n30641 | n30643;
  assign n56105 = n31096 & n55907;
  assign n56106 = n30641 & n31096;
  assign n56107 = (n55676 & n56105) | (n55676 & n56106) | (n56105 & n56106);
  assign n56108 = n31096 | n55907;
  assign n56109 = n30641 | n31096;
  assign n56110 = (n55676 & n56108) | (n55676 & n56109) | (n56108 & n56109);
  assign n31099 = ~n56107 & n56110;
  assign n31100 = x128 & x218;
  assign n31101 = n31099 & n31100;
  assign n31102 = n31099 | n31100;
  assign n31103 = ~n31101 & n31102;
  assign n55905 = n30648 | n30650;
  assign n70197 = n31103 & n55905;
  assign n70198 = n30648 & n31103;
  assign n70199 = (n55674 & n70197) | (n55674 & n70198) | (n70197 & n70198);
  assign n70200 = n31103 | n55905;
  assign n70201 = n30648 | n31103;
  assign n70202 = (n55674 & n70200) | (n55674 & n70201) | (n70200 & n70201);
  assign n31106 = ~n70199 & n70202;
  assign n31107 = x127 & x219;
  assign n31108 = n31106 & n31107;
  assign n31109 = n31106 | n31107;
  assign n31110 = ~n31108 & n31109;
  assign n55903 = n30655 | n30657;
  assign n70203 = n31110 & n55903;
  assign n70204 = n30655 & n31110;
  assign n70205 = (n55672 & n70203) | (n55672 & n70204) | (n70203 & n70204);
  assign n70206 = n31110 | n55903;
  assign n70207 = n30655 | n31110;
  assign n70208 = (n55672 & n70206) | (n55672 & n70207) | (n70206 & n70207);
  assign n31113 = ~n70205 & n70208;
  assign n31114 = x126 & x220;
  assign n31115 = n31113 & n31114;
  assign n31116 = n31113 | n31114;
  assign n31117 = ~n31115 & n31116;
  assign n31118 = n55902 & n31117;
  assign n31119 = n55902 | n31117;
  assign n31120 = ~n31118 & n31119;
  assign n31121 = x125 & x221;
  assign n31122 = n31120 & n31121;
  assign n31123 = n31120 | n31121;
  assign n31124 = ~n31122 & n31123;
  assign n31125 = n55900 & n31124;
  assign n31126 = n55900 | n31124;
  assign n31127 = ~n31125 & n31126;
  assign n31128 = x124 & x222;
  assign n31129 = n31127 & n31128;
  assign n31130 = n31127 | n31128;
  assign n31131 = ~n31129 & n31130;
  assign n31132 = n55898 & n31131;
  assign n31133 = n55898 | n31131;
  assign n31134 = ~n31132 & n31133;
  assign n31135 = x123 & x223;
  assign n31136 = n31134 & n31135;
  assign n31137 = n31134 | n31135;
  assign n31138 = ~n31136 & n31137;
  assign n31139 = n30765 & n31138;
  assign n31140 = n30765 | n31138;
  assign n31141 = ~n31139 & n31140;
  assign n31142 = x122 & x224;
  assign n31143 = n31141 & n31142;
  assign n31144 = n31141 | n31142;
  assign n31145 = ~n31143 & n31144;
  assign n31146 = n30764 & n31145;
  assign n31147 = n30764 | n31145;
  assign n31148 = ~n31146 & n31147;
  assign n31149 = x121 & x225;
  assign n31150 = n31148 & n31149;
  assign n31151 = n31148 | n31149;
  assign n31152 = ~n31150 & n31151;
  assign n31153 = n30763 & n31152;
  assign n31154 = n30763 | n31152;
  assign n31155 = ~n31153 & n31154;
  assign n31156 = x120 & x226;
  assign n31157 = n31155 & n31156;
  assign n31158 = n31155 | n31156;
  assign n31159 = ~n31157 & n31158;
  assign n31160 = n30762 & n31159;
  assign n31161 = n30762 | n31159;
  assign n31162 = ~n31160 & n31161;
  assign n31163 = x119 & x227;
  assign n31164 = n31162 & n31163;
  assign n31165 = n31162 | n31163;
  assign n31166 = ~n31164 & n31165;
  assign n31167 = n70096 & n31166;
  assign n31168 = n70096 | n31166;
  assign n31169 = ~n31167 & n31168;
  assign n31170 = x118 & x228;
  assign n31171 = n31169 & n31170;
  assign n31172 = n31169 | n31170;
  assign n31173 = ~n31171 & n31172;
  assign n31174 = n55896 & n31173;
  assign n31175 = n55896 | n31173;
  assign n31176 = ~n31174 & n31175;
  assign n31177 = x117 & x229;
  assign n31178 = n31176 & n31177;
  assign n31179 = n31176 | n31177;
  assign n31180 = ~n31178 & n31179;
  assign n31181 = n55894 & n31180;
  assign n31182 = n55894 | n31180;
  assign n31183 = ~n31181 & n31182;
  assign n31184 = x116 & x230;
  assign n31185 = n31183 & n31184;
  assign n31186 = n31183 | n31184;
  assign n31187 = ~n31185 & n31186;
  assign n31188 = n55892 & n31187;
  assign n31189 = n55892 | n31187;
  assign n31190 = ~n31188 & n31189;
  assign n31191 = x115 & x231;
  assign n31192 = n31190 & n31191;
  assign n31193 = n31190 | n31191;
  assign n31194 = ~n31192 & n31193;
  assign n31195 = n55890 & n31194;
  assign n31196 = n55890 | n31194;
  assign n31197 = ~n31195 & n31196;
  assign n31198 = x114 & x232;
  assign n31199 = n31197 & n31198;
  assign n31200 = n31197 | n31198;
  assign n31201 = ~n31199 & n31200;
  assign n31202 = n55888 & n31201;
  assign n31203 = n55888 | n31201;
  assign n31204 = ~n31202 & n31203;
  assign n31205 = x113 & x233;
  assign n31206 = n31204 & n31205;
  assign n31207 = n31204 | n31205;
  assign n31208 = ~n31206 & n31207;
  assign n31209 = n30753 & n31208;
  assign n31210 = n30753 | n31208;
  assign n31211 = ~n31209 & n31210;
  assign n31212 = x112 & x234;
  assign n31213 = n31211 & n31212;
  assign n31214 = n31211 | n31212;
  assign n31215 = ~n31213 & n31214;
  assign n70209 = n30753 | n31205;
  assign n70210 = (n30753 & n31204) | (n30753 & n70209) | (n31204 & n70209);
  assign n56112 = (n31206 & n31208) | (n31206 & n70210) | (n31208 & n70210);
  assign n56113 = n31199 | n55888;
  assign n56114 = (n31199 & n31201) | (n31199 & n56113) | (n31201 & n56113);
  assign n56115 = n31192 | n55890;
  assign n56116 = (n31192 & n31194) | (n31192 & n56115) | (n31194 & n56115);
  assign n56117 = n31185 | n55892;
  assign n56118 = (n31185 & n31187) | (n31185 & n56117) | (n31187 & n56117);
  assign n56119 = n31178 | n55894;
  assign n56120 = (n31178 & n31180) | (n31178 & n56119) | (n31180 & n56119);
  assign n56121 = n31171 | n55896;
  assign n56122 = (n31171 & n31173) | (n31171 & n56121) | (n31173 & n56121);
  assign n70211 = n31164 | n70096;
  assign n70212 = (n31164 & n31166) | (n31164 & n70211) | (n31166 & n70211);
  assign n31223 = n31157 | n31160;
  assign n31224 = n31150 | n31153;
  assign n31225 = n31143 | n31146;
  assign n56123 = n31136 | n31138;
  assign n56124 = (n30765 & n31136) | (n30765 & n56123) | (n31136 & n56123);
  assign n56125 = n31129 | n31131;
  assign n56126 = (n31129 & n55898) | (n31129 & n56125) | (n55898 & n56125);
  assign n56127 = n31122 | n31124;
  assign n56128 = (n31122 & n55900) | (n31122 & n56127) | (n55900 & n56127);
  assign n55904 = (n30655 & n55672) | (n30655 & n55903) | (n55672 & n55903);
  assign n55906 = (n30648 & n55674) | (n30648 & n55905) | (n55674 & n55905);
  assign n55911 = (n69954 & n70098) | (n69954 & n55910) | (n70098 & n55910);
  assign n56138 = n30968 | n30970;
  assign n70213 = n30515 | n30968;
  assign n70214 = (n30968 & n30970) | (n30968 & n70213) | (n30970 & n70213);
  assign n70215 = (n55812 & n56138) | (n55812 & n70214) | (n56138 & n70214);
  assign n70216 = (n55811 & n56138) | (n55811 & n70214) | (n56138 & n70214);
  assign n70217 = (n55465 & n70215) | (n55465 & n70216) | (n70215 & n70216);
  assign n56143 = n30947 | n30949;
  assign n70218 = n30494 | n30947;
  assign n70219 = (n30947 & n30949) | (n30947 & n70218) | (n30949 & n70218);
  assign n70220 = (n55802 & n56143) | (n55802 & n70219) | (n56143 & n70219);
  assign n70221 = (n55801 & n56143) | (n55801 & n70219) | (n56143 & n70219);
  assign n70222 = (n69860 & n70220) | (n69860 & n70221) | (n70220 & n70221);
  assign n70229 = n30863 | n30865;
  assign n70230 = (n30863 & n55940) | (n30863 & n70229) | (n55940 & n70229);
  assign n70231 = n30410 | n30863;
  assign n70232 = (n30863 & n30865) | (n30863 & n70231) | (n30865 & n70231);
  assign n70233 = (n55707 & n70230) | (n55707 & n70232) | (n70230 & n70232);
  assign n70234 = (n69996 & n70230) | (n69996 & n70232) | (n70230 & n70232);
  assign n70235 = (n69730 & n70233) | (n69730 & n70234) | (n70233 & n70234);
  assign n31273 = x171 & x176;
  assign n31274 = x170 & x177;
  assign n31275 = n31273 & n31274;
  assign n31276 = n31273 | n31274;
  assign n31277 = ~n31275 & n31276;
  assign n70239 = n30814 & n31277;
  assign n70240 = (n31277 & n70138) | (n31277 & n70239) | (n70138 & n70239);
  assign n70241 = n30814 | n30816;
  assign n70243 = n31277 & n70241;
  assign n70244 = (n70139 & n70239) | (n70139 & n70243) | (n70239 & n70243);
  assign n70245 = (n69747 & n70240) | (n69747 & n70244) | (n70240 & n70244);
  assign n70246 = (n69746 & n70240) | (n69746 & n70244) | (n70240 & n70244);
  assign n70247 = (n68195 & n70245) | (n68195 & n70246) | (n70245 & n70246);
  assign n70248 = n30814 | n31277;
  assign n70249 = n70138 | n70248;
  assign n70250 = n31277 | n70241;
  assign n70251 = (n70139 & n70248) | (n70139 & n70250) | (n70248 & n70250);
  assign n70252 = (n69747 & n70249) | (n69747 & n70251) | (n70249 & n70251);
  assign n70253 = (n69746 & n70249) | (n69746 & n70251) | (n70249 & n70251);
  assign n70254 = (n68195 & n70252) | (n68195 & n70253) | (n70252 & n70253);
  assign n31280 = ~n70247 & n70254;
  assign n31281 = x169 & x178;
  assign n31282 = n31280 & n31281;
  assign n31283 = n31280 | n31281;
  assign n31284 = ~n31282 & n31283;
  assign n70255 = n30821 | n30823;
  assign n70257 = n31284 & n70255;
  assign n70258 = n30821 & n31284;
  assign n70259 = (n70150 & n70257) | (n70150 & n70258) | (n70257 & n70258);
  assign n70260 = (n30821 & n70152) | (n30821 & n70255) | (n70152 & n70255);
  assign n56191 = n31284 & n70260;
  assign n56192 = (n69887 & n70259) | (n69887 & n56191) | (n70259 & n56191);
  assign n70261 = n31284 | n70255;
  assign n70262 = n30821 | n31284;
  assign n70263 = (n70150 & n70261) | (n70150 & n70262) | (n70261 & n70262);
  assign n56194 = n31284 | n70260;
  assign n56195 = (n69887 & n70263) | (n69887 & n56194) | (n70263 & n56194);
  assign n31287 = ~n56192 & n56195;
  assign n31288 = x168 & x179;
  assign n31289 = n31287 & n31288;
  assign n31290 = n31287 | n31288;
  assign n31291 = ~n31289 & n31290;
  assign n70264 = n30375 | n30828;
  assign n70265 = (n30828 & n30830) | (n30828 & n70264) | (n30830 & n70264);
  assign n56196 = n31291 & n70265;
  assign n56176 = n30828 | n30830;
  assign n56197 = n31291 & n56176;
  assign n56198 = (n70013 & n56196) | (n70013 & n56197) | (n56196 & n56197);
  assign n56199 = n31291 | n70265;
  assign n56200 = n31291 | n56176;
  assign n56201 = (n70013 & n56199) | (n70013 & n56200) | (n56199 & n56200);
  assign n31294 = ~n56198 & n56201;
  assign n31295 = x167 & x180;
  assign n31296 = n31294 & n31295;
  assign n31297 = n31294 | n31295;
  assign n31298 = ~n31296 & n31297;
  assign n56173 = n30835 | n30837;
  assign n56202 = n31298 & n56173;
  assign n56203 = n30835 & n31298;
  assign n56204 = (n70133 & n56202) | (n70133 & n56203) | (n56202 & n56203);
  assign n56205 = n31298 | n56173;
  assign n56206 = n30835 | n31298;
  assign n56207 = (n70133 & n56205) | (n70133 & n56206) | (n56205 & n56206);
  assign n31301 = ~n56204 & n56207;
  assign n31302 = x166 & x181;
  assign n31303 = n31301 & n31302;
  assign n31304 = n31301 | n31302;
  assign n31305 = ~n31303 & n31304;
  assign n70266 = n30389 | n30842;
  assign n70267 = (n30842 & n30844) | (n30842 & n70266) | (n30844 & n70266);
  assign n56208 = n31305 & n70267;
  assign n56171 = n30842 | n30844;
  assign n56209 = n31305 & n56171;
  assign n70268 = (n55749 & n56208) | (n55749 & n56209) | (n56208 & n56209);
  assign n70269 = (n55750 & n56208) | (n55750 & n56209) | (n56208 & n56209);
  assign n70270 = (n69736 & n70268) | (n69736 & n70269) | (n70268 & n70269);
  assign n56211 = n31305 | n70267;
  assign n56212 = n31305 | n56171;
  assign n70271 = (n55749 & n56211) | (n55749 & n56212) | (n56211 & n56212);
  assign n70272 = (n55750 & n56211) | (n55750 & n56212) | (n56211 & n56212);
  assign n70273 = (n69736 & n70271) | (n69736 & n70272) | (n70271 & n70272);
  assign n31308 = ~n70270 & n70273;
  assign n31309 = x165 & x182;
  assign n31310 = n31308 & n31309;
  assign n31311 = n31308 | n31309;
  assign n31312 = ~n31310 & n31311;
  assign n70236 = n30849 | n30851;
  assign n70238 = (n30849 & n55946) | (n30849 & n70236) | (n55946 & n70236);
  assign n70274 = n31312 & n70238;
  assign n70237 = (n30849 & n70160) | (n30849 & n70236) | (n70160 & n70236);
  assign n70275 = n31312 & n70237;
  assign n70276 = (n69916 & n70274) | (n69916 & n70275) | (n70274 & n70275);
  assign n70277 = n31312 | n70238;
  assign n70278 = n31312 | n70237;
  assign n70279 = (n69916 & n70277) | (n69916 & n70278) | (n70277 & n70278);
  assign n31315 = ~n70276 & n70279;
  assign n31316 = x164 & x183;
  assign n31317 = n31315 & n31316;
  assign n31318 = n31315 | n31316;
  assign n31319 = ~n31317 & n31318;
  assign n56214 = n30856 & n31319;
  assign n70280 = (n31319 & n55984) | (n31319 & n56214) | (n55984 & n56214);
  assign n70281 = (n31319 & n56214) | (n31319 & n70162) | (n56214 & n70162);
  assign n70282 = (n69884 & n70280) | (n69884 & n70281) | (n70280 & n70281);
  assign n56216 = n30856 | n31319;
  assign n70283 = n55984 | n56216;
  assign n70284 = n56216 | n70162;
  assign n70285 = (n69884 & n70283) | (n69884 & n70284) | (n70283 & n70284);
  assign n31322 = ~n70282 & n70285;
  assign n31323 = x163 & x184;
  assign n31324 = n31322 & n31323;
  assign n31325 = n31322 | n31323;
  assign n31326 = ~n31324 & n31325;
  assign n31327 = n70235 & n31326;
  assign n31328 = n70235 | n31326;
  assign n31329 = ~n31327 & n31328;
  assign n31330 = x162 & x185;
  assign n31331 = n31329 & n31330;
  assign n31332 = n31329 | n31330;
  assign n31333 = ~n31331 & n31332;
  assign n56162 = n30870 | n30872;
  assign n56218 = n31333 & n56162;
  assign n56219 = n30870 & n31333;
  assign n56220 = (n70127 & n56218) | (n70127 & n56219) | (n56218 & n56219);
  assign n56221 = n31333 | n56162;
  assign n56222 = n30870 | n31333;
  assign n56223 = (n70127 & n56221) | (n70127 & n56222) | (n56221 & n56222);
  assign n31336 = ~n56220 & n56223;
  assign n31337 = x161 & x186;
  assign n31338 = n31336 & n31337;
  assign n31339 = n31336 | n31337;
  assign n31340 = ~n31338 & n31339;
  assign n56160 = n30877 | n55995;
  assign n70286 = n31340 & n56160;
  assign n70227 = n30424 | n30877;
  assign n70228 = (n30877 & n30879) | (n30877 & n70227) | (n30879 & n70227);
  assign n70287 = n31340 & n70228;
  assign n70288 = (n69994 & n70286) | (n69994 & n70287) | (n70286 & n70287);
  assign n70289 = n31340 | n56160;
  assign n70290 = n31340 | n70228;
  assign n70291 = (n69994 & n70289) | (n69994 & n70290) | (n70289 & n70290);
  assign n31343 = ~n70288 & n70291;
  assign n31344 = x160 & x187;
  assign n31345 = n31343 & n31344;
  assign n31346 = n31343 | n31344;
  assign n31347 = ~n31345 & n31346;
  assign n56157 = n30884 | n30886;
  assign n56224 = n31347 & n56157;
  assign n56225 = n30884 & n31347;
  assign n56226 = (n55934 & n56224) | (n55934 & n56225) | (n56224 & n56225);
  assign n56227 = n31347 | n56157;
  assign n56228 = n30884 | n31347;
  assign n56229 = (n55934 & n56227) | (n55934 & n56228) | (n56227 & n56228);
  assign n31350 = ~n56226 & n56229;
  assign n31351 = x159 & x188;
  assign n31352 = n31350 & n31351;
  assign n31353 = n31350 | n31351;
  assign n31354 = ~n31352 & n31353;
  assign n56155 = n30891 | n30893;
  assign n56230 = n31354 & n56155;
  assign n56231 = n30891 & n31354;
  assign n56232 = (n70118 & n56230) | (n70118 & n56231) | (n56230 & n56231);
  assign n56233 = n31354 | n56155;
  assign n56234 = n30891 | n31354;
  assign n56235 = (n70118 & n56233) | (n70118 & n56234) | (n56233 & n56234);
  assign n31357 = ~n56232 & n56235;
  assign n31358 = x158 & x189;
  assign n31359 = n31357 & n31358;
  assign n31360 = n31357 | n31358;
  assign n31361 = ~n31359 & n31360;
  assign n56236 = n30898 & n31361;
  assign n70292 = (n31361 & n56002) | (n31361 & n56236) | (n56002 & n56236);
  assign n70293 = (n31361 & n56001) | (n31361 & n56236) | (n56001 & n56236);
  assign n70294 = (n55698 & n70292) | (n55698 & n70293) | (n70292 & n70293);
  assign n56238 = n30898 | n31361;
  assign n70295 = n56002 | n56238;
  assign n70296 = n56001 | n56238;
  assign n70297 = (n55698 & n70295) | (n55698 & n70296) | (n70295 & n70296);
  assign n31364 = ~n70294 & n70297;
  assign n31365 = x157 & x190;
  assign n31366 = n31364 & n31365;
  assign n31367 = n31364 | n31365;
  assign n31368 = ~n31366 & n31367;
  assign n56153 = n30905 | n30907;
  assign n70298 = n31368 & n56153;
  assign n70225 = n30452 | n30905;
  assign n70226 = (n30905 & n30907) | (n30905 & n70225) | (n30907 & n70225);
  assign n70299 = n31368 & n70226;
  assign n70300 = (n55783 & n70298) | (n55783 & n70299) | (n70298 & n70299);
  assign n70301 = n31368 | n56153;
  assign n70302 = n31368 | n70226;
  assign n70303 = (n55783 & n70301) | (n55783 & n70302) | (n70301 & n70302);
  assign n31371 = ~n70300 & n70303;
  assign n31372 = x156 & x191;
  assign n31373 = n31371 & n31372;
  assign n31374 = n31371 | n31372;
  assign n31375 = ~n31373 & n31374;
  assign n56150 = n30912 | n30914;
  assign n56240 = n31375 & n56150;
  assign n56241 = n30912 & n31375;
  assign n56242 = (n70113 & n56240) | (n70113 & n56241) | (n56240 & n56241);
  assign n56243 = n31375 | n56150;
  assign n56244 = n30912 | n31375;
  assign n56245 = (n70113 & n56243) | (n70113 & n56244) | (n56243 & n56244);
  assign n31378 = ~n56242 & n56245;
  assign n31379 = x155 & x192;
  assign n31380 = n31378 & n31379;
  assign n31381 = n31378 | n31379;
  assign n31382 = ~n31380 & n31381;
  assign n56246 = n30919 & n31382;
  assign n70304 = (n31382 & n56012) | (n31382 & n56246) | (n56012 & n56246);
  assign n70305 = (n31382 & n56011) | (n31382 & n56246) | (n56011 & n56246);
  assign n70306 = (n55693 & n70304) | (n55693 & n70305) | (n70304 & n70305);
  assign n56248 = n30919 | n31382;
  assign n70307 = n56012 | n56248;
  assign n70308 = n56011 | n56248;
  assign n70309 = (n55693 & n70307) | (n55693 & n70308) | (n70307 & n70308);
  assign n31385 = ~n70306 & n70309;
  assign n31386 = x154 & x193;
  assign n31387 = n31385 & n31386;
  assign n31388 = n31385 | n31386;
  assign n31389 = ~n31387 & n31388;
  assign n56148 = n30926 | n30928;
  assign n70310 = n31389 & n56148;
  assign n70223 = n30473 | n30926;
  assign n70224 = (n30926 & n30928) | (n30926 & n70223) | (n30928 & n70223);
  assign n70311 = n31389 & n70224;
  assign n70312 = (n55793 & n70310) | (n55793 & n70311) | (n70310 & n70311);
  assign n70313 = n31389 | n56148;
  assign n70314 = n31389 | n70224;
  assign n70315 = (n55793 & n70313) | (n55793 & n70314) | (n70313 & n70314);
  assign n31392 = ~n70312 & n70315;
  assign n31393 = x153 & x194;
  assign n31394 = n31392 & n31393;
  assign n31395 = n31392 | n31393;
  assign n31396 = ~n31394 & n31395;
  assign n56145 = n30933 | n30935;
  assign n56250 = n31396 & n56145;
  assign n56251 = n30933 & n31396;
  assign n56252 = (n70108 & n56250) | (n70108 & n56251) | (n56250 & n56251);
  assign n56253 = n31396 | n56145;
  assign n56254 = n30933 | n31396;
  assign n56255 = (n70108 & n56253) | (n70108 & n56254) | (n56253 & n56254);
  assign n31399 = ~n56252 & n56255;
  assign n31400 = x152 & x195;
  assign n31401 = n31399 & n31400;
  assign n31402 = n31399 | n31400;
  assign n31403 = ~n31401 & n31402;
  assign n56256 = n30940 & n31403;
  assign n70316 = (n31403 & n56022) | (n31403 & n56256) | (n56022 & n56256);
  assign n70317 = (n31403 & n56021) | (n31403 & n56256) | (n56021 & n56256);
  assign n70318 = (n69983 & n70316) | (n69983 & n70317) | (n70316 & n70317);
  assign n56258 = n30940 | n31403;
  assign n70319 = n56022 | n56258;
  assign n70320 = n56021 | n56258;
  assign n70321 = (n69983 & n70319) | (n69983 & n70320) | (n70319 & n70320);
  assign n31406 = ~n70318 & n70321;
  assign n31407 = x151 & x196;
  assign n31408 = n31406 & n31407;
  assign n31409 = n31406 | n31407;
  assign n31410 = ~n31408 & n31409;
  assign n31411 = n70222 & n31410;
  assign n31412 = n70222 | n31410;
  assign n31413 = ~n31411 & n31412;
  assign n31414 = x150 & x197;
  assign n31415 = n31413 & n31414;
  assign n31416 = n31413 | n31414;
  assign n31417 = ~n31415 & n31416;
  assign n56140 = n30954 | n30956;
  assign n56260 = n31417 & n56140;
  assign n56261 = n30954 & n31417;
  assign n56262 = (n70103 & n56260) | (n70103 & n56261) | (n56260 & n56261);
  assign n56263 = n31417 | n56140;
  assign n56264 = n30954 | n31417;
  assign n56265 = (n70103 & n56263) | (n70103 & n56264) | (n56263 & n56264);
  assign n31420 = ~n56262 & n56265;
  assign n31421 = x149 & x198;
  assign n31422 = n31420 & n31421;
  assign n31423 = n31420 | n31421;
  assign n31424 = ~n31422 & n31423;
  assign n56266 = n30961 & n31424;
  assign n70322 = (n31424 & n56032) | (n31424 & n56266) | (n56032 & n56266);
  assign n70323 = (n31424 & n56031) | (n31424 & n56266) | (n56031 & n56266);
  assign n70324 = (n69978 & n70322) | (n69978 & n70323) | (n70322 & n70323);
  assign n56268 = n30961 | n31424;
  assign n70325 = n56032 | n56268;
  assign n70326 = n56031 | n56268;
  assign n70327 = (n69978 & n70325) | (n69978 & n70326) | (n70325 & n70326);
  assign n31427 = ~n70324 & n70327;
  assign n31428 = x148 & x199;
  assign n31429 = n31427 & n31428;
  assign n31430 = n31427 | n31428;
  assign n31431 = ~n31429 & n31430;
  assign n31432 = n70217 & n31431;
  assign n31433 = n70217 | n31431;
  assign n31434 = ~n31432 & n31433;
  assign n31435 = x147 & x200;
  assign n31436 = n31434 & n31435;
  assign n31437 = n31434 | n31435;
  assign n31438 = ~n31436 & n31437;
  assign n56135 = n30975 | n30977;
  assign n56270 = n31438 & n56135;
  assign n56271 = n30975 & n31438;
  assign n56272 = (n55911 & n56270) | (n55911 & n56271) | (n56270 & n56271);
  assign n56273 = n31438 | n56135;
  assign n56274 = n30975 | n31438;
  assign n56275 = (n55911 & n56273) | (n55911 & n56274) | (n56273 & n56274);
  assign n31441 = ~n56272 & n56275;
  assign n31442 = x146 & x201;
  assign n31443 = n31441 & n31442;
  assign n31444 = n31441 | n31442;
  assign n31445 = ~n31443 & n31444;
  assign n56276 = n30982 & n31445;
  assign n56277 = (n31445 & n70193) | (n31445 & n56276) | (n70193 & n56276);
  assign n56278 = n30982 | n31445;
  assign n56279 = n70193 | n56278;
  assign n31448 = ~n56277 & n56279;
  assign n31449 = x145 & x202;
  assign n31450 = n31448 & n31449;
  assign n31451 = n31448 | n31449;
  assign n31452 = ~n31450 & n31451;
  assign n56280 = n30989 & n31452;
  assign n56281 = (n31452 & n56046) | (n31452 & n56280) | (n56046 & n56280);
  assign n56282 = n30989 | n31452;
  assign n56283 = n56046 | n56282;
  assign n31455 = ~n56281 & n56283;
  assign n31456 = x144 & x203;
  assign n31457 = n31455 & n31456;
  assign n31458 = n31455 | n31456;
  assign n31459 = ~n31457 & n31458;
  assign n56284 = n30996 & n31459;
  assign n56285 = (n31459 & n56050) | (n31459 & n56284) | (n56050 & n56284);
  assign n56286 = n30996 | n31459;
  assign n56287 = n56050 | n56286;
  assign n31462 = ~n56285 & n56287;
  assign n31463 = x143 & x204;
  assign n31464 = n31462 & n31463;
  assign n31465 = n31462 | n31463;
  assign n31466 = ~n31464 & n31465;
  assign n56288 = n31003 & n31466;
  assign n56289 = (n31466 & n56054) | (n31466 & n56288) | (n56054 & n56288);
  assign n56290 = n31003 | n31466;
  assign n56291 = n56054 | n56290;
  assign n31469 = ~n56289 & n56291;
  assign n31470 = x142 & x205;
  assign n31471 = n31469 & n31470;
  assign n31472 = n31469 | n31470;
  assign n31473 = ~n31471 & n31472;
  assign n56292 = n31010 & n31473;
  assign n56293 = (n31473 & n56058) | (n31473 & n56292) | (n56058 & n56292);
  assign n56294 = n31010 | n31473;
  assign n56295 = n56058 | n56294;
  assign n31476 = ~n56293 & n56295;
  assign n31477 = x141 & x206;
  assign n31478 = n31476 & n31477;
  assign n31479 = n31476 | n31477;
  assign n31480 = ~n31478 & n31479;
  assign n56296 = n31017 & n31480;
  assign n56297 = (n31480 & n56062) | (n31480 & n56296) | (n56062 & n56296);
  assign n56298 = n31017 | n31480;
  assign n56299 = n56062 | n56298;
  assign n31483 = ~n56297 & n56299;
  assign n31484 = x140 & x207;
  assign n31485 = n31483 & n31484;
  assign n31486 = n31483 | n31484;
  assign n31487 = ~n31485 & n31486;
  assign n56300 = n31024 & n31487;
  assign n56301 = (n31487 & n56066) | (n31487 & n56300) | (n56066 & n56300);
  assign n56302 = n31024 | n31487;
  assign n56303 = n56066 | n56302;
  assign n31490 = ~n56301 & n56303;
  assign n31491 = x139 & x208;
  assign n31492 = n31490 & n31491;
  assign n31493 = n31490 | n31491;
  assign n31494 = ~n31492 & n31493;
  assign n56304 = n31031 & n31494;
  assign n56305 = (n31494 & n56070) | (n31494 & n56304) | (n56070 & n56304);
  assign n56306 = n31031 | n31494;
  assign n56307 = n56070 | n56306;
  assign n31497 = ~n56305 & n56307;
  assign n31498 = x138 & x209;
  assign n31499 = n31497 & n31498;
  assign n31500 = n31497 | n31498;
  assign n31501 = ~n31499 & n31500;
  assign n56308 = n31038 & n31501;
  assign n56309 = (n31501 & n56074) | (n31501 & n56308) | (n56074 & n56308);
  assign n56310 = n31038 | n31501;
  assign n56311 = n56074 | n56310;
  assign n31504 = ~n56309 & n56311;
  assign n31505 = x137 & x210;
  assign n31506 = n31504 & n31505;
  assign n31507 = n31504 | n31505;
  assign n31508 = ~n31506 & n31507;
  assign n56312 = n31045 & n31508;
  assign n56313 = (n31508 & n56078) | (n31508 & n56312) | (n56078 & n56312);
  assign n56314 = n31045 | n31508;
  assign n56315 = n56078 | n56314;
  assign n31511 = ~n56313 & n56315;
  assign n31512 = x136 & x211;
  assign n31513 = n31511 & n31512;
  assign n31514 = n31511 | n31512;
  assign n31515 = ~n31513 & n31514;
  assign n56316 = n31052 & n31515;
  assign n56317 = (n31515 & n56082) | (n31515 & n56316) | (n56082 & n56316);
  assign n56318 = n31052 | n31515;
  assign n56319 = n56082 | n56318;
  assign n31518 = ~n56317 & n56319;
  assign n31519 = x135 & x212;
  assign n31520 = n31518 & n31519;
  assign n31521 = n31518 | n31519;
  assign n31522 = ~n31520 & n31521;
  assign n56320 = n31059 & n31522;
  assign n56321 = (n31522 & n56086) | (n31522 & n56320) | (n56086 & n56320);
  assign n56322 = n31059 | n31522;
  assign n56323 = n56086 | n56322;
  assign n31525 = ~n56321 & n56323;
  assign n31526 = x134 & x213;
  assign n31527 = n31525 & n31526;
  assign n31528 = n31525 | n31526;
  assign n31529 = ~n31527 & n31528;
  assign n56324 = n31066 & n31529;
  assign n56325 = (n31529 & n56090) | (n31529 & n56324) | (n56090 & n56324);
  assign n56326 = n31066 | n31529;
  assign n56327 = n56090 | n56326;
  assign n31532 = ~n56325 & n56327;
  assign n31533 = x133 & x214;
  assign n31534 = n31532 & n31533;
  assign n31535 = n31532 | n31533;
  assign n31536 = ~n31534 & n31535;
  assign n56328 = n31073 & n31536;
  assign n56329 = (n31536 & n56094) | (n31536 & n56328) | (n56094 & n56328);
  assign n56330 = n31073 | n31536;
  assign n56331 = n56094 | n56330;
  assign n31539 = ~n56329 & n56331;
  assign n31540 = x132 & x215;
  assign n31541 = n31539 & n31540;
  assign n31542 = n31539 | n31540;
  assign n31543 = ~n31541 & n31542;
  assign n56332 = n31080 & n31543;
  assign n56333 = (n31543 & n56098) | (n31543 & n56332) | (n56098 & n56332);
  assign n56334 = n31080 | n31543;
  assign n56335 = n56098 | n56334;
  assign n31546 = ~n56333 & n56335;
  assign n31547 = x131 & x216;
  assign n31548 = n31546 & n31547;
  assign n31549 = n31546 | n31547;
  assign n31550 = ~n31548 & n31549;
  assign n56336 = n31087 & n31550;
  assign n56337 = (n31550 & n56102) | (n31550 & n56336) | (n56102 & n56336);
  assign n56338 = n31087 | n31550;
  assign n56339 = n56102 | n56338;
  assign n31553 = ~n56337 & n56339;
  assign n31554 = x130 & x217;
  assign n31555 = n31553 & n31554;
  assign n31556 = n31553 | n31554;
  assign n31557 = ~n31555 & n31556;
  assign n56340 = n31094 & n31557;
  assign n56341 = (n31557 & n56107) | (n31557 & n56340) | (n56107 & n56340);
  assign n56342 = n31094 | n31557;
  assign n56343 = n56107 | n56342;
  assign n31560 = ~n56341 & n56343;
  assign n31561 = x129 & x218;
  assign n31562 = n31560 & n31561;
  assign n31563 = n31560 | n31561;
  assign n31564 = ~n31562 & n31563;
  assign n56133 = n31101 | n31103;
  assign n56344 = n31564 & n56133;
  assign n56345 = n31101 & n31564;
  assign n56346 = (n55906 & n56344) | (n55906 & n56345) | (n56344 & n56345);
  assign n56347 = n31564 | n56133;
  assign n56348 = n31101 | n31564;
  assign n56349 = (n55906 & n56347) | (n55906 & n56348) | (n56347 & n56348);
  assign n31567 = ~n56346 & n56349;
  assign n31568 = x128 & x219;
  assign n31569 = n31567 & n31568;
  assign n31570 = n31567 | n31568;
  assign n31571 = ~n31569 & n31570;
  assign n56131 = n31108 | n31110;
  assign n70328 = n31571 & n56131;
  assign n70329 = n31108 & n31571;
  assign n70330 = (n55904 & n70328) | (n55904 & n70329) | (n70328 & n70329);
  assign n70331 = n31571 | n56131;
  assign n70332 = n31108 | n31571;
  assign n70333 = (n55904 & n70331) | (n55904 & n70332) | (n70331 & n70332);
  assign n31574 = ~n70330 & n70333;
  assign n31575 = x127 & x220;
  assign n31576 = n31574 & n31575;
  assign n31577 = n31574 | n31575;
  assign n31578 = ~n31576 & n31577;
  assign n56129 = n31115 | n31117;
  assign n70334 = n31578 & n56129;
  assign n70335 = n31115 & n31578;
  assign n70336 = (n55902 & n70334) | (n55902 & n70335) | (n70334 & n70335);
  assign n70337 = n31578 | n56129;
  assign n70338 = n31115 | n31578;
  assign n70339 = (n55902 & n70337) | (n55902 & n70338) | (n70337 & n70338);
  assign n31581 = ~n70336 & n70339;
  assign n31582 = x126 & x221;
  assign n31583 = n31581 & n31582;
  assign n31584 = n31581 | n31582;
  assign n31585 = ~n31583 & n31584;
  assign n31586 = n56128 & n31585;
  assign n31587 = n56128 | n31585;
  assign n31588 = ~n31586 & n31587;
  assign n31589 = x125 & x222;
  assign n31590 = n31588 & n31589;
  assign n31591 = n31588 | n31589;
  assign n31592 = ~n31590 & n31591;
  assign n31593 = n56126 & n31592;
  assign n31594 = n56126 | n31592;
  assign n31595 = ~n31593 & n31594;
  assign n31596 = x124 & x223;
  assign n31597 = n31595 & n31596;
  assign n31598 = n31595 | n31596;
  assign n31599 = ~n31597 & n31598;
  assign n31600 = n56124 & n31599;
  assign n31601 = n56124 | n31599;
  assign n31602 = ~n31600 & n31601;
  assign n31603 = x123 & x224;
  assign n31604 = n31602 & n31603;
  assign n31605 = n31602 | n31603;
  assign n31606 = ~n31604 & n31605;
  assign n31607 = n31225 & n31606;
  assign n31608 = n31225 | n31606;
  assign n31609 = ~n31607 & n31608;
  assign n31610 = x122 & x225;
  assign n31611 = n31609 & n31610;
  assign n31612 = n31609 | n31610;
  assign n31613 = ~n31611 & n31612;
  assign n31614 = n31224 & n31613;
  assign n31615 = n31224 | n31613;
  assign n31616 = ~n31614 & n31615;
  assign n31617 = x121 & x226;
  assign n31618 = n31616 & n31617;
  assign n31619 = n31616 | n31617;
  assign n31620 = ~n31618 & n31619;
  assign n31621 = n31223 & n31620;
  assign n31622 = n31223 | n31620;
  assign n31623 = ~n31621 & n31622;
  assign n31624 = x120 & x227;
  assign n31625 = n31623 & n31624;
  assign n31626 = n31623 | n31624;
  assign n31627 = ~n31625 & n31626;
  assign n31628 = n70212 & n31627;
  assign n31629 = n70212 | n31627;
  assign n31630 = ~n31628 & n31629;
  assign n31631 = x119 & x228;
  assign n31632 = n31630 & n31631;
  assign n31633 = n31630 | n31631;
  assign n31634 = ~n31632 & n31633;
  assign n31635 = n56122 & n31634;
  assign n31636 = n56122 | n31634;
  assign n31637 = ~n31635 & n31636;
  assign n31638 = x118 & x229;
  assign n31639 = n31637 & n31638;
  assign n31640 = n31637 | n31638;
  assign n31641 = ~n31639 & n31640;
  assign n31642 = n56120 & n31641;
  assign n31643 = n56120 | n31641;
  assign n31644 = ~n31642 & n31643;
  assign n31645 = x117 & x230;
  assign n31646 = n31644 & n31645;
  assign n31647 = n31644 | n31645;
  assign n31648 = ~n31646 & n31647;
  assign n31649 = n56118 & n31648;
  assign n31650 = n56118 | n31648;
  assign n31651 = ~n31649 & n31650;
  assign n31652 = x116 & x231;
  assign n31653 = n31651 & n31652;
  assign n31654 = n31651 | n31652;
  assign n31655 = ~n31653 & n31654;
  assign n31656 = n56116 & n31655;
  assign n31657 = n56116 | n31655;
  assign n31658 = ~n31656 & n31657;
  assign n31659 = x115 & x232;
  assign n31660 = n31658 & n31659;
  assign n31661 = n31658 | n31659;
  assign n31662 = ~n31660 & n31661;
  assign n31663 = n56114 & n31662;
  assign n31664 = n56114 | n31662;
  assign n31665 = ~n31663 & n31664;
  assign n31666 = x114 & x233;
  assign n31667 = n31665 & n31666;
  assign n31668 = n31665 | n31666;
  assign n31669 = ~n31667 & n31668;
  assign n31670 = n56112 & n31669;
  assign n31671 = n56112 | n31669;
  assign n31672 = ~n31670 & n31671;
  assign n31673 = x113 & x234;
  assign n31674 = n31672 & n31673;
  assign n31675 = n31672 | n31673;
  assign n31676 = ~n31674 & n31675;
  assign n31677 = n31213 & n31676;
  assign n31678 = n31213 | n31676;
  assign n31679 = ~n31677 & n31678;
  assign n31680 = x112 & x235;
  assign n31681 = n31679 & n31680;
  assign n31682 = n31679 | n31680;
  assign n31683 = ~n31681 & n31682;
  assign n70340 = n31213 | n31673;
  assign n70341 = (n31213 & n31672) | (n31213 & n70340) | (n31672 & n70340);
  assign n56351 = (n31674 & n31676) | (n31674 & n70341) | (n31676 & n70341);
  assign n56352 = n31667 | n56112;
  assign n56353 = (n31667 & n31669) | (n31667 & n56352) | (n31669 & n56352);
  assign n56354 = n31660 | n56114;
  assign n56355 = (n31660 & n31662) | (n31660 & n56354) | (n31662 & n56354);
  assign n56356 = n31653 | n56116;
  assign n56357 = (n31653 & n31655) | (n31653 & n56356) | (n31655 & n56356);
  assign n56358 = n31646 | n56118;
  assign n56359 = (n31646 & n31648) | (n31646 & n56358) | (n31648 & n56358);
  assign n56360 = n31639 | n56120;
  assign n56361 = (n31639 & n31641) | (n31639 & n56360) | (n31641 & n56360);
  assign n56362 = n31632 | n56122;
  assign n56363 = (n31632 & n31634) | (n31632 & n56362) | (n31634 & n56362);
  assign n70342 = n31625 | n70212;
  assign n70343 = (n31625 & n31627) | (n31625 & n70342) | (n31627 & n70342);
  assign n31692 = n31618 | n31621;
  assign n31693 = n31611 | n31614;
  assign n56364 = n31604 | n31606;
  assign n56365 = (n31225 & n31604) | (n31225 & n56364) | (n31604 & n56364);
  assign n56366 = n31597 | n31599;
  assign n56367 = (n31597 & n56124) | (n31597 & n56366) | (n56124 & n56366);
  assign n56368 = n31590 | n31592;
  assign n56369 = (n31590 & n56126) | (n31590 & n56368) | (n56126 & n56368);
  assign n56130 = (n31115 & n55902) | (n31115 & n56129) | (n55902 & n56129);
  assign n56132 = (n31108 & n55904) | (n31108 & n56131) | (n55904 & n56131);
  assign n56382 = n31422 | n31424;
  assign n70346 = n30961 | n31422;
  assign n70347 = (n31422 & n31424) | (n31422 & n70346) | (n31424 & n70346);
  assign n70348 = (n56032 & n56382) | (n56032 & n70347) | (n56382 & n70347);
  assign n70349 = (n56031 & n56382) | (n56031 & n70347) | (n56382 & n70347);
  assign n70350 = (n69978 & n70348) | (n69978 & n70349) | (n70348 & n70349);
  assign n56387 = n31401 | n31403;
  assign n70351 = n30940 | n31401;
  assign n70352 = (n31401 & n31403) | (n31401 & n70351) | (n31403 & n70351);
  assign n70353 = (n56022 & n56387) | (n56022 & n70352) | (n56387 & n70352);
  assign n70354 = (n56021 & n56387) | (n56021 & n70352) | (n56387 & n70352);
  assign n70355 = (n69983 & n70353) | (n69983 & n70354) | (n70353 & n70354);
  assign n56149 = (n55793 & n70224) | (n55793 & n56148) | (n70224 & n56148);
  assign n56392 = n31380 | n31382;
  assign n70356 = n30919 | n31380;
  assign n70357 = (n31380 & n31382) | (n31380 & n70356) | (n31382 & n70356);
  assign n70358 = (n56012 & n56392) | (n56012 & n70357) | (n56392 & n70357);
  assign n70359 = (n56011 & n56392) | (n56011 & n70357) | (n56392 & n70357);
  assign n70360 = (n55693 & n70358) | (n55693 & n70359) | (n70358 & n70359);
  assign n56154 = (n55783 & n70226) | (n55783 & n56153) | (n70226 & n56153);
  assign n56397 = n31359 | n31361;
  assign n70361 = n30898 | n31359;
  assign n70362 = (n31359 & n31361) | (n31359 & n70361) | (n31361 & n70361);
  assign n70363 = (n56002 & n56397) | (n56002 & n70362) | (n56397 & n70362);
  assign n70364 = (n56001 & n56397) | (n56001 & n70362) | (n56397 & n70362);
  assign n70365 = (n55698 & n70363) | (n55698 & n70364) | (n70363 & n70364);
  assign n31742 = x172 & x176;
  assign n31743 = x171 & x177;
  assign n31744 = n31742 & n31743;
  assign n31745 = n31742 | n31743;
  assign n31746 = ~n31744 & n31745;
  assign n70378 = n31275 | n70239;
  assign n70381 = n31746 & n70378;
  assign n70379 = n31275 | n31277;
  assign n70382 = n31746 & n70379;
  assign n70383 = (n70138 & n70381) | (n70138 & n70382) | (n70381 & n70382);
  assign n70384 = n31275 & n31746;
  assign n70385 = (n31746 & n70244) | (n31746 & n70384) | (n70244 & n70384);
  assign n70386 = (n69747 & n70383) | (n69747 & n70385) | (n70383 & n70385);
  assign n70387 = (n69746 & n70383) | (n69746 & n70385) | (n70383 & n70385);
  assign n70388 = (n68195 & n70386) | (n68195 & n70387) | (n70386 & n70387);
  assign n70389 = n31746 | n70378;
  assign n70390 = n31746 | n70379;
  assign n70391 = (n70138 & n70389) | (n70138 & n70390) | (n70389 & n70390);
  assign n70392 = n31275 | n31746;
  assign n70393 = n70244 | n70392;
  assign n70394 = (n69747 & n70391) | (n69747 & n70393) | (n70391 & n70393);
  assign n70395 = (n69746 & n70391) | (n69746 & n70393) | (n70391 & n70393);
  assign n70396 = (n68195 & n70394) | (n68195 & n70395) | (n70394 & n70395);
  assign n31749 = ~n70388 & n70396;
  assign n31750 = x170 & x178;
  assign n31751 = n31749 & n31750;
  assign n31752 = n31749 | n31750;
  assign n31753 = ~n31751 & n31752;
  assign n70397 = n31282 & n31753;
  assign n70398 = (n31753 & n70259) | (n31753 & n70397) | (n70259 & n70397);
  assign n70399 = n31282 | n31284;
  assign n70401 = n31753 & n70399;
  assign n70402 = (n70260 & n70397) | (n70260 & n70401) | (n70397 & n70401);
  assign n56437 = (n69887 & n70398) | (n69887 & n70402) | (n70398 & n70402);
  assign n70403 = n31282 | n31753;
  assign n70404 = n70259 | n70403;
  assign n70405 = n31753 | n70399;
  assign n70406 = (n70260 & n70403) | (n70260 & n70405) | (n70403 & n70405);
  assign n56440 = (n69887 & n70404) | (n69887 & n70406) | (n70404 & n70406);
  assign n31756 = ~n56437 & n56440;
  assign n31757 = x169 & x179;
  assign n31758 = n31756 & n31757;
  assign n31759 = n31756 | n31757;
  assign n31760 = ~n31758 & n31759;
  assign n70407 = n31289 | n31291;
  assign n70408 = (n31289 & n70265) | (n31289 & n70407) | (n70265 & n70407);
  assign n56441 = n31760 & n70408;
  assign n70409 = (n31289 & n56176) | (n31289 & n70407) | (n56176 & n70407);
  assign n56442 = n31760 & n70409;
  assign n56443 = (n70013 & n56441) | (n70013 & n56442) | (n56441 & n56442);
  assign n56444 = n31760 | n70408;
  assign n56445 = n31760 | n70409;
  assign n56446 = (n70013 & n56444) | (n70013 & n56445) | (n56444 & n56445);
  assign n31763 = ~n56443 & n56446;
  assign n31764 = x168 & x180;
  assign n31765 = n31763 & n31764;
  assign n31766 = n31763 | n31764;
  assign n31767 = ~n31765 & n31766;
  assign n70410 = n31296 | n31298;
  assign n70411 = (n31296 & n56173) | (n31296 & n70410) | (n56173 & n70410);
  assign n56447 = n31767 & n70411;
  assign n70412 = n30835 | n31296;
  assign n70413 = (n31296 & n31298) | (n31296 & n70412) | (n31298 & n70412);
  assign n56448 = n31767 & n70413;
  assign n56449 = (n70133 & n56447) | (n70133 & n56448) | (n56447 & n56448);
  assign n56450 = n31767 | n70411;
  assign n56451 = n31767 | n70413;
  assign n56452 = (n70133 & n56450) | (n70133 & n56451) | (n56450 & n56451);
  assign n31770 = ~n56449 & n56452;
  assign n31771 = x167 & x181;
  assign n31772 = n31770 & n31771;
  assign n31773 = n31770 | n31771;
  assign n31774 = ~n31772 & n31773;
  assign n70372 = n31303 | n31305;
  assign n70373 = (n31303 & n70267) | (n31303 & n70372) | (n70267 & n70372);
  assign n70374 = (n31303 & n56171) | (n31303 & n70372) | (n56171 & n70372);
  assign n70376 = (n55750 & n70373) | (n55750 & n70374) | (n70373 & n70374);
  assign n70414 = n31774 & n70376;
  assign n70375 = (n55749 & n70373) | (n55749 & n70374) | (n70373 & n70374);
  assign n70415 = n31774 & n70375;
  assign n70416 = (n69736 & n70414) | (n69736 & n70415) | (n70414 & n70415);
  assign n70417 = n31774 | n70376;
  assign n70418 = n31774 | n70375;
  assign n70419 = (n69736 & n70417) | (n69736 & n70418) | (n70417 & n70418);
  assign n31777 = ~n70416 & n70419;
  assign n31778 = x166 & x182;
  assign n31779 = n31777 & n31778;
  assign n31780 = n31777 | n31778;
  assign n31781 = ~n31779 & n31780;
  assign n56412 = n31310 | n31312;
  assign n56453 = n31781 & n56412;
  assign n56454 = n31310 & n31781;
  assign n70420 = (n56453 & n56454) | (n56453 & n70238) | (n56454 & n70238);
  assign n70421 = (n56453 & n56454) | (n56453 & n70237) | (n56454 & n70237);
  assign n70422 = (n69916 & n70420) | (n69916 & n70421) | (n70420 & n70421);
  assign n56456 = n31781 | n56412;
  assign n56457 = n31310 | n31781;
  assign n70423 = (n56456 & n56457) | (n56456 & n70238) | (n56457 & n70238);
  assign n70424 = (n56456 & n56457) | (n56456 & n70237) | (n56457 & n70237);
  assign n70425 = (n69916 & n70423) | (n69916 & n70424) | (n70423 & n70424);
  assign n31784 = ~n70422 & n70425;
  assign n31785 = x165 & x183;
  assign n31786 = n31784 & n31785;
  assign n31787 = n31784 | n31785;
  assign n31788 = ~n31786 & n31787;
  assign n70426 = n30856 | n31317;
  assign n70427 = (n31317 & n31319) | (n31317 & n70426) | (n31319 & n70426);
  assign n56459 = n31788 & n70427;
  assign n56410 = n31317 | n31319;
  assign n56460 = n31788 & n56410;
  assign n70428 = (n55984 & n56459) | (n55984 & n56460) | (n56459 & n56460);
  assign n70429 = (n56459 & n56460) | (n56459 & n70162) | (n56460 & n70162);
  assign n70430 = (n69884 & n70428) | (n69884 & n70429) | (n70428 & n70429);
  assign n56462 = n31788 | n70427;
  assign n56463 = n31788 | n56410;
  assign n70431 = (n55984 & n56462) | (n55984 & n56463) | (n56462 & n56463);
  assign n70432 = (n56462 & n56463) | (n56462 & n70162) | (n56463 & n70162);
  assign n70433 = (n69884 & n70431) | (n69884 & n70432) | (n70431 & n70432);
  assign n31791 = ~n70430 & n70433;
  assign n31792 = x164 & x184;
  assign n31793 = n31791 & n31792;
  assign n31794 = n31791 | n31792;
  assign n31795 = ~n31793 & n31794;
  assign n56407 = n31324 | n31326;
  assign n56465 = n31795 & n56407;
  assign n56466 = n31324 & n31795;
  assign n56467 = (n70235 & n56465) | (n70235 & n56466) | (n56465 & n56466);
  assign n56468 = n31795 | n56407;
  assign n56469 = n31324 | n31795;
  assign n56470 = (n70235 & n56468) | (n70235 & n56469) | (n56468 & n56469);
  assign n31798 = ~n56467 & n56470;
  assign n31799 = x163 & x185;
  assign n31800 = n31798 & n31799;
  assign n31801 = n31798 | n31799;
  assign n31802 = ~n31800 & n31801;
  assign n56405 = n31331 | n56218;
  assign n70434 = n31802 & n56405;
  assign n70370 = n30870 | n31331;
  assign n70371 = (n31331 & n31333) | (n31331 & n70370) | (n31333 & n70370);
  assign n70435 = n31802 & n70371;
  assign n70436 = (n70127 & n70434) | (n70127 & n70435) | (n70434 & n70435);
  assign n70437 = n31802 | n56405;
  assign n70438 = n31802 | n70371;
  assign n70439 = (n70127 & n70437) | (n70127 & n70438) | (n70437 & n70438);
  assign n31805 = ~n70436 & n70439;
  assign n31806 = x162 & x186;
  assign n31807 = n31805 & n31806;
  assign n31808 = n31805 | n31806;
  assign n31809 = ~n31807 & n31808;
  assign n56402 = n31338 | n31340;
  assign n56471 = n31809 & n56402;
  assign n56472 = n31338 & n31809;
  assign n70440 = (n56160 & n56471) | (n56160 & n56472) | (n56471 & n56472);
  assign n70441 = (n56471 & n56472) | (n56471 & n70228) | (n56472 & n70228);
  assign n70442 = (n69994 & n70440) | (n69994 & n70441) | (n70440 & n70441);
  assign n56474 = n31809 | n56402;
  assign n56475 = n31338 | n31809;
  assign n70443 = (n56160 & n56474) | (n56160 & n56475) | (n56474 & n56475);
  assign n70444 = (n56474 & n56475) | (n56474 & n70228) | (n56475 & n70228);
  assign n70445 = (n69994 & n70443) | (n69994 & n70444) | (n70443 & n70444);
  assign n31812 = ~n70442 & n70445;
  assign n31813 = x161 & x187;
  assign n31814 = n31812 & n31813;
  assign n31815 = n31812 | n31813;
  assign n31816 = ~n31814 & n31815;
  assign n70368 = n31345 | n31347;
  assign n70369 = (n31345 & n56157) | (n31345 & n70368) | (n56157 & n70368);
  assign n70446 = n31816 & n70369;
  assign n70366 = n30884 | n31345;
  assign n70367 = (n31345 & n31347) | (n31345 & n70366) | (n31347 & n70366);
  assign n70447 = n31816 & n70367;
  assign n70448 = (n55934 & n70446) | (n55934 & n70447) | (n70446 & n70447);
  assign n70449 = n31816 | n70369;
  assign n70450 = n31816 | n70367;
  assign n70451 = (n55934 & n70449) | (n55934 & n70450) | (n70449 & n70450);
  assign n31819 = ~n70448 & n70451;
  assign n31820 = x160 & x188;
  assign n31821 = n31819 & n31820;
  assign n31822 = n31819 | n31820;
  assign n31823 = ~n31821 & n31822;
  assign n56477 = n31352 & n31823;
  assign n56478 = (n31823 & n56232) | (n31823 & n56477) | (n56232 & n56477);
  assign n56479 = n31352 | n31823;
  assign n56480 = n56232 | n56479;
  assign n31826 = ~n56478 & n56480;
  assign n31827 = x159 & x189;
  assign n31828 = n31826 & n31827;
  assign n31829 = n31826 | n31827;
  assign n31830 = ~n31828 & n31829;
  assign n31831 = n70365 & n31830;
  assign n31832 = n70365 | n31830;
  assign n31833 = ~n31831 & n31832;
  assign n31834 = x158 & x190;
  assign n31835 = n31833 & n31834;
  assign n31836 = n31833 | n31834;
  assign n31837 = ~n31835 & n31836;
  assign n56394 = n31366 | n31368;
  assign n56481 = n31837 & n56394;
  assign n56482 = n31366 & n31837;
  assign n56483 = (n56154 & n56481) | (n56154 & n56482) | (n56481 & n56482);
  assign n56484 = n31837 | n56394;
  assign n56485 = n31366 | n31837;
  assign n56486 = (n56154 & n56484) | (n56154 & n56485) | (n56484 & n56485);
  assign n31840 = ~n56483 & n56486;
  assign n31841 = x157 & x191;
  assign n31842 = n31840 & n31841;
  assign n31843 = n31840 | n31841;
  assign n31844 = ~n31842 & n31843;
  assign n56487 = n31373 & n31844;
  assign n56488 = (n31844 & n56242) | (n31844 & n56487) | (n56242 & n56487);
  assign n56489 = n31373 | n31844;
  assign n56490 = n56242 | n56489;
  assign n31847 = ~n56488 & n56490;
  assign n31848 = x156 & x192;
  assign n31849 = n31847 & n31848;
  assign n31850 = n31847 | n31848;
  assign n31851 = ~n31849 & n31850;
  assign n31852 = n70360 & n31851;
  assign n31853 = n70360 | n31851;
  assign n31854 = ~n31852 & n31853;
  assign n31855 = x155 & x193;
  assign n31856 = n31854 & n31855;
  assign n31857 = n31854 | n31855;
  assign n31858 = ~n31856 & n31857;
  assign n56389 = n31387 | n31389;
  assign n56491 = n31858 & n56389;
  assign n56492 = n31387 & n31858;
  assign n56493 = (n56149 & n56491) | (n56149 & n56492) | (n56491 & n56492);
  assign n56494 = n31858 | n56389;
  assign n56495 = n31387 | n31858;
  assign n56496 = (n56149 & n56494) | (n56149 & n56495) | (n56494 & n56495);
  assign n31861 = ~n56493 & n56496;
  assign n31862 = x154 & x194;
  assign n31863 = n31861 & n31862;
  assign n31864 = n31861 | n31862;
  assign n31865 = ~n31863 & n31864;
  assign n56497 = n31394 & n31865;
  assign n56498 = (n31865 & n56252) | (n31865 & n56497) | (n56252 & n56497);
  assign n56499 = n31394 | n31865;
  assign n56500 = n56252 | n56499;
  assign n31868 = ~n56498 & n56500;
  assign n31869 = x153 & x195;
  assign n31870 = n31868 & n31869;
  assign n31871 = n31868 | n31869;
  assign n31872 = ~n31870 & n31871;
  assign n31873 = n70355 & n31872;
  assign n31874 = n70355 | n31872;
  assign n31875 = ~n31873 & n31874;
  assign n31876 = x152 & x196;
  assign n31877 = n31875 & n31876;
  assign n31878 = n31875 | n31876;
  assign n31879 = ~n31877 & n31878;
  assign n56384 = n31408 | n31410;
  assign n56501 = n31879 & n56384;
  assign n56502 = n31408 & n31879;
  assign n56503 = (n70222 & n56501) | (n70222 & n56502) | (n56501 & n56502);
  assign n56504 = n31879 | n56384;
  assign n56505 = n31408 | n31879;
  assign n56506 = (n70222 & n56504) | (n70222 & n56505) | (n56504 & n56505);
  assign n31882 = ~n56503 & n56506;
  assign n31883 = x151 & x197;
  assign n31884 = n31882 & n31883;
  assign n31885 = n31882 | n31883;
  assign n31886 = ~n31884 & n31885;
  assign n56507 = n31415 & n31886;
  assign n70452 = (n31886 & n56261) | (n31886 & n56507) | (n56261 & n56507);
  assign n70453 = (n31886 & n56260) | (n31886 & n56507) | (n56260 & n56507);
  assign n70454 = (n70103 & n70452) | (n70103 & n70453) | (n70452 & n70453);
  assign n56509 = n31415 | n31886;
  assign n70455 = n56261 | n56509;
  assign n70456 = n56260 | n56509;
  assign n70457 = (n70103 & n70455) | (n70103 & n70456) | (n70455 & n70456);
  assign n31889 = ~n70454 & n70457;
  assign n31890 = x150 & x198;
  assign n31891 = n31889 & n31890;
  assign n31892 = n31889 | n31890;
  assign n31893 = ~n31891 & n31892;
  assign n31894 = n70350 & n31893;
  assign n31895 = n70350 | n31893;
  assign n31896 = ~n31894 & n31895;
  assign n31897 = x149 & x199;
  assign n31898 = n31896 & n31897;
  assign n31899 = n31896 | n31897;
  assign n31900 = ~n31898 & n31899;
  assign n56379 = n31429 | n31431;
  assign n56511 = n31900 & n56379;
  assign n56512 = n31429 & n31900;
  assign n56513 = (n70217 & n56511) | (n70217 & n56512) | (n56511 & n56512);
  assign n56514 = n31900 | n56379;
  assign n56515 = n31429 | n31900;
  assign n56516 = (n70217 & n56514) | (n70217 & n56515) | (n56514 & n56515);
  assign n31903 = ~n56513 & n56516;
  assign n31904 = x148 & x200;
  assign n31905 = n31903 & n31904;
  assign n31906 = n31903 | n31904;
  assign n31907 = ~n31905 & n31906;
  assign n56517 = n31436 & n31907;
  assign n70458 = (n31907 & n56271) | (n31907 & n56517) | (n56271 & n56517);
  assign n70459 = (n31907 & n56270) | (n31907 & n56517) | (n56270 & n56517);
  assign n70460 = (n55911 & n70458) | (n55911 & n70459) | (n70458 & n70459);
  assign n56519 = n31436 | n31907;
  assign n70461 = n56271 | n56519;
  assign n70462 = n56270 | n56519;
  assign n70463 = (n55911 & n70461) | (n55911 & n70462) | (n70461 & n70462);
  assign n31910 = ~n70460 & n70463;
  assign n31911 = x147 & x201;
  assign n31912 = n31910 & n31911;
  assign n31913 = n31910 | n31911;
  assign n31914 = ~n31912 & n31913;
  assign n56377 = n31443 | n31445;
  assign n70464 = n31914 & n56377;
  assign n70344 = n30982 | n31443;
  assign n70345 = (n31443 & n31445) | (n31443 & n70344) | (n31445 & n70344);
  assign n70465 = n31914 & n70345;
  assign n70466 = (n70193 & n70464) | (n70193 & n70465) | (n70464 & n70465);
  assign n70467 = n31914 | n56377;
  assign n70468 = n31914 | n70345;
  assign n70469 = (n70193 & n70467) | (n70193 & n70468) | (n70467 & n70468);
  assign n31917 = ~n70466 & n70469;
  assign n31918 = x146 & x202;
  assign n31919 = n31917 & n31918;
  assign n31920 = n31917 | n31918;
  assign n31921 = ~n31919 & n31920;
  assign n56521 = n31450 & n31921;
  assign n70470 = (n31921 & n56280) | (n31921 & n56521) | (n56280 & n56521);
  assign n70471 = (n31452 & n31921) | (n31452 & n56521) | (n31921 & n56521);
  assign n70472 = (n56046 & n70470) | (n56046 & n70471) | (n70470 & n70471);
  assign n56523 = n31450 | n31921;
  assign n70473 = n56280 | n56523;
  assign n70474 = n31452 | n56523;
  assign n70475 = (n56046 & n70473) | (n56046 & n70474) | (n70473 & n70474);
  assign n31924 = ~n70472 & n70475;
  assign n31925 = x145 & x203;
  assign n31926 = n31924 & n31925;
  assign n31927 = n31924 | n31925;
  assign n31928 = ~n31926 & n31927;
  assign n56525 = n31457 & n31928;
  assign n56526 = (n31928 & n56285) | (n31928 & n56525) | (n56285 & n56525);
  assign n56527 = n31457 | n31928;
  assign n56528 = n56285 | n56527;
  assign n31931 = ~n56526 & n56528;
  assign n31932 = x144 & x204;
  assign n31933 = n31931 & n31932;
  assign n31934 = n31931 | n31932;
  assign n31935 = ~n31933 & n31934;
  assign n56529 = n31464 & n31935;
  assign n56530 = (n31935 & n56289) | (n31935 & n56529) | (n56289 & n56529);
  assign n56531 = n31464 | n31935;
  assign n56532 = n56289 | n56531;
  assign n31938 = ~n56530 & n56532;
  assign n31939 = x143 & x205;
  assign n31940 = n31938 & n31939;
  assign n31941 = n31938 | n31939;
  assign n31942 = ~n31940 & n31941;
  assign n56533 = n31471 & n31942;
  assign n56534 = (n31942 & n56293) | (n31942 & n56533) | (n56293 & n56533);
  assign n56535 = n31471 | n31942;
  assign n56536 = n56293 | n56535;
  assign n31945 = ~n56534 & n56536;
  assign n31946 = x142 & x206;
  assign n31947 = n31945 & n31946;
  assign n31948 = n31945 | n31946;
  assign n31949 = ~n31947 & n31948;
  assign n56537 = n31478 & n31949;
  assign n56538 = (n31949 & n56297) | (n31949 & n56537) | (n56297 & n56537);
  assign n56539 = n31478 | n31949;
  assign n56540 = n56297 | n56539;
  assign n31952 = ~n56538 & n56540;
  assign n31953 = x141 & x207;
  assign n31954 = n31952 & n31953;
  assign n31955 = n31952 | n31953;
  assign n31956 = ~n31954 & n31955;
  assign n56541 = n31485 & n31956;
  assign n56542 = (n31956 & n56301) | (n31956 & n56541) | (n56301 & n56541);
  assign n56543 = n31485 | n31956;
  assign n56544 = n56301 | n56543;
  assign n31959 = ~n56542 & n56544;
  assign n31960 = x140 & x208;
  assign n31961 = n31959 & n31960;
  assign n31962 = n31959 | n31960;
  assign n31963 = ~n31961 & n31962;
  assign n56545 = n31492 & n31963;
  assign n56546 = (n31963 & n56305) | (n31963 & n56545) | (n56305 & n56545);
  assign n56547 = n31492 | n31963;
  assign n56548 = n56305 | n56547;
  assign n31966 = ~n56546 & n56548;
  assign n31967 = x139 & x209;
  assign n31968 = n31966 & n31967;
  assign n31969 = n31966 | n31967;
  assign n31970 = ~n31968 & n31969;
  assign n56549 = n31499 & n31970;
  assign n56550 = (n31970 & n56309) | (n31970 & n56549) | (n56309 & n56549);
  assign n56551 = n31499 | n31970;
  assign n56552 = n56309 | n56551;
  assign n31973 = ~n56550 & n56552;
  assign n31974 = x138 & x210;
  assign n31975 = n31973 & n31974;
  assign n31976 = n31973 | n31974;
  assign n31977 = ~n31975 & n31976;
  assign n56553 = n31506 & n31977;
  assign n56554 = (n31977 & n56313) | (n31977 & n56553) | (n56313 & n56553);
  assign n56555 = n31506 | n31977;
  assign n56556 = n56313 | n56555;
  assign n31980 = ~n56554 & n56556;
  assign n31981 = x137 & x211;
  assign n31982 = n31980 & n31981;
  assign n31983 = n31980 | n31981;
  assign n31984 = ~n31982 & n31983;
  assign n56557 = n31513 & n31984;
  assign n56558 = (n31984 & n56317) | (n31984 & n56557) | (n56317 & n56557);
  assign n56559 = n31513 | n31984;
  assign n56560 = n56317 | n56559;
  assign n31987 = ~n56558 & n56560;
  assign n31988 = x136 & x212;
  assign n31989 = n31987 & n31988;
  assign n31990 = n31987 | n31988;
  assign n31991 = ~n31989 & n31990;
  assign n56561 = n31520 & n31991;
  assign n56562 = (n31991 & n56321) | (n31991 & n56561) | (n56321 & n56561);
  assign n56563 = n31520 | n31991;
  assign n56564 = n56321 | n56563;
  assign n31994 = ~n56562 & n56564;
  assign n31995 = x135 & x213;
  assign n31996 = n31994 & n31995;
  assign n31997 = n31994 | n31995;
  assign n31998 = ~n31996 & n31997;
  assign n56565 = n31527 & n31998;
  assign n56566 = (n31998 & n56325) | (n31998 & n56565) | (n56325 & n56565);
  assign n56567 = n31527 | n31998;
  assign n56568 = n56325 | n56567;
  assign n32001 = ~n56566 & n56568;
  assign n32002 = x134 & x214;
  assign n32003 = n32001 & n32002;
  assign n32004 = n32001 | n32002;
  assign n32005 = ~n32003 & n32004;
  assign n56569 = n31534 & n32005;
  assign n56570 = (n32005 & n56329) | (n32005 & n56569) | (n56329 & n56569);
  assign n56571 = n31534 | n32005;
  assign n56572 = n56329 | n56571;
  assign n32008 = ~n56570 & n56572;
  assign n32009 = x133 & x215;
  assign n32010 = n32008 & n32009;
  assign n32011 = n32008 | n32009;
  assign n32012 = ~n32010 & n32011;
  assign n56573 = n31541 & n32012;
  assign n56574 = (n32012 & n56333) | (n32012 & n56573) | (n56333 & n56573);
  assign n56575 = n31541 | n32012;
  assign n56576 = n56333 | n56575;
  assign n32015 = ~n56574 & n56576;
  assign n32016 = x132 & x216;
  assign n32017 = n32015 & n32016;
  assign n32018 = n32015 | n32016;
  assign n32019 = ~n32017 & n32018;
  assign n56577 = n31548 & n32019;
  assign n56578 = (n32019 & n56337) | (n32019 & n56577) | (n56337 & n56577);
  assign n56579 = n31548 | n32019;
  assign n56580 = n56337 | n56579;
  assign n32022 = ~n56578 & n56580;
  assign n32023 = x131 & x217;
  assign n32024 = n32022 & n32023;
  assign n32025 = n32022 | n32023;
  assign n32026 = ~n32024 & n32025;
  assign n56581 = n31555 & n32026;
  assign n56582 = (n32026 & n56341) | (n32026 & n56581) | (n56341 & n56581);
  assign n56583 = n31555 | n32026;
  assign n56584 = n56341 | n56583;
  assign n32029 = ~n56582 & n56584;
  assign n32030 = x130 & x218;
  assign n32031 = n32029 & n32030;
  assign n32032 = n32029 | n32030;
  assign n32033 = ~n32031 & n32032;
  assign n56585 = n31562 & n32033;
  assign n56586 = (n32033 & n56346) | (n32033 & n56585) | (n56346 & n56585);
  assign n56587 = n31562 | n32033;
  assign n56588 = n56346 | n56587;
  assign n32036 = ~n56586 & n56588;
  assign n32037 = x129 & x219;
  assign n32038 = n32036 & n32037;
  assign n32039 = n32036 | n32037;
  assign n32040 = ~n32038 & n32039;
  assign n56374 = n31569 | n31571;
  assign n56589 = n32040 & n56374;
  assign n56590 = n31569 & n32040;
  assign n56591 = (n56132 & n56589) | (n56132 & n56590) | (n56589 & n56590);
  assign n56592 = n32040 | n56374;
  assign n56593 = n31569 | n32040;
  assign n56594 = (n56132 & n56592) | (n56132 & n56593) | (n56592 & n56593);
  assign n32043 = ~n56591 & n56594;
  assign n32044 = x128 & x220;
  assign n32045 = n32043 & n32044;
  assign n32046 = n32043 | n32044;
  assign n32047 = ~n32045 & n32046;
  assign n56372 = n31576 | n31578;
  assign n70476 = n32047 & n56372;
  assign n70477 = n31576 & n32047;
  assign n70478 = (n56130 & n70476) | (n56130 & n70477) | (n70476 & n70477);
  assign n70479 = n32047 | n56372;
  assign n70480 = n31576 | n32047;
  assign n70481 = (n56130 & n70479) | (n56130 & n70480) | (n70479 & n70480);
  assign n32050 = ~n70478 & n70481;
  assign n32051 = x127 & x221;
  assign n32052 = n32050 & n32051;
  assign n32053 = n32050 | n32051;
  assign n32054 = ~n32052 & n32053;
  assign n56370 = n31583 | n31585;
  assign n70482 = n32054 & n56370;
  assign n70483 = n31583 & n32054;
  assign n70484 = (n56128 & n70482) | (n56128 & n70483) | (n70482 & n70483);
  assign n70485 = n32054 | n56370;
  assign n70486 = n31583 | n32054;
  assign n70487 = (n56128 & n70485) | (n56128 & n70486) | (n70485 & n70486);
  assign n32057 = ~n70484 & n70487;
  assign n32058 = x126 & x222;
  assign n32059 = n32057 & n32058;
  assign n32060 = n32057 | n32058;
  assign n32061 = ~n32059 & n32060;
  assign n32062 = n56369 & n32061;
  assign n32063 = n56369 | n32061;
  assign n32064 = ~n32062 & n32063;
  assign n32065 = x125 & x223;
  assign n32066 = n32064 & n32065;
  assign n32067 = n32064 | n32065;
  assign n32068 = ~n32066 & n32067;
  assign n32069 = n56367 & n32068;
  assign n32070 = n56367 | n32068;
  assign n32071 = ~n32069 & n32070;
  assign n32072 = x124 & x224;
  assign n32073 = n32071 & n32072;
  assign n32074 = n32071 | n32072;
  assign n32075 = ~n32073 & n32074;
  assign n32076 = n56365 & n32075;
  assign n32077 = n56365 | n32075;
  assign n32078 = ~n32076 & n32077;
  assign n32079 = x123 & x225;
  assign n32080 = n32078 & n32079;
  assign n32081 = n32078 | n32079;
  assign n32082 = ~n32080 & n32081;
  assign n32083 = n31693 & n32082;
  assign n32084 = n31693 | n32082;
  assign n32085 = ~n32083 & n32084;
  assign n32086 = x122 & x226;
  assign n32087 = n32085 & n32086;
  assign n32088 = n32085 | n32086;
  assign n32089 = ~n32087 & n32088;
  assign n32090 = n31692 & n32089;
  assign n32091 = n31692 | n32089;
  assign n32092 = ~n32090 & n32091;
  assign n32093 = x121 & x227;
  assign n32094 = n32092 & n32093;
  assign n32095 = n32092 | n32093;
  assign n32096 = ~n32094 & n32095;
  assign n32097 = n70343 & n32096;
  assign n32098 = n70343 | n32096;
  assign n32099 = ~n32097 & n32098;
  assign n32100 = x120 & x228;
  assign n32101 = n32099 & n32100;
  assign n32102 = n32099 | n32100;
  assign n32103 = ~n32101 & n32102;
  assign n32104 = n56363 & n32103;
  assign n32105 = n56363 | n32103;
  assign n32106 = ~n32104 & n32105;
  assign n32107 = x119 & x229;
  assign n32108 = n32106 & n32107;
  assign n32109 = n32106 | n32107;
  assign n32110 = ~n32108 & n32109;
  assign n32111 = n56361 & n32110;
  assign n32112 = n56361 | n32110;
  assign n32113 = ~n32111 & n32112;
  assign n32114 = x118 & x230;
  assign n32115 = n32113 & n32114;
  assign n32116 = n32113 | n32114;
  assign n32117 = ~n32115 & n32116;
  assign n32118 = n56359 & n32117;
  assign n32119 = n56359 | n32117;
  assign n32120 = ~n32118 & n32119;
  assign n32121 = x117 & x231;
  assign n32122 = n32120 & n32121;
  assign n32123 = n32120 | n32121;
  assign n32124 = ~n32122 & n32123;
  assign n32125 = n56357 & n32124;
  assign n32126 = n56357 | n32124;
  assign n32127 = ~n32125 & n32126;
  assign n32128 = x116 & x232;
  assign n32129 = n32127 & n32128;
  assign n32130 = n32127 | n32128;
  assign n32131 = ~n32129 & n32130;
  assign n32132 = n56355 & n32131;
  assign n32133 = n56355 | n32131;
  assign n32134 = ~n32132 & n32133;
  assign n32135 = x115 & x233;
  assign n32136 = n32134 & n32135;
  assign n32137 = n32134 | n32135;
  assign n32138 = ~n32136 & n32137;
  assign n32139 = n56353 & n32138;
  assign n32140 = n56353 | n32138;
  assign n32141 = ~n32139 & n32140;
  assign n32142 = x114 & x234;
  assign n32143 = n32141 & n32142;
  assign n32144 = n32141 | n32142;
  assign n32145 = ~n32143 & n32144;
  assign n32146 = n56351 & n32145;
  assign n32147 = n56351 | n32145;
  assign n32148 = ~n32146 & n32147;
  assign n32149 = x113 & x235;
  assign n32150 = n32148 & n32149;
  assign n32151 = n32148 | n32149;
  assign n32152 = ~n32150 & n32151;
  assign n32153 = n31681 & n32152;
  assign n32154 = n31681 | n32152;
  assign n32155 = ~n32153 & n32154;
  assign n32156 = x112 & x236;
  assign n32157 = n32155 & n32156;
  assign n32158 = n32155 | n32156;
  assign n32159 = ~n32157 & n32158;
  assign n70488 = n31681 | n32149;
  assign n70489 = (n31681 & n32148) | (n31681 & n70488) | (n32148 & n70488);
  assign n56596 = (n32150 & n32152) | (n32150 & n70489) | (n32152 & n70489);
  assign n56597 = n32143 | n56351;
  assign n56598 = (n32143 & n32145) | (n32143 & n56597) | (n32145 & n56597);
  assign n56599 = n32136 | n56353;
  assign n56600 = (n32136 & n32138) | (n32136 & n56599) | (n32138 & n56599);
  assign n56601 = n32129 | n56355;
  assign n56602 = (n32129 & n32131) | (n32129 & n56601) | (n32131 & n56601);
  assign n56603 = n32122 | n56357;
  assign n56604 = (n32122 & n32124) | (n32122 & n56603) | (n32124 & n56603);
  assign n56605 = n32115 | n56359;
  assign n56606 = (n32115 & n32117) | (n32115 & n56605) | (n32117 & n56605);
  assign n56607 = n32108 | n56361;
  assign n56608 = (n32108 & n32110) | (n32108 & n56607) | (n32110 & n56607);
  assign n56609 = n32101 | n56363;
  assign n56610 = (n32101 & n32103) | (n32101 & n56609) | (n32103 & n56609);
  assign n70490 = n32094 | n70343;
  assign n70491 = (n32094 & n32096) | (n32094 & n70490) | (n32096 & n70490);
  assign n32169 = n32087 | n32090;
  assign n56611 = n32080 | n32082;
  assign n56612 = (n31693 & n32080) | (n31693 & n56611) | (n32080 & n56611);
  assign n56613 = n32073 | n32075;
  assign n56614 = (n32073 & n56365) | (n32073 & n56613) | (n56365 & n56613);
  assign n56615 = n32066 | n32068;
  assign n56616 = (n32066 & n56367) | (n32066 & n56615) | (n56367 & n56615);
  assign n56371 = (n31583 & n56128) | (n31583 & n56370) | (n56128 & n56370);
  assign n56373 = (n31576 & n56130) | (n31576 & n56372) | (n56130 & n56372);
  assign n56378 = (n70193 & n70345) | (n70193 & n56377) | (n70345 & n56377);
  assign n56626 = n31905 | n31907;
  assign n70492 = n31436 | n31905;
  assign n70493 = (n31905 & n31907) | (n31905 & n70492) | (n31907 & n70492);
  assign n70494 = (n56271 & n56626) | (n56271 & n70493) | (n56626 & n70493);
  assign n70495 = (n56270 & n56626) | (n56270 & n70493) | (n56626 & n70493);
  assign n70496 = (n55911 & n70494) | (n55911 & n70495) | (n70494 & n70495);
  assign n56631 = n31884 | n31886;
  assign n70497 = n31415 | n31884;
  assign n70498 = (n31884 & n31886) | (n31884 & n70497) | (n31886 & n70497);
  assign n70499 = (n56261 & n56631) | (n56261 & n70498) | (n56631 & n70498);
  assign n70500 = (n56260 & n56631) | (n56260 & n70498) | (n56631 & n70498);
  assign n70501 = (n70103 & n70499) | (n70103 & n70500) | (n70499 & n70500);
  assign n70508 = n31338 | n31807;
  assign n70509 = (n31807 & n31809) | (n31807 & n70508) | (n31809 & n70508);
  assign n70510 = n31807 | n31809;
  assign n70511 = (n31807 & n56402) | (n31807 & n70510) | (n56402 & n70510);
  assign n70512 = (n56160 & n70509) | (n56160 & n70511) | (n70509 & n70511);
  assign n70513 = (n70228 & n70509) | (n70228 & n70511) | (n70509 & n70511);
  assign n70514 = (n69994 & n70512) | (n69994 & n70513) | (n70512 & n70513);
  assign n32219 = x173 & x176;
  assign n32220 = x172 & x177;
  assign n32221 = n32219 & n32220;
  assign n32222 = n32219 | n32220;
  assign n32223 = ~n32221 & n32222;
  assign n70525 = n31744 & n32223;
  assign n70526 = (n32223 & n70383) | (n32223 & n70525) | (n70383 & n70525);
  assign n70527 = n31744 | n70384;
  assign n70530 = n32223 & n70527;
  assign n70528 = n31744 | n31746;
  assign n70531 = n32223 & n70528;
  assign n70532 = (n70244 & n70530) | (n70244 & n70531) | (n70530 & n70531);
  assign n70533 = (n69747 & n70526) | (n69747 & n70532) | (n70526 & n70532);
  assign n70534 = (n69746 & n70526) | (n69746 & n70532) | (n70526 & n70532);
  assign n70535 = (n68195 & n70533) | (n68195 & n70534) | (n70533 & n70534);
  assign n70536 = n31744 | n32223;
  assign n70537 = n70383 | n70536;
  assign n70538 = n32223 | n70527;
  assign n70539 = n32223 | n70528;
  assign n70540 = (n70244 & n70538) | (n70244 & n70539) | (n70538 & n70539);
  assign n70541 = (n69747 & n70537) | (n69747 & n70540) | (n70537 & n70540);
  assign n70542 = (n69746 & n70537) | (n69746 & n70540) | (n70537 & n70540);
  assign n70543 = (n68195 & n70541) | (n68195 & n70542) | (n70541 & n70542);
  assign n32226 = ~n70535 & n70543;
  assign n32227 = x171 & x178;
  assign n32228 = n32226 & n32227;
  assign n32229 = n32226 | n32227;
  assign n32230 = ~n32228 & n32229;
  assign n56678 = n31751 & n32230;
  assign n70544 = (n32230 & n56678) | (n32230 & n70398) | (n56678 & n70398);
  assign n70545 = (n32230 & n56678) | (n32230 & n70402) | (n56678 & n70402);
  assign n70546 = (n69887 & n70544) | (n69887 & n70545) | (n70544 & n70545);
  assign n56680 = n31751 | n32230;
  assign n70547 = n56680 | n70398;
  assign n70548 = n56680 | n70402;
  assign n70549 = (n69887 & n70547) | (n69887 & n70548) | (n70547 & n70548);
  assign n32233 = ~n70546 & n70549;
  assign n32234 = x170 & x179;
  assign n32235 = n32233 & n32234;
  assign n32236 = n32233 | n32234;
  assign n32237 = ~n32235 & n32236;
  assign n70522 = n31758 | n31760;
  assign n70524 = (n31758 & n70409) | (n31758 & n70522) | (n70409 & n70522);
  assign n70550 = n32237 & n70524;
  assign n70523 = (n31758 & n70408) | (n31758 & n70522) | (n70408 & n70522);
  assign n70551 = n32237 & n70523;
  assign n70552 = (n70013 & n70550) | (n70013 & n70551) | (n70550 & n70551);
  assign n70553 = n32237 | n70524;
  assign n70554 = n32237 | n70523;
  assign n70555 = (n70013 & n70553) | (n70013 & n70554) | (n70553 & n70554);
  assign n32240 = ~n70552 & n70555;
  assign n32241 = x169 & x180;
  assign n32242 = n32240 & n32241;
  assign n32243 = n32240 | n32241;
  assign n32244 = ~n32242 & n32243;
  assign n70519 = n31765 | n31767;
  assign n70520 = (n31765 & n70411) | (n31765 & n70519) | (n70411 & n70519);
  assign n70556 = n32244 & n70520;
  assign n70521 = (n31765 & n70413) | (n31765 & n70519) | (n70413 & n70519);
  assign n70557 = n32244 & n70521;
  assign n70558 = (n70133 & n70556) | (n70133 & n70557) | (n70556 & n70557);
  assign n70559 = n32244 | n70520;
  assign n70560 = n32244 | n70521;
  assign n70561 = (n70133 & n70559) | (n70133 & n70560) | (n70559 & n70560);
  assign n32247 = ~n70558 & n70561;
  assign n32248 = x168 & x181;
  assign n32249 = n32247 & n32248;
  assign n32250 = n32247 | n32248;
  assign n32251 = ~n32249 & n32250;
  assign n56661 = n31772 | n31774;
  assign n56682 = n32251 & n56661;
  assign n56683 = n31772 & n32251;
  assign n70562 = (n56682 & n56683) | (n56682 & n70376) | (n56683 & n70376);
  assign n70563 = (n56682 & n56683) | (n56682 & n70375) | (n56683 & n70375);
  assign n70564 = (n69736 & n70562) | (n69736 & n70563) | (n70562 & n70563);
  assign n56685 = n32251 | n56661;
  assign n56686 = n31772 | n32251;
  assign n70565 = (n56685 & n56686) | (n56685 & n70376) | (n56686 & n70376);
  assign n70566 = (n56685 & n56686) | (n56685 & n70375) | (n56686 & n70375);
  assign n70567 = (n69736 & n70565) | (n69736 & n70566) | (n70565 & n70566);
  assign n32254 = ~n70564 & n70567;
  assign n32255 = x167 & x182;
  assign n32256 = n32254 & n32255;
  assign n32257 = n32254 | n32255;
  assign n32258 = ~n32256 & n32257;
  assign n70568 = n31779 | n31781;
  assign n70569 = (n31779 & n56412) | (n31779 & n70568) | (n56412 & n70568);
  assign n56688 = n32258 & n70569;
  assign n70570 = n31310 | n31779;
  assign n70571 = (n31779 & n31781) | (n31779 & n70570) | (n31781 & n70570);
  assign n56689 = n32258 & n70571;
  assign n70572 = (n56688 & n56689) | (n56688 & n70238) | (n56689 & n70238);
  assign n70573 = (n56688 & n56689) | (n56688 & n70237) | (n56689 & n70237);
  assign n70574 = (n69916 & n70572) | (n69916 & n70573) | (n70572 & n70573);
  assign n56691 = n32258 | n70569;
  assign n56692 = n32258 | n70571;
  assign n70575 = (n56691 & n56692) | (n56691 & n70238) | (n56692 & n70238);
  assign n70576 = (n56691 & n56692) | (n56691 & n70237) | (n56692 & n70237);
  assign n70577 = (n69916 & n70575) | (n69916 & n70576) | (n70575 & n70576);
  assign n32261 = ~n70574 & n70577;
  assign n32262 = x166 & x183;
  assign n32263 = n32261 & n32262;
  assign n32264 = n32261 | n32262;
  assign n32265 = ~n32263 & n32264;
  assign n56694 = n31786 & n32265;
  assign n56695 = (n32265 & n70430) | (n32265 & n56694) | (n70430 & n56694);
  assign n56696 = n31786 | n32265;
  assign n56697 = n70430 | n56696;
  assign n32268 = ~n56695 & n56697;
  assign n32269 = x165 & x184;
  assign n32270 = n32268 & n32269;
  assign n32271 = n32268 | n32269;
  assign n32272 = ~n32270 & n32271;
  assign n70515 = n31793 | n31795;
  assign n70516 = (n31793 & n56407) | (n31793 & n70515) | (n56407 & n70515);
  assign n70578 = n32272 & n70516;
  assign n70517 = n31324 | n31793;
  assign n70518 = (n31793 & n31795) | (n31793 & n70517) | (n31795 & n70517);
  assign n70579 = n32272 & n70518;
  assign n70580 = (n70235 & n70578) | (n70235 & n70579) | (n70578 & n70579);
  assign n70581 = n32272 | n70516;
  assign n70582 = n32272 | n70518;
  assign n70583 = (n70235 & n70581) | (n70235 & n70582) | (n70581 & n70582);
  assign n32275 = ~n70580 & n70583;
  assign n32276 = x164 & x185;
  assign n32277 = n32275 & n32276;
  assign n32278 = n32275 | n32276;
  assign n32279 = ~n32277 & n32278;
  assign n56653 = n31800 | n31802;
  assign n56698 = n32279 & n56653;
  assign n56699 = n31800 & n32279;
  assign n70584 = (n56405 & n56698) | (n56405 & n56699) | (n56698 & n56699);
  assign n70585 = (n56698 & n56699) | (n56698 & n70371) | (n56699 & n70371);
  assign n70586 = (n70127 & n70584) | (n70127 & n70585) | (n70584 & n70585);
  assign n56701 = n32279 | n56653;
  assign n56702 = n31800 | n32279;
  assign n70587 = (n56405 & n56701) | (n56405 & n56702) | (n56701 & n56702);
  assign n70588 = (n56701 & n56702) | (n56701 & n70371) | (n56702 & n70371);
  assign n70589 = (n70127 & n70587) | (n70127 & n70588) | (n70587 & n70588);
  assign n32282 = ~n70586 & n70589;
  assign n32283 = x163 & x186;
  assign n32284 = n32282 & n32283;
  assign n32285 = n32282 | n32283;
  assign n32286 = ~n32284 & n32285;
  assign n32287 = n70514 & n32286;
  assign n32288 = n70514 | n32286;
  assign n32289 = ~n32287 & n32288;
  assign n32290 = x162 & x187;
  assign n32291 = n32289 & n32290;
  assign n32292 = n32289 | n32290;
  assign n32293 = ~n32291 & n32292;
  assign n56648 = n31814 | n31816;
  assign n56704 = n32293 & n56648;
  assign n56705 = n31814 & n32293;
  assign n70590 = (n56704 & n56705) | (n56704 & n70369) | (n56705 & n70369);
  assign n70591 = (n56704 & n56705) | (n56704 & n70367) | (n56705 & n70367);
  assign n70592 = (n55934 & n70590) | (n55934 & n70591) | (n70590 & n70591);
  assign n56707 = n32293 | n56648;
  assign n56708 = n31814 | n32293;
  assign n70593 = (n56707 & n56708) | (n56707 & n70369) | (n56708 & n70369);
  assign n70594 = (n56707 & n56708) | (n56707 & n70367) | (n56708 & n70367);
  assign n70595 = (n55934 & n70593) | (n55934 & n70594) | (n70593 & n70594);
  assign n32296 = ~n70592 & n70595;
  assign n32297 = x161 & x188;
  assign n32298 = n32296 & n32297;
  assign n32299 = n32296 | n32297;
  assign n32300 = ~n32298 & n32299;
  assign n56646 = n31821 | n31823;
  assign n70596 = n32300 & n56646;
  assign n70506 = n31352 | n31821;
  assign n70507 = (n31821 & n31823) | (n31821 & n70506) | (n31823 & n70506);
  assign n70597 = n32300 & n70507;
  assign n70598 = (n56232 & n70596) | (n56232 & n70597) | (n70596 & n70597);
  assign n70599 = n32300 | n56646;
  assign n70600 = n32300 | n70507;
  assign n70601 = (n56232 & n70599) | (n56232 & n70600) | (n70599 & n70600);
  assign n32303 = ~n70598 & n70601;
  assign n32304 = x160 & x189;
  assign n32305 = n32303 & n32304;
  assign n32306 = n32303 | n32304;
  assign n32307 = ~n32305 & n32306;
  assign n56643 = n31828 | n31830;
  assign n56710 = n32307 & n56643;
  assign n56711 = n31828 & n32307;
  assign n56712 = (n70365 & n56710) | (n70365 & n56711) | (n56710 & n56711);
  assign n56713 = n32307 | n56643;
  assign n56714 = n31828 | n32307;
  assign n56715 = (n70365 & n56713) | (n70365 & n56714) | (n56713 & n56714);
  assign n32310 = ~n56712 & n56715;
  assign n32311 = x159 & x190;
  assign n32312 = n32310 & n32311;
  assign n32313 = n32310 | n32311;
  assign n32314 = ~n32312 & n32313;
  assign n56716 = n31835 & n32314;
  assign n70602 = (n32314 & n56482) | (n32314 & n56716) | (n56482 & n56716);
  assign n70603 = (n32314 & n56481) | (n32314 & n56716) | (n56481 & n56716);
  assign n70604 = (n56154 & n70602) | (n56154 & n70603) | (n70602 & n70603);
  assign n56718 = n31835 | n32314;
  assign n70605 = n56482 | n56718;
  assign n70606 = n56481 | n56718;
  assign n70607 = (n56154 & n70605) | (n56154 & n70606) | (n70605 & n70606);
  assign n32317 = ~n70604 & n70607;
  assign n32318 = x158 & x191;
  assign n32319 = n32317 & n32318;
  assign n32320 = n32317 | n32318;
  assign n32321 = ~n32319 & n32320;
  assign n56641 = n31842 | n31844;
  assign n70608 = n32321 & n56641;
  assign n70504 = n31373 | n31842;
  assign n70505 = (n31842 & n31844) | (n31842 & n70504) | (n31844 & n70504);
  assign n70609 = n32321 & n70505;
  assign n70610 = (n56242 & n70608) | (n56242 & n70609) | (n70608 & n70609);
  assign n70611 = n32321 | n56641;
  assign n70612 = n32321 | n70505;
  assign n70613 = (n56242 & n70611) | (n56242 & n70612) | (n70611 & n70612);
  assign n32324 = ~n70610 & n70613;
  assign n32325 = x157 & x192;
  assign n32326 = n32324 & n32325;
  assign n32327 = n32324 | n32325;
  assign n32328 = ~n32326 & n32327;
  assign n56638 = n31849 | n31851;
  assign n56720 = n32328 & n56638;
  assign n56721 = n31849 & n32328;
  assign n56722 = (n70360 & n56720) | (n70360 & n56721) | (n56720 & n56721);
  assign n56723 = n32328 | n56638;
  assign n56724 = n31849 | n32328;
  assign n56725 = (n70360 & n56723) | (n70360 & n56724) | (n56723 & n56724);
  assign n32331 = ~n56722 & n56725;
  assign n32332 = x156 & x193;
  assign n32333 = n32331 & n32332;
  assign n32334 = n32331 | n32332;
  assign n32335 = ~n32333 & n32334;
  assign n56726 = n31856 & n32335;
  assign n70614 = (n32335 & n56492) | (n32335 & n56726) | (n56492 & n56726);
  assign n70615 = (n32335 & n56491) | (n32335 & n56726) | (n56491 & n56726);
  assign n70616 = (n56149 & n70614) | (n56149 & n70615) | (n70614 & n70615);
  assign n56728 = n31856 | n32335;
  assign n70617 = n56492 | n56728;
  assign n70618 = n56491 | n56728;
  assign n70619 = (n56149 & n70617) | (n56149 & n70618) | (n70617 & n70618);
  assign n32338 = ~n70616 & n70619;
  assign n32339 = x155 & x194;
  assign n32340 = n32338 & n32339;
  assign n32341 = n32338 | n32339;
  assign n32342 = ~n32340 & n32341;
  assign n56636 = n31863 | n31865;
  assign n70620 = n32342 & n56636;
  assign n70502 = n31394 | n31863;
  assign n70503 = (n31863 & n31865) | (n31863 & n70502) | (n31865 & n70502);
  assign n70621 = n32342 & n70503;
  assign n70622 = (n56252 & n70620) | (n56252 & n70621) | (n70620 & n70621);
  assign n70623 = n32342 | n56636;
  assign n70624 = n32342 | n70503;
  assign n70625 = (n56252 & n70623) | (n56252 & n70624) | (n70623 & n70624);
  assign n32345 = ~n70622 & n70625;
  assign n32346 = x154 & x195;
  assign n32347 = n32345 & n32346;
  assign n32348 = n32345 | n32346;
  assign n32349 = ~n32347 & n32348;
  assign n56633 = n31870 | n31872;
  assign n56730 = n32349 & n56633;
  assign n56731 = n31870 & n32349;
  assign n56732 = (n70355 & n56730) | (n70355 & n56731) | (n56730 & n56731);
  assign n56733 = n32349 | n56633;
  assign n56734 = n31870 | n32349;
  assign n56735 = (n70355 & n56733) | (n70355 & n56734) | (n56733 & n56734);
  assign n32352 = ~n56732 & n56735;
  assign n32353 = x153 & x196;
  assign n32354 = n32352 & n32353;
  assign n32355 = n32352 | n32353;
  assign n32356 = ~n32354 & n32355;
  assign n56736 = n31877 & n32356;
  assign n70626 = (n32356 & n56502) | (n32356 & n56736) | (n56502 & n56736);
  assign n70627 = (n32356 & n56501) | (n32356 & n56736) | (n56501 & n56736);
  assign n70628 = (n70222 & n70626) | (n70222 & n70627) | (n70626 & n70627);
  assign n56738 = n31877 | n32356;
  assign n70629 = n56502 | n56738;
  assign n70630 = n56501 | n56738;
  assign n70631 = (n70222 & n70629) | (n70222 & n70630) | (n70629 & n70630);
  assign n32359 = ~n70628 & n70631;
  assign n32360 = x152 & x197;
  assign n32361 = n32359 & n32360;
  assign n32362 = n32359 | n32360;
  assign n32363 = ~n32361 & n32362;
  assign n32364 = n70501 & n32363;
  assign n32365 = n70501 | n32363;
  assign n32366 = ~n32364 & n32365;
  assign n32367 = x151 & x198;
  assign n32368 = n32366 & n32367;
  assign n32369 = n32366 | n32367;
  assign n32370 = ~n32368 & n32369;
  assign n56628 = n31891 | n31893;
  assign n56740 = n32370 & n56628;
  assign n56741 = n31891 & n32370;
  assign n56742 = (n70350 & n56740) | (n70350 & n56741) | (n56740 & n56741);
  assign n56743 = n32370 | n56628;
  assign n56744 = n31891 | n32370;
  assign n56745 = (n70350 & n56743) | (n70350 & n56744) | (n56743 & n56744);
  assign n32373 = ~n56742 & n56745;
  assign n32374 = x150 & x199;
  assign n32375 = n32373 & n32374;
  assign n32376 = n32373 | n32374;
  assign n32377 = ~n32375 & n32376;
  assign n56746 = n31898 & n32377;
  assign n70632 = (n32377 & n56512) | (n32377 & n56746) | (n56512 & n56746);
  assign n70633 = (n32377 & n56511) | (n32377 & n56746) | (n56511 & n56746);
  assign n70634 = (n70217 & n70632) | (n70217 & n70633) | (n70632 & n70633);
  assign n56748 = n31898 | n32377;
  assign n70635 = n56512 | n56748;
  assign n70636 = n56511 | n56748;
  assign n70637 = (n70217 & n70635) | (n70217 & n70636) | (n70635 & n70636);
  assign n32380 = ~n70634 & n70637;
  assign n32381 = x149 & x200;
  assign n32382 = n32380 & n32381;
  assign n32383 = n32380 | n32381;
  assign n32384 = ~n32382 & n32383;
  assign n32385 = n70496 & n32384;
  assign n32386 = n70496 | n32384;
  assign n32387 = ~n32385 & n32386;
  assign n32388 = x148 & x201;
  assign n32389 = n32387 & n32388;
  assign n32390 = n32387 | n32388;
  assign n32391 = ~n32389 & n32390;
  assign n56623 = n31912 | n31914;
  assign n56750 = n32391 & n56623;
  assign n56751 = n31912 & n32391;
  assign n56752 = (n56378 & n56750) | (n56378 & n56751) | (n56750 & n56751);
  assign n56753 = n32391 | n56623;
  assign n56754 = n31912 | n32391;
  assign n56755 = (n56378 & n56753) | (n56378 & n56754) | (n56753 & n56754);
  assign n32394 = ~n56752 & n56755;
  assign n32395 = x147 & x202;
  assign n32396 = n32394 & n32395;
  assign n32397 = n32394 | n32395;
  assign n32398 = ~n32396 & n32397;
  assign n56756 = n31919 & n32398;
  assign n56757 = (n32398 & n70472) | (n32398 & n56756) | (n70472 & n56756);
  assign n56758 = n31919 | n32398;
  assign n56759 = n70472 | n56758;
  assign n32401 = ~n56757 & n56759;
  assign n32402 = x146 & x203;
  assign n32403 = n32401 & n32402;
  assign n32404 = n32401 | n32402;
  assign n32405 = ~n32403 & n32404;
  assign n56760 = n31926 & n32405;
  assign n56761 = (n32405 & n56526) | (n32405 & n56760) | (n56526 & n56760);
  assign n56762 = n31926 | n32405;
  assign n56763 = n56526 | n56762;
  assign n32408 = ~n56761 & n56763;
  assign n32409 = x145 & x204;
  assign n32410 = n32408 & n32409;
  assign n32411 = n32408 | n32409;
  assign n32412 = ~n32410 & n32411;
  assign n56764 = n31933 & n32412;
  assign n56765 = (n32412 & n56530) | (n32412 & n56764) | (n56530 & n56764);
  assign n56766 = n31933 | n32412;
  assign n56767 = n56530 | n56766;
  assign n32415 = ~n56765 & n56767;
  assign n32416 = x144 & x205;
  assign n32417 = n32415 & n32416;
  assign n32418 = n32415 | n32416;
  assign n32419 = ~n32417 & n32418;
  assign n56768 = n31940 & n32419;
  assign n56769 = (n32419 & n56534) | (n32419 & n56768) | (n56534 & n56768);
  assign n56770 = n31940 | n32419;
  assign n56771 = n56534 | n56770;
  assign n32422 = ~n56769 & n56771;
  assign n32423 = x143 & x206;
  assign n32424 = n32422 & n32423;
  assign n32425 = n32422 | n32423;
  assign n32426 = ~n32424 & n32425;
  assign n56772 = n31947 & n32426;
  assign n56773 = (n32426 & n56538) | (n32426 & n56772) | (n56538 & n56772);
  assign n56774 = n31947 | n32426;
  assign n56775 = n56538 | n56774;
  assign n32429 = ~n56773 & n56775;
  assign n32430 = x142 & x207;
  assign n32431 = n32429 & n32430;
  assign n32432 = n32429 | n32430;
  assign n32433 = ~n32431 & n32432;
  assign n56776 = n31954 & n32433;
  assign n56777 = (n32433 & n56542) | (n32433 & n56776) | (n56542 & n56776);
  assign n56778 = n31954 | n32433;
  assign n56779 = n56542 | n56778;
  assign n32436 = ~n56777 & n56779;
  assign n32437 = x141 & x208;
  assign n32438 = n32436 & n32437;
  assign n32439 = n32436 | n32437;
  assign n32440 = ~n32438 & n32439;
  assign n56780 = n31961 & n32440;
  assign n56781 = (n32440 & n56546) | (n32440 & n56780) | (n56546 & n56780);
  assign n56782 = n31961 | n32440;
  assign n56783 = n56546 | n56782;
  assign n32443 = ~n56781 & n56783;
  assign n32444 = x140 & x209;
  assign n32445 = n32443 & n32444;
  assign n32446 = n32443 | n32444;
  assign n32447 = ~n32445 & n32446;
  assign n56784 = n31968 & n32447;
  assign n56785 = (n32447 & n56550) | (n32447 & n56784) | (n56550 & n56784);
  assign n56786 = n31968 | n32447;
  assign n56787 = n56550 | n56786;
  assign n32450 = ~n56785 & n56787;
  assign n32451 = x139 & x210;
  assign n32452 = n32450 & n32451;
  assign n32453 = n32450 | n32451;
  assign n32454 = ~n32452 & n32453;
  assign n56788 = n31975 & n32454;
  assign n56789 = (n32454 & n56554) | (n32454 & n56788) | (n56554 & n56788);
  assign n56790 = n31975 | n32454;
  assign n56791 = n56554 | n56790;
  assign n32457 = ~n56789 & n56791;
  assign n32458 = x138 & x211;
  assign n32459 = n32457 & n32458;
  assign n32460 = n32457 | n32458;
  assign n32461 = ~n32459 & n32460;
  assign n56792 = n31982 & n32461;
  assign n56793 = (n32461 & n56558) | (n32461 & n56792) | (n56558 & n56792);
  assign n56794 = n31982 | n32461;
  assign n56795 = n56558 | n56794;
  assign n32464 = ~n56793 & n56795;
  assign n32465 = x137 & x212;
  assign n32466 = n32464 & n32465;
  assign n32467 = n32464 | n32465;
  assign n32468 = ~n32466 & n32467;
  assign n56796 = n31989 & n32468;
  assign n56797 = (n32468 & n56562) | (n32468 & n56796) | (n56562 & n56796);
  assign n56798 = n31989 | n32468;
  assign n56799 = n56562 | n56798;
  assign n32471 = ~n56797 & n56799;
  assign n32472 = x136 & x213;
  assign n32473 = n32471 & n32472;
  assign n32474 = n32471 | n32472;
  assign n32475 = ~n32473 & n32474;
  assign n56800 = n31996 & n32475;
  assign n56801 = (n32475 & n56566) | (n32475 & n56800) | (n56566 & n56800);
  assign n56802 = n31996 | n32475;
  assign n56803 = n56566 | n56802;
  assign n32478 = ~n56801 & n56803;
  assign n32479 = x135 & x214;
  assign n32480 = n32478 & n32479;
  assign n32481 = n32478 | n32479;
  assign n32482 = ~n32480 & n32481;
  assign n56804 = n32003 & n32482;
  assign n56805 = (n32482 & n56570) | (n32482 & n56804) | (n56570 & n56804);
  assign n56806 = n32003 | n32482;
  assign n56807 = n56570 | n56806;
  assign n32485 = ~n56805 & n56807;
  assign n32486 = x134 & x215;
  assign n32487 = n32485 & n32486;
  assign n32488 = n32485 | n32486;
  assign n32489 = ~n32487 & n32488;
  assign n56808 = n32010 & n32489;
  assign n56809 = (n32489 & n56574) | (n32489 & n56808) | (n56574 & n56808);
  assign n56810 = n32010 | n32489;
  assign n56811 = n56574 | n56810;
  assign n32492 = ~n56809 & n56811;
  assign n32493 = x133 & x216;
  assign n32494 = n32492 & n32493;
  assign n32495 = n32492 | n32493;
  assign n32496 = ~n32494 & n32495;
  assign n56812 = n32017 & n32496;
  assign n56813 = (n32496 & n56578) | (n32496 & n56812) | (n56578 & n56812);
  assign n56814 = n32017 | n32496;
  assign n56815 = n56578 | n56814;
  assign n32499 = ~n56813 & n56815;
  assign n32500 = x132 & x217;
  assign n32501 = n32499 & n32500;
  assign n32502 = n32499 | n32500;
  assign n32503 = ~n32501 & n32502;
  assign n56816 = n32024 & n32503;
  assign n56817 = (n32503 & n56582) | (n32503 & n56816) | (n56582 & n56816);
  assign n56818 = n32024 | n32503;
  assign n56819 = n56582 | n56818;
  assign n32506 = ~n56817 & n56819;
  assign n32507 = x131 & x218;
  assign n32508 = n32506 & n32507;
  assign n32509 = n32506 | n32507;
  assign n32510 = ~n32508 & n32509;
  assign n56820 = n32031 & n32510;
  assign n56821 = (n32510 & n56586) | (n32510 & n56820) | (n56586 & n56820);
  assign n56822 = n32031 | n32510;
  assign n56823 = n56586 | n56822;
  assign n32513 = ~n56821 & n56823;
  assign n32514 = x130 & x219;
  assign n32515 = n32513 & n32514;
  assign n32516 = n32513 | n32514;
  assign n32517 = ~n32515 & n32516;
  assign n56824 = n32038 & n32517;
  assign n56825 = (n32517 & n56591) | (n32517 & n56824) | (n56591 & n56824);
  assign n56826 = n32038 | n32517;
  assign n56827 = n56591 | n56826;
  assign n32520 = ~n56825 & n56827;
  assign n32521 = x129 & x220;
  assign n32522 = n32520 & n32521;
  assign n32523 = n32520 | n32521;
  assign n32524 = ~n32522 & n32523;
  assign n56621 = n32045 | n32047;
  assign n56828 = n32524 & n56621;
  assign n56829 = n32045 & n32524;
  assign n56830 = (n56373 & n56828) | (n56373 & n56829) | (n56828 & n56829);
  assign n56831 = n32524 | n56621;
  assign n56832 = n32045 | n32524;
  assign n56833 = (n56373 & n56831) | (n56373 & n56832) | (n56831 & n56832);
  assign n32527 = ~n56830 & n56833;
  assign n32528 = x128 & x221;
  assign n32529 = n32527 & n32528;
  assign n32530 = n32527 | n32528;
  assign n32531 = ~n32529 & n32530;
  assign n56619 = n32052 | n32054;
  assign n70638 = n32531 & n56619;
  assign n70639 = n32052 & n32531;
  assign n70640 = (n56371 & n70638) | (n56371 & n70639) | (n70638 & n70639);
  assign n70641 = n32531 | n56619;
  assign n70642 = n32052 | n32531;
  assign n70643 = (n56371 & n70641) | (n56371 & n70642) | (n70641 & n70642);
  assign n32534 = ~n70640 & n70643;
  assign n32535 = x127 & x222;
  assign n32536 = n32534 & n32535;
  assign n32537 = n32534 | n32535;
  assign n32538 = ~n32536 & n32537;
  assign n56617 = n32059 | n32061;
  assign n70644 = n32538 & n56617;
  assign n70645 = n32059 & n32538;
  assign n70646 = (n56369 & n70644) | (n56369 & n70645) | (n70644 & n70645);
  assign n70647 = n32538 | n56617;
  assign n70648 = n32059 | n32538;
  assign n70649 = (n56369 & n70647) | (n56369 & n70648) | (n70647 & n70648);
  assign n32541 = ~n70646 & n70649;
  assign n32542 = x126 & x223;
  assign n32543 = n32541 & n32542;
  assign n32544 = n32541 | n32542;
  assign n32545 = ~n32543 & n32544;
  assign n32546 = n56616 & n32545;
  assign n32547 = n56616 | n32545;
  assign n32548 = ~n32546 & n32547;
  assign n32549 = x125 & x224;
  assign n32550 = n32548 & n32549;
  assign n32551 = n32548 | n32549;
  assign n32552 = ~n32550 & n32551;
  assign n32553 = n56614 & n32552;
  assign n32554 = n56614 | n32552;
  assign n32555 = ~n32553 & n32554;
  assign n32556 = x124 & x225;
  assign n32557 = n32555 & n32556;
  assign n32558 = n32555 | n32556;
  assign n32559 = ~n32557 & n32558;
  assign n32560 = n56612 & n32559;
  assign n32561 = n56612 | n32559;
  assign n32562 = ~n32560 & n32561;
  assign n32563 = x123 & x226;
  assign n32564 = n32562 & n32563;
  assign n32565 = n32562 | n32563;
  assign n32566 = ~n32564 & n32565;
  assign n32567 = n32169 & n32566;
  assign n32568 = n32169 | n32566;
  assign n32569 = ~n32567 & n32568;
  assign n32570 = x122 & x227;
  assign n32571 = n32569 & n32570;
  assign n32572 = n32569 | n32570;
  assign n32573 = ~n32571 & n32572;
  assign n32574 = n70491 & n32573;
  assign n32575 = n70491 | n32573;
  assign n32576 = ~n32574 & n32575;
  assign n32577 = x121 & x228;
  assign n32578 = n32576 & n32577;
  assign n32579 = n32576 | n32577;
  assign n32580 = ~n32578 & n32579;
  assign n32581 = n56610 & n32580;
  assign n32582 = n56610 | n32580;
  assign n32583 = ~n32581 & n32582;
  assign n32584 = x120 & x229;
  assign n32585 = n32583 & n32584;
  assign n32586 = n32583 | n32584;
  assign n32587 = ~n32585 & n32586;
  assign n32588 = n56608 & n32587;
  assign n32589 = n56608 | n32587;
  assign n32590 = ~n32588 & n32589;
  assign n32591 = x119 & x230;
  assign n32592 = n32590 & n32591;
  assign n32593 = n32590 | n32591;
  assign n32594 = ~n32592 & n32593;
  assign n32595 = n56606 & n32594;
  assign n32596 = n56606 | n32594;
  assign n32597 = ~n32595 & n32596;
  assign n32598 = x118 & x231;
  assign n32599 = n32597 & n32598;
  assign n32600 = n32597 | n32598;
  assign n32601 = ~n32599 & n32600;
  assign n32602 = n56604 & n32601;
  assign n32603 = n56604 | n32601;
  assign n32604 = ~n32602 & n32603;
  assign n32605 = x117 & x232;
  assign n32606 = n32604 & n32605;
  assign n32607 = n32604 | n32605;
  assign n32608 = ~n32606 & n32607;
  assign n32609 = n56602 & n32608;
  assign n32610 = n56602 | n32608;
  assign n32611 = ~n32609 & n32610;
  assign n32612 = x116 & x233;
  assign n32613 = n32611 & n32612;
  assign n32614 = n32611 | n32612;
  assign n32615 = ~n32613 & n32614;
  assign n32616 = n56600 & n32615;
  assign n32617 = n56600 | n32615;
  assign n32618 = ~n32616 & n32617;
  assign n32619 = x115 & x234;
  assign n32620 = n32618 & n32619;
  assign n32621 = n32618 | n32619;
  assign n32622 = ~n32620 & n32621;
  assign n32623 = n56598 & n32622;
  assign n32624 = n56598 | n32622;
  assign n32625 = ~n32623 & n32624;
  assign n32626 = x114 & x235;
  assign n32627 = n32625 & n32626;
  assign n32628 = n32625 | n32626;
  assign n32629 = ~n32627 & n32628;
  assign n32630 = n56596 & n32629;
  assign n32631 = n56596 | n32629;
  assign n32632 = ~n32630 & n32631;
  assign n32633 = x113 & x236;
  assign n32634 = n32632 & n32633;
  assign n32635 = n32632 | n32633;
  assign n32636 = ~n32634 & n32635;
  assign n32637 = n32157 & n32636;
  assign n32638 = n32157 | n32636;
  assign n32639 = ~n32637 & n32638;
  assign n32640 = x112 & x237;
  assign n32641 = n32639 & n32640;
  assign n32642 = n32639 | n32640;
  assign n32643 = ~n32641 & n32642;
  assign n70650 = n32157 | n32633;
  assign n70651 = (n32157 & n32632) | (n32157 & n70650) | (n32632 & n70650);
  assign n56835 = (n32634 & n32636) | (n32634 & n70651) | (n32636 & n70651);
  assign n56836 = n32627 | n56596;
  assign n56837 = (n32627 & n32629) | (n32627 & n56836) | (n32629 & n56836);
  assign n56838 = n32620 | n56598;
  assign n56839 = (n32620 & n32622) | (n32620 & n56838) | (n32622 & n56838);
  assign n56840 = n32613 | n56600;
  assign n56841 = (n32613 & n32615) | (n32613 & n56840) | (n32615 & n56840);
  assign n56842 = n32606 | n56602;
  assign n56843 = (n32606 & n32608) | (n32606 & n56842) | (n32608 & n56842);
  assign n56844 = n32599 | n56604;
  assign n56845 = (n32599 & n32601) | (n32599 & n56844) | (n32601 & n56844);
  assign n56846 = n32592 | n56606;
  assign n56847 = (n32592 & n32594) | (n32592 & n56846) | (n32594 & n56846);
  assign n56848 = n32585 | n56608;
  assign n56849 = (n32585 & n32587) | (n32585 & n56848) | (n32587 & n56848);
  assign n56850 = n32578 | n56610;
  assign n56851 = (n32578 & n32580) | (n32578 & n56850) | (n32580 & n56850);
  assign n70652 = n32571 | n70491;
  assign n70653 = (n32571 & n32573) | (n32571 & n70652) | (n32573 & n70652);
  assign n56852 = n32564 | n32566;
  assign n56853 = (n32169 & n32564) | (n32169 & n56852) | (n32564 & n56852);
  assign n56854 = n32557 | n32559;
  assign n56855 = (n32557 & n56612) | (n32557 & n56854) | (n56612 & n56854);
  assign n56856 = n32550 | n32552;
  assign n56857 = (n32550 & n56614) | (n32550 & n56856) | (n56614 & n56856);
  assign n56618 = (n32059 & n56369) | (n32059 & n56617) | (n56369 & n56617);
  assign n56620 = (n32052 & n56371) | (n32052 & n56619) | (n56371 & n56619);
  assign n56870 = n32375 | n32377;
  assign n70656 = n31898 | n32375;
  assign n70657 = (n32375 & n32377) | (n32375 & n70656) | (n32377 & n70656);
  assign n70658 = (n56512 & n56870) | (n56512 & n70657) | (n56870 & n70657);
  assign n70659 = (n56511 & n56870) | (n56511 & n70657) | (n56870 & n70657);
  assign n70660 = (n70217 & n70658) | (n70217 & n70659) | (n70658 & n70659);
  assign n56875 = n32354 | n32356;
  assign n70661 = n31877 | n32354;
  assign n70662 = (n32354 & n32356) | (n32354 & n70661) | (n32356 & n70661);
  assign n70663 = (n56502 & n56875) | (n56502 & n70662) | (n56875 & n70662);
  assign n70664 = (n56501 & n56875) | (n56501 & n70662) | (n56875 & n70662);
  assign n70665 = (n70222 & n70663) | (n70222 & n70664) | (n70663 & n70664);
  assign n56637 = (n56252 & n70503) | (n56252 & n56636) | (n70503 & n56636);
  assign n56880 = n32333 | n32335;
  assign n70666 = n31856 | n32333;
  assign n70667 = (n32333 & n32335) | (n32333 & n70666) | (n32335 & n70666);
  assign n70668 = (n56492 & n56880) | (n56492 & n70667) | (n56880 & n70667);
  assign n70669 = (n56491 & n56880) | (n56491 & n70667) | (n56880 & n70667);
  assign n70670 = (n56149 & n70668) | (n56149 & n70669) | (n70668 & n70669);
  assign n56642 = (n56242 & n70505) | (n56242 & n56641) | (n70505 & n56641);
  assign n56885 = n32312 | n32314;
  assign n70671 = n31835 | n32312;
  assign n70672 = (n32312 & n32314) | (n32312 & n70671) | (n32314 & n70671);
  assign n70673 = (n56482 & n56885) | (n56482 & n70672) | (n56885 & n70672);
  assign n70674 = (n56481 & n56885) | (n56481 & n70672) | (n56885 & n70672);
  assign n70675 = (n56154 & n70673) | (n56154 & n70674) | (n70673 & n70674);
  assign n56401 = (n55934 & n70367) | (n55934 & n70369) | (n70367 & n70369);
  assign n70678 = n31800 | n32277;
  assign n70679 = (n32277 & n32279) | (n32277 & n70678) | (n32279 & n70678);
  assign n70680 = n32277 | n32279;
  assign n70681 = (n32277 & n56653) | (n32277 & n70680) | (n56653 & n70680);
  assign n70682 = (n56405 & n70679) | (n56405 & n70681) | (n70679 & n70681);
  assign n70683 = (n70371 & n70679) | (n70371 & n70681) | (n70679 & n70681);
  assign n70684 = (n70127 & n70682) | (n70127 & n70683) | (n70682 & n70683);
  assign n32704 = x174 & x176;
  assign n32705 = x173 & x177;
  assign n32706 = n32704 & n32705;
  assign n32707 = n32704 | n32705;
  assign n32708 = ~n32706 & n32707;
  assign n70685 = n32221 | n70525;
  assign n70688 = n32708 & n70685;
  assign n70686 = n32221 | n32223;
  assign n70689 = n32708 & n70686;
  assign n70690 = (n70383 & n70688) | (n70383 & n70689) | (n70688 & n70689);
  assign n70691 = n32221 & n32708;
  assign n70692 = (n32708 & n70532) | (n32708 & n70691) | (n70532 & n70691);
  assign n70693 = (n69747 & n70690) | (n69747 & n70692) | (n70690 & n70692);
  assign n70694 = (n69746 & n70690) | (n69746 & n70692) | (n70690 & n70692);
  assign n70695 = (n68195 & n70693) | (n68195 & n70694) | (n70693 & n70694);
  assign n70696 = n32708 | n70685;
  assign n70697 = n32708 | n70686;
  assign n70698 = (n70383 & n70696) | (n70383 & n70697) | (n70696 & n70697);
  assign n70699 = n32221 | n32708;
  assign n70700 = n70532 | n70699;
  assign n70701 = (n69747 & n70698) | (n69747 & n70700) | (n70698 & n70700);
  assign n70702 = (n69746 & n70698) | (n69746 & n70700) | (n70698 & n70700);
  assign n70703 = (n68195 & n70701) | (n68195 & n70702) | (n70701 & n70702);
  assign n32711 = ~n70695 & n70703;
  assign n32712 = x172 & x178;
  assign n32713 = n32711 & n32712;
  assign n32714 = n32711 | n32712;
  assign n32715 = ~n32713 & n32714;
  assign n70704 = n31751 | n32228;
  assign n70705 = (n32228 & n32230) | (n32228 & n70704) | (n32230 & n70704);
  assign n56921 = n32715 & n70705;
  assign n56910 = n32228 | n32230;
  assign n56922 = n32715 & n56910;
  assign n70706 = (n56921 & n56922) | (n56921 & n70398) | (n56922 & n70398);
  assign n70707 = (n56921 & n56922) | (n56921 & n70402) | (n56922 & n70402);
  assign n70708 = (n69887 & n70706) | (n69887 & n70707) | (n70706 & n70707);
  assign n56924 = n32715 | n70705;
  assign n56925 = n32715 | n56910;
  assign n70709 = (n56924 & n56925) | (n56924 & n70398) | (n56925 & n70398);
  assign n70710 = (n56924 & n56925) | (n56924 & n70402) | (n56925 & n70402);
  assign n70711 = (n69887 & n70709) | (n69887 & n70710) | (n70709 & n70710);
  assign n32718 = ~n70708 & n70711;
  assign n32719 = x171 & x179;
  assign n32720 = n32718 & n32719;
  assign n32721 = n32718 | n32719;
  assign n32722 = ~n32720 & n32721;
  assign n56907 = n32235 | n32237;
  assign n56927 = n32722 & n56907;
  assign n56928 = n32235 & n32722;
  assign n70712 = (n56927 & n56928) | (n56927 & n70524) | (n56928 & n70524);
  assign n70713 = (n56927 & n56928) | (n56927 & n70523) | (n56928 & n70523);
  assign n70714 = (n70013 & n70712) | (n70013 & n70713) | (n70712 & n70713);
  assign n56930 = n32722 | n56907;
  assign n56931 = n32235 | n32722;
  assign n70715 = (n56930 & n56931) | (n56930 & n70524) | (n56931 & n70524);
  assign n70716 = (n56930 & n56931) | (n56930 & n70523) | (n56931 & n70523);
  assign n70717 = (n70013 & n70715) | (n70013 & n70716) | (n70715 & n70716);
  assign n32725 = ~n70714 & n70717;
  assign n32726 = x170 & x180;
  assign n32727 = n32725 & n32726;
  assign n32728 = n32725 | n32726;
  assign n32729 = ~n32727 & n32728;
  assign n56905 = n32242 | n32244;
  assign n56933 = n32729 & n56905;
  assign n56934 = n32242 & n32729;
  assign n70718 = (n56933 & n56934) | (n56933 & n70520) | (n56934 & n70520);
  assign n70719 = (n56933 & n56934) | (n56933 & n70521) | (n56934 & n70521);
  assign n70720 = (n70133 & n70718) | (n70133 & n70719) | (n70718 & n70719);
  assign n56936 = n32729 | n56905;
  assign n56937 = n32242 | n32729;
  assign n70721 = (n56936 & n56937) | (n56936 & n70520) | (n56937 & n70520);
  assign n70722 = (n56936 & n56937) | (n56936 & n70521) | (n56937 & n70521);
  assign n70723 = (n70133 & n70721) | (n70133 & n70722) | (n70721 & n70722);
  assign n32732 = ~n70720 & n70723;
  assign n32733 = x169 & x181;
  assign n32734 = n32732 & n32733;
  assign n32735 = n32732 | n32733;
  assign n32736 = ~n32734 & n32735;
  assign n70724 = n32249 | n32251;
  assign n70725 = (n32249 & n56661) | (n32249 & n70724) | (n56661 & n70724);
  assign n56939 = n32736 & n70725;
  assign n70726 = n31772 | n32249;
  assign n70727 = (n32249 & n32251) | (n32249 & n70726) | (n32251 & n70726);
  assign n56940 = n32736 & n70727;
  assign n70728 = (n56939 & n56940) | (n56939 & n70376) | (n56940 & n70376);
  assign n70729 = (n56939 & n56940) | (n56939 & n70375) | (n56940 & n70375);
  assign n70730 = (n69736 & n70728) | (n69736 & n70729) | (n70728 & n70729);
  assign n56942 = n32736 | n70725;
  assign n56943 = n32736 | n70727;
  assign n70731 = (n56942 & n56943) | (n56942 & n70376) | (n56943 & n70376);
  assign n70732 = (n56942 & n56943) | (n56942 & n70375) | (n56943 & n70375);
  assign n70733 = (n69736 & n70731) | (n69736 & n70732) | (n70731 & n70732);
  assign n32739 = ~n70730 & n70733;
  assign n32740 = x168 & x182;
  assign n32741 = n32739 & n32740;
  assign n32742 = n32739 | n32740;
  assign n32743 = ~n32741 & n32742;
  assign n56945 = n32256 & n32743;
  assign n56946 = (n32743 & n70574) | (n32743 & n56945) | (n70574 & n56945);
  assign n56947 = n32256 | n32743;
  assign n56948 = n70574 | n56947;
  assign n32746 = ~n56946 & n56948;
  assign n32747 = x167 & x183;
  assign n32748 = n32746 & n32747;
  assign n32749 = n32746 | n32747;
  assign n32750 = ~n32748 & n32749;
  assign n70734 = n31786 | n32263;
  assign n70735 = (n32263 & n32265) | (n32263 & n70734) | (n32265 & n70734);
  assign n56949 = n32750 & n70735;
  assign n56900 = n32263 | n32265;
  assign n56950 = n32750 & n56900;
  assign n56951 = (n70430 & n56949) | (n70430 & n56950) | (n56949 & n56950);
  assign n56952 = n32750 | n70735;
  assign n56953 = n32750 | n56900;
  assign n56954 = (n70430 & n56952) | (n70430 & n56953) | (n56952 & n56953);
  assign n32753 = ~n56951 & n56954;
  assign n32754 = x166 & x184;
  assign n32755 = n32753 & n32754;
  assign n32756 = n32753 | n32754;
  assign n32757 = ~n32755 & n32756;
  assign n56897 = n32270 | n32272;
  assign n56955 = n32757 & n56897;
  assign n56956 = n32270 & n32757;
  assign n70736 = (n56955 & n56956) | (n56955 & n70516) | (n56956 & n70516);
  assign n70737 = (n56955 & n56956) | (n56955 & n70518) | (n56956 & n70518);
  assign n70738 = (n70235 & n70736) | (n70235 & n70737) | (n70736 & n70737);
  assign n56958 = n32757 | n56897;
  assign n56959 = n32270 | n32757;
  assign n70739 = (n56958 & n56959) | (n56958 & n70516) | (n56959 & n70516);
  assign n70740 = (n56958 & n56959) | (n56958 & n70518) | (n56959 & n70518);
  assign n70741 = (n70235 & n70739) | (n70235 & n70740) | (n70739 & n70740);
  assign n32760 = ~n70738 & n70741;
  assign n32761 = x165 & x185;
  assign n32762 = n32760 & n32761;
  assign n32763 = n32760 | n32761;
  assign n32764 = ~n32762 & n32763;
  assign n32765 = n70684 & n32764;
  assign n32766 = n70684 | n32764;
  assign n32767 = ~n32765 & n32766;
  assign n32768 = x164 & x186;
  assign n32769 = n32767 & n32768;
  assign n32770 = n32767 | n32768;
  assign n32771 = ~n32769 & n32770;
  assign n56892 = n32284 | n32286;
  assign n56961 = n32771 & n56892;
  assign n56962 = n32284 & n32771;
  assign n56963 = (n70514 & n56961) | (n70514 & n56962) | (n56961 & n56962);
  assign n56964 = n32771 | n56892;
  assign n56965 = n32284 | n32771;
  assign n56966 = (n70514 & n56964) | (n70514 & n56965) | (n56964 & n56965);
  assign n32774 = ~n56963 & n56966;
  assign n32775 = x163 & x187;
  assign n32776 = n32774 & n32775;
  assign n32777 = n32774 | n32775;
  assign n32778 = ~n32776 & n32777;
  assign n56890 = n32291 | n56704;
  assign n70742 = n32778 & n56890;
  assign n70676 = n31814 | n32291;
  assign n70677 = (n32291 & n32293) | (n32291 & n70676) | (n32293 & n70676);
  assign n70743 = n32778 & n70677;
  assign n70744 = (n56401 & n70742) | (n56401 & n70743) | (n70742 & n70743);
  assign n70745 = n32778 | n56890;
  assign n70746 = n32778 | n70677;
  assign n70747 = (n56401 & n70745) | (n56401 & n70746) | (n70745 & n70746);
  assign n32781 = ~n70744 & n70747;
  assign n32782 = x162 & x188;
  assign n32783 = n32781 & n32782;
  assign n32784 = n32781 | n32782;
  assign n32785 = ~n32783 & n32784;
  assign n56887 = n32298 | n32300;
  assign n56967 = n32785 & n56887;
  assign n56968 = n32298 & n32785;
  assign n70748 = (n56646 & n56967) | (n56646 & n56968) | (n56967 & n56968);
  assign n70749 = (n56967 & n56968) | (n56967 & n70507) | (n56968 & n70507);
  assign n70750 = (n56232 & n70748) | (n56232 & n70749) | (n70748 & n70749);
  assign n56970 = n32785 | n56887;
  assign n56971 = n32298 | n32785;
  assign n70751 = (n56646 & n56970) | (n56646 & n56971) | (n56970 & n56971);
  assign n70752 = (n56970 & n56971) | (n56970 & n70507) | (n56971 & n70507);
  assign n70753 = (n56232 & n70751) | (n56232 & n70752) | (n70751 & n70752);
  assign n32788 = ~n70750 & n70753;
  assign n32789 = x161 & x189;
  assign n32790 = n32788 & n32789;
  assign n32791 = n32788 | n32789;
  assign n32792 = ~n32790 & n32791;
  assign n56973 = n32305 & n32792;
  assign n56974 = (n32792 & n56712) | (n32792 & n56973) | (n56712 & n56973);
  assign n56975 = n32305 | n32792;
  assign n56976 = n56712 | n56975;
  assign n32795 = ~n56974 & n56976;
  assign n32796 = x160 & x190;
  assign n32797 = n32795 & n32796;
  assign n32798 = n32795 | n32796;
  assign n32799 = ~n32797 & n32798;
  assign n32800 = n70675 & n32799;
  assign n32801 = n70675 | n32799;
  assign n32802 = ~n32800 & n32801;
  assign n32803 = x159 & x191;
  assign n32804 = n32802 & n32803;
  assign n32805 = n32802 | n32803;
  assign n32806 = ~n32804 & n32805;
  assign n56882 = n32319 | n32321;
  assign n56977 = n32806 & n56882;
  assign n56978 = n32319 & n32806;
  assign n56979 = (n56642 & n56977) | (n56642 & n56978) | (n56977 & n56978);
  assign n56980 = n32806 | n56882;
  assign n56981 = n32319 | n32806;
  assign n56982 = (n56642 & n56980) | (n56642 & n56981) | (n56980 & n56981);
  assign n32809 = ~n56979 & n56982;
  assign n32810 = x158 & x192;
  assign n32811 = n32809 & n32810;
  assign n32812 = n32809 | n32810;
  assign n32813 = ~n32811 & n32812;
  assign n56983 = n32326 & n32813;
  assign n56984 = (n32813 & n56722) | (n32813 & n56983) | (n56722 & n56983);
  assign n56985 = n32326 | n32813;
  assign n56986 = n56722 | n56985;
  assign n32816 = ~n56984 & n56986;
  assign n32817 = x157 & x193;
  assign n32818 = n32816 & n32817;
  assign n32819 = n32816 | n32817;
  assign n32820 = ~n32818 & n32819;
  assign n32821 = n70670 & n32820;
  assign n32822 = n70670 | n32820;
  assign n32823 = ~n32821 & n32822;
  assign n32824 = x156 & x194;
  assign n32825 = n32823 & n32824;
  assign n32826 = n32823 | n32824;
  assign n32827 = ~n32825 & n32826;
  assign n56877 = n32340 | n32342;
  assign n56987 = n32827 & n56877;
  assign n56988 = n32340 & n32827;
  assign n56989 = (n56637 & n56987) | (n56637 & n56988) | (n56987 & n56988);
  assign n56990 = n32827 | n56877;
  assign n56991 = n32340 | n32827;
  assign n56992 = (n56637 & n56990) | (n56637 & n56991) | (n56990 & n56991);
  assign n32830 = ~n56989 & n56992;
  assign n32831 = x155 & x195;
  assign n32832 = n32830 & n32831;
  assign n32833 = n32830 | n32831;
  assign n32834 = ~n32832 & n32833;
  assign n56993 = n32347 & n32834;
  assign n56994 = (n32834 & n56732) | (n32834 & n56993) | (n56732 & n56993);
  assign n56995 = n32347 | n32834;
  assign n56996 = n56732 | n56995;
  assign n32837 = ~n56994 & n56996;
  assign n32838 = x154 & x196;
  assign n32839 = n32837 & n32838;
  assign n32840 = n32837 | n32838;
  assign n32841 = ~n32839 & n32840;
  assign n32842 = n70665 & n32841;
  assign n32843 = n70665 | n32841;
  assign n32844 = ~n32842 & n32843;
  assign n32845 = x153 & x197;
  assign n32846 = n32844 & n32845;
  assign n32847 = n32844 | n32845;
  assign n32848 = ~n32846 & n32847;
  assign n56872 = n32361 | n32363;
  assign n56997 = n32848 & n56872;
  assign n56998 = n32361 & n32848;
  assign n56999 = (n70501 & n56997) | (n70501 & n56998) | (n56997 & n56998);
  assign n57000 = n32848 | n56872;
  assign n57001 = n32361 | n32848;
  assign n57002 = (n70501 & n57000) | (n70501 & n57001) | (n57000 & n57001);
  assign n32851 = ~n56999 & n57002;
  assign n32852 = x152 & x198;
  assign n32853 = n32851 & n32852;
  assign n32854 = n32851 | n32852;
  assign n32855 = ~n32853 & n32854;
  assign n57003 = n32368 & n32855;
  assign n70754 = (n32855 & n56741) | (n32855 & n57003) | (n56741 & n57003);
  assign n70755 = (n32855 & n56740) | (n32855 & n57003) | (n56740 & n57003);
  assign n70756 = (n70350 & n70754) | (n70350 & n70755) | (n70754 & n70755);
  assign n57005 = n32368 | n32855;
  assign n70757 = n56741 | n57005;
  assign n70758 = n56740 | n57005;
  assign n70759 = (n70350 & n70757) | (n70350 & n70758) | (n70757 & n70758);
  assign n32858 = ~n70756 & n70759;
  assign n32859 = x151 & x199;
  assign n32860 = n32858 & n32859;
  assign n32861 = n32858 | n32859;
  assign n32862 = ~n32860 & n32861;
  assign n32863 = n70660 & n32862;
  assign n32864 = n70660 | n32862;
  assign n32865 = ~n32863 & n32864;
  assign n32866 = x150 & x200;
  assign n32867 = n32865 & n32866;
  assign n32868 = n32865 | n32866;
  assign n32869 = ~n32867 & n32868;
  assign n56867 = n32382 | n32384;
  assign n57007 = n32869 & n56867;
  assign n57008 = n32382 & n32869;
  assign n57009 = (n70496 & n57007) | (n70496 & n57008) | (n57007 & n57008);
  assign n57010 = n32869 | n56867;
  assign n57011 = n32382 | n32869;
  assign n57012 = (n70496 & n57010) | (n70496 & n57011) | (n57010 & n57011);
  assign n32872 = ~n57009 & n57012;
  assign n32873 = x149 & x201;
  assign n32874 = n32872 & n32873;
  assign n32875 = n32872 | n32873;
  assign n32876 = ~n32874 & n32875;
  assign n57013 = n32389 & n32876;
  assign n70760 = (n32876 & n56751) | (n32876 & n57013) | (n56751 & n57013);
  assign n70761 = (n32876 & n56750) | (n32876 & n57013) | (n56750 & n57013);
  assign n70762 = (n56378 & n70760) | (n56378 & n70761) | (n70760 & n70761);
  assign n57015 = n32389 | n32876;
  assign n70763 = n56751 | n57015;
  assign n70764 = n56750 | n57015;
  assign n70765 = (n56378 & n70763) | (n56378 & n70764) | (n70763 & n70764);
  assign n32879 = ~n70762 & n70765;
  assign n32880 = x148 & x202;
  assign n32881 = n32879 & n32880;
  assign n32882 = n32879 | n32880;
  assign n32883 = ~n32881 & n32882;
  assign n56865 = n32396 | n32398;
  assign n70766 = n32883 & n56865;
  assign n70654 = n31919 | n32396;
  assign n70655 = (n32396 & n32398) | (n32396 & n70654) | (n32398 & n70654);
  assign n70767 = n32883 & n70655;
  assign n70768 = (n70472 & n70766) | (n70472 & n70767) | (n70766 & n70767);
  assign n70769 = n32883 | n56865;
  assign n70770 = n32883 | n70655;
  assign n70771 = (n70472 & n70769) | (n70472 & n70770) | (n70769 & n70770);
  assign n32886 = ~n70768 & n70771;
  assign n32887 = x147 & x203;
  assign n32888 = n32886 & n32887;
  assign n32889 = n32886 | n32887;
  assign n32890 = ~n32888 & n32889;
  assign n57017 = n32403 & n32890;
  assign n70772 = (n32890 & n56760) | (n32890 & n57017) | (n56760 & n57017);
  assign n70773 = (n32405 & n32890) | (n32405 & n57017) | (n32890 & n57017);
  assign n70774 = (n56526 & n70772) | (n56526 & n70773) | (n70772 & n70773);
  assign n57019 = n32403 | n32890;
  assign n70775 = n56760 | n57019;
  assign n70776 = n32405 | n57019;
  assign n70777 = (n56526 & n70775) | (n56526 & n70776) | (n70775 & n70776);
  assign n32893 = ~n70774 & n70777;
  assign n32894 = x146 & x204;
  assign n32895 = n32893 & n32894;
  assign n32896 = n32893 | n32894;
  assign n32897 = ~n32895 & n32896;
  assign n57021 = n32410 & n32897;
  assign n57022 = (n32897 & n56765) | (n32897 & n57021) | (n56765 & n57021);
  assign n57023 = n32410 | n32897;
  assign n57024 = n56765 | n57023;
  assign n32900 = ~n57022 & n57024;
  assign n32901 = x145 & x205;
  assign n32902 = n32900 & n32901;
  assign n32903 = n32900 | n32901;
  assign n32904 = ~n32902 & n32903;
  assign n57025 = n32417 & n32904;
  assign n57026 = (n32904 & n56769) | (n32904 & n57025) | (n56769 & n57025);
  assign n57027 = n32417 | n32904;
  assign n57028 = n56769 | n57027;
  assign n32907 = ~n57026 & n57028;
  assign n32908 = x144 & x206;
  assign n32909 = n32907 & n32908;
  assign n32910 = n32907 | n32908;
  assign n32911 = ~n32909 & n32910;
  assign n57029 = n32424 & n32911;
  assign n57030 = (n32911 & n56773) | (n32911 & n57029) | (n56773 & n57029);
  assign n57031 = n32424 | n32911;
  assign n57032 = n56773 | n57031;
  assign n32914 = ~n57030 & n57032;
  assign n32915 = x143 & x207;
  assign n32916 = n32914 & n32915;
  assign n32917 = n32914 | n32915;
  assign n32918 = ~n32916 & n32917;
  assign n57033 = n32431 & n32918;
  assign n57034 = (n32918 & n56777) | (n32918 & n57033) | (n56777 & n57033);
  assign n57035 = n32431 | n32918;
  assign n57036 = n56777 | n57035;
  assign n32921 = ~n57034 & n57036;
  assign n32922 = x142 & x208;
  assign n32923 = n32921 & n32922;
  assign n32924 = n32921 | n32922;
  assign n32925 = ~n32923 & n32924;
  assign n57037 = n32438 & n32925;
  assign n57038 = (n32925 & n56781) | (n32925 & n57037) | (n56781 & n57037);
  assign n57039 = n32438 | n32925;
  assign n57040 = n56781 | n57039;
  assign n32928 = ~n57038 & n57040;
  assign n32929 = x141 & x209;
  assign n32930 = n32928 & n32929;
  assign n32931 = n32928 | n32929;
  assign n32932 = ~n32930 & n32931;
  assign n57041 = n32445 & n32932;
  assign n57042 = (n32932 & n56785) | (n32932 & n57041) | (n56785 & n57041);
  assign n57043 = n32445 | n32932;
  assign n57044 = n56785 | n57043;
  assign n32935 = ~n57042 & n57044;
  assign n32936 = x140 & x210;
  assign n32937 = n32935 & n32936;
  assign n32938 = n32935 | n32936;
  assign n32939 = ~n32937 & n32938;
  assign n57045 = n32452 & n32939;
  assign n57046 = (n32939 & n56789) | (n32939 & n57045) | (n56789 & n57045);
  assign n57047 = n32452 | n32939;
  assign n57048 = n56789 | n57047;
  assign n32942 = ~n57046 & n57048;
  assign n32943 = x139 & x211;
  assign n32944 = n32942 & n32943;
  assign n32945 = n32942 | n32943;
  assign n32946 = ~n32944 & n32945;
  assign n57049 = n32459 & n32946;
  assign n57050 = (n32946 & n56793) | (n32946 & n57049) | (n56793 & n57049);
  assign n57051 = n32459 | n32946;
  assign n57052 = n56793 | n57051;
  assign n32949 = ~n57050 & n57052;
  assign n32950 = x138 & x212;
  assign n32951 = n32949 & n32950;
  assign n32952 = n32949 | n32950;
  assign n32953 = ~n32951 & n32952;
  assign n57053 = n32466 & n32953;
  assign n57054 = (n32953 & n56797) | (n32953 & n57053) | (n56797 & n57053);
  assign n57055 = n32466 | n32953;
  assign n57056 = n56797 | n57055;
  assign n32956 = ~n57054 & n57056;
  assign n32957 = x137 & x213;
  assign n32958 = n32956 & n32957;
  assign n32959 = n32956 | n32957;
  assign n32960 = ~n32958 & n32959;
  assign n57057 = n32473 & n32960;
  assign n57058 = (n32960 & n56801) | (n32960 & n57057) | (n56801 & n57057);
  assign n57059 = n32473 | n32960;
  assign n57060 = n56801 | n57059;
  assign n32963 = ~n57058 & n57060;
  assign n32964 = x136 & x214;
  assign n32965 = n32963 & n32964;
  assign n32966 = n32963 | n32964;
  assign n32967 = ~n32965 & n32966;
  assign n57061 = n32480 & n32967;
  assign n57062 = (n32967 & n56805) | (n32967 & n57061) | (n56805 & n57061);
  assign n57063 = n32480 | n32967;
  assign n57064 = n56805 | n57063;
  assign n32970 = ~n57062 & n57064;
  assign n32971 = x135 & x215;
  assign n32972 = n32970 & n32971;
  assign n32973 = n32970 | n32971;
  assign n32974 = ~n32972 & n32973;
  assign n57065 = n32487 & n32974;
  assign n57066 = (n32974 & n56809) | (n32974 & n57065) | (n56809 & n57065);
  assign n57067 = n32487 | n32974;
  assign n57068 = n56809 | n57067;
  assign n32977 = ~n57066 & n57068;
  assign n32978 = x134 & x216;
  assign n32979 = n32977 & n32978;
  assign n32980 = n32977 | n32978;
  assign n32981 = ~n32979 & n32980;
  assign n57069 = n32494 & n32981;
  assign n57070 = (n32981 & n56813) | (n32981 & n57069) | (n56813 & n57069);
  assign n57071 = n32494 | n32981;
  assign n57072 = n56813 | n57071;
  assign n32984 = ~n57070 & n57072;
  assign n32985 = x133 & x217;
  assign n32986 = n32984 & n32985;
  assign n32987 = n32984 | n32985;
  assign n32988 = ~n32986 & n32987;
  assign n57073 = n32501 & n32988;
  assign n57074 = (n32988 & n56817) | (n32988 & n57073) | (n56817 & n57073);
  assign n57075 = n32501 | n32988;
  assign n57076 = n56817 | n57075;
  assign n32991 = ~n57074 & n57076;
  assign n32992 = x132 & x218;
  assign n32993 = n32991 & n32992;
  assign n32994 = n32991 | n32992;
  assign n32995 = ~n32993 & n32994;
  assign n57077 = n32508 & n32995;
  assign n57078 = (n32995 & n56821) | (n32995 & n57077) | (n56821 & n57077);
  assign n57079 = n32508 | n32995;
  assign n57080 = n56821 | n57079;
  assign n32998 = ~n57078 & n57080;
  assign n32999 = x131 & x219;
  assign n33000 = n32998 & n32999;
  assign n33001 = n32998 | n32999;
  assign n33002 = ~n33000 & n33001;
  assign n57081 = n32515 & n33002;
  assign n57082 = (n33002 & n56825) | (n33002 & n57081) | (n56825 & n57081);
  assign n57083 = n32515 | n33002;
  assign n57084 = n56825 | n57083;
  assign n33005 = ~n57082 & n57084;
  assign n33006 = x130 & x220;
  assign n33007 = n33005 & n33006;
  assign n33008 = n33005 | n33006;
  assign n33009 = ~n33007 & n33008;
  assign n57085 = n32522 & n33009;
  assign n57086 = (n33009 & n56830) | (n33009 & n57085) | (n56830 & n57085);
  assign n57087 = n32522 | n33009;
  assign n57088 = n56830 | n57087;
  assign n33012 = ~n57086 & n57088;
  assign n33013 = x129 & x221;
  assign n33014 = n33012 & n33013;
  assign n33015 = n33012 | n33013;
  assign n33016 = ~n33014 & n33015;
  assign n56862 = n32529 | n32531;
  assign n57089 = n33016 & n56862;
  assign n57090 = n32529 & n33016;
  assign n57091 = (n56620 & n57089) | (n56620 & n57090) | (n57089 & n57090);
  assign n57092 = n33016 | n56862;
  assign n57093 = n32529 | n33016;
  assign n57094 = (n56620 & n57092) | (n56620 & n57093) | (n57092 & n57093);
  assign n33019 = ~n57091 & n57094;
  assign n33020 = x128 & x222;
  assign n33021 = n33019 & n33020;
  assign n33022 = n33019 | n33020;
  assign n33023 = ~n33021 & n33022;
  assign n56860 = n32536 | n32538;
  assign n70778 = n33023 & n56860;
  assign n70779 = n32536 & n33023;
  assign n70780 = (n56618 & n70778) | (n56618 & n70779) | (n70778 & n70779);
  assign n70781 = n33023 | n56860;
  assign n70782 = n32536 | n33023;
  assign n70783 = (n56618 & n70781) | (n56618 & n70782) | (n70781 & n70782);
  assign n33026 = ~n70780 & n70783;
  assign n33027 = x127 & x223;
  assign n33028 = n33026 & n33027;
  assign n33029 = n33026 | n33027;
  assign n33030 = ~n33028 & n33029;
  assign n56858 = n32543 | n32545;
  assign n70784 = n33030 & n56858;
  assign n70785 = n32543 & n33030;
  assign n70786 = (n56616 & n70784) | (n56616 & n70785) | (n70784 & n70785);
  assign n70787 = n33030 | n56858;
  assign n70788 = n32543 | n33030;
  assign n70789 = (n56616 & n70787) | (n56616 & n70788) | (n70787 & n70788);
  assign n33033 = ~n70786 & n70789;
  assign n33034 = x126 & x224;
  assign n33035 = n33033 & n33034;
  assign n33036 = n33033 | n33034;
  assign n33037 = ~n33035 & n33036;
  assign n33038 = n56857 & n33037;
  assign n33039 = n56857 | n33037;
  assign n33040 = ~n33038 & n33039;
  assign n33041 = x125 & x225;
  assign n33042 = n33040 & n33041;
  assign n33043 = n33040 | n33041;
  assign n33044 = ~n33042 & n33043;
  assign n33045 = n56855 & n33044;
  assign n33046 = n56855 | n33044;
  assign n33047 = ~n33045 & n33046;
  assign n33048 = x124 & x226;
  assign n33049 = n33047 & n33048;
  assign n33050 = n33047 | n33048;
  assign n33051 = ~n33049 & n33050;
  assign n33052 = n56853 & n33051;
  assign n33053 = n56853 | n33051;
  assign n33054 = ~n33052 & n33053;
  assign n33055 = x123 & x227;
  assign n33056 = n33054 & n33055;
  assign n33057 = n33054 | n33055;
  assign n33058 = ~n33056 & n33057;
  assign n33059 = n70653 & n33058;
  assign n33060 = n70653 | n33058;
  assign n33061 = ~n33059 & n33060;
  assign n33062 = x122 & x228;
  assign n33063 = n33061 & n33062;
  assign n33064 = n33061 | n33062;
  assign n33065 = ~n33063 & n33064;
  assign n33066 = n56851 & n33065;
  assign n33067 = n56851 | n33065;
  assign n33068 = ~n33066 & n33067;
  assign n33069 = x121 & x229;
  assign n33070 = n33068 & n33069;
  assign n33071 = n33068 | n33069;
  assign n33072 = ~n33070 & n33071;
  assign n33073 = n56849 & n33072;
  assign n33074 = n56849 | n33072;
  assign n33075 = ~n33073 & n33074;
  assign n33076 = x120 & x230;
  assign n33077 = n33075 & n33076;
  assign n33078 = n33075 | n33076;
  assign n33079 = ~n33077 & n33078;
  assign n33080 = n56847 & n33079;
  assign n33081 = n56847 | n33079;
  assign n33082 = ~n33080 & n33081;
  assign n33083 = x119 & x231;
  assign n33084 = n33082 & n33083;
  assign n33085 = n33082 | n33083;
  assign n33086 = ~n33084 & n33085;
  assign n33087 = n56845 & n33086;
  assign n33088 = n56845 | n33086;
  assign n33089 = ~n33087 & n33088;
  assign n33090 = x118 & x232;
  assign n33091 = n33089 & n33090;
  assign n33092 = n33089 | n33090;
  assign n33093 = ~n33091 & n33092;
  assign n33094 = n56843 & n33093;
  assign n33095 = n56843 | n33093;
  assign n33096 = ~n33094 & n33095;
  assign n33097 = x117 & x233;
  assign n33098 = n33096 & n33097;
  assign n33099 = n33096 | n33097;
  assign n33100 = ~n33098 & n33099;
  assign n33101 = n56841 & n33100;
  assign n33102 = n56841 | n33100;
  assign n33103 = ~n33101 & n33102;
  assign n33104 = x116 & x234;
  assign n33105 = n33103 & n33104;
  assign n33106 = n33103 | n33104;
  assign n33107 = ~n33105 & n33106;
  assign n33108 = n56839 & n33107;
  assign n33109 = n56839 | n33107;
  assign n33110 = ~n33108 & n33109;
  assign n33111 = x115 & x235;
  assign n33112 = n33110 & n33111;
  assign n33113 = n33110 | n33111;
  assign n33114 = ~n33112 & n33113;
  assign n33115 = n56837 & n33114;
  assign n33116 = n56837 | n33114;
  assign n33117 = ~n33115 & n33116;
  assign n33118 = x114 & x236;
  assign n33119 = n33117 & n33118;
  assign n33120 = n33117 | n33118;
  assign n33121 = ~n33119 & n33120;
  assign n33122 = n56835 & n33121;
  assign n33123 = n56835 | n33121;
  assign n33124 = ~n33122 & n33123;
  assign n33125 = x113 & x237;
  assign n33126 = n33124 & n33125;
  assign n33127 = n33124 | n33125;
  assign n33128 = ~n33126 & n33127;
  assign n33129 = n32641 & n33128;
  assign n33130 = n32641 | n33128;
  assign n33131 = ~n33129 & n33130;
  assign n33132 = x112 & x238;
  assign n33133 = n33131 & n33132;
  assign n33134 = n33131 | n33132;
  assign n33135 = ~n33133 & n33134;
  assign n57095 = n32641 | n33126;
  assign n57096 = (n33126 & n33128) | (n33126 & n57095) | (n33128 & n57095);
  assign n57097 = n33119 | n56835;
  assign n57098 = (n33119 & n33121) | (n33119 & n57097) | (n33121 & n57097);
  assign n57099 = n33112 | n56837;
  assign n57100 = (n33112 & n33114) | (n33112 & n57099) | (n33114 & n57099);
  assign n57101 = n33105 | n56839;
  assign n57102 = (n33105 & n33107) | (n33105 & n57101) | (n33107 & n57101);
  assign n57103 = n33098 | n56841;
  assign n57104 = (n33098 & n33100) | (n33098 & n57103) | (n33100 & n57103);
  assign n57105 = n33091 | n56843;
  assign n57106 = (n33091 & n33093) | (n33091 & n57105) | (n33093 & n57105);
  assign n57107 = n33084 | n56845;
  assign n57108 = (n33084 & n33086) | (n33084 & n57107) | (n33086 & n57107);
  assign n57109 = n33077 | n56847;
  assign n57110 = (n33077 & n33079) | (n33077 & n57109) | (n33079 & n57109);
  assign n57111 = n33070 | n56849;
  assign n57112 = (n33070 & n33072) | (n33070 & n57111) | (n33072 & n57111);
  assign n57113 = n33063 | n56851;
  assign n57114 = (n33063 & n33065) | (n33063 & n57113) | (n33065 & n57113);
  assign n57115 = n33056 | n33058;
  assign n57116 = (n70653 & n33056) | (n70653 & n57115) | (n33056 & n57115);
  assign n57117 = n33049 | n33051;
  assign n57118 = (n33049 & n56853) | (n33049 & n57117) | (n56853 & n57117);
  assign n57119 = n33042 | n33044;
  assign n57120 = (n33042 & n56855) | (n33042 & n57119) | (n56855 & n57119);
  assign n56859 = (n32543 & n56616) | (n32543 & n56858) | (n56616 & n56858);
  assign n56861 = (n32536 & n56618) | (n32536 & n56860) | (n56618 & n56860);
  assign n56866 = (n70472 & n70655) | (n70472 & n56865) | (n70655 & n56865);
  assign n57130 = n32874 | n32876;
  assign n70790 = n32389 | n32874;
  assign n70791 = (n32874 & n32876) | (n32874 & n70790) | (n32876 & n70790);
  assign n70792 = (n56751 & n57130) | (n56751 & n70791) | (n57130 & n70791);
  assign n70793 = (n56750 & n57130) | (n56750 & n70791) | (n57130 & n70791);
  assign n70794 = (n56378 & n70792) | (n56378 & n70793) | (n70792 & n70793);
  assign n57135 = n32853 | n32855;
  assign n70795 = n32368 | n32853;
  assign n70796 = (n32853 & n32855) | (n32853 & n70795) | (n32855 & n70795);
  assign n70797 = (n56741 & n57135) | (n56741 & n70796) | (n57135 & n70796);
  assign n70798 = (n56740 & n57135) | (n56740 & n70796) | (n57135 & n70796);
  assign n70799 = (n70350 & n70797) | (n70350 & n70798) | (n70797 & n70798);
  assign n56647 = (n56232 & n70507) | (n56232 & n56646) | (n70507 & n56646);
  assign n70810 = n32755 | n32757;
  assign n70811 = (n32755 & n56897) | (n32755 & n70810) | (n56897 & n70810);
  assign n70812 = n32270 | n32755;
  assign n70813 = (n32755 & n32757) | (n32755 & n70812) | (n32757 & n70812);
  assign n70814 = (n70516 & n70811) | (n70516 & n70813) | (n70811 & n70813);
  assign n70815 = (n70518 & n70811) | (n70518 & n70813) | (n70811 & n70813);
  assign n70816 = (n70235 & n70814) | (n70235 & n70815) | (n70814 & n70815);
  assign n70817 = n32734 | n32736;
  assign n70818 = (n32734 & n70727) | (n32734 & n70817) | (n70727 & n70817);
  assign n70819 = (n32734 & n70725) | (n32734 & n70817) | (n70725 & n70817);
  assign n70820 = (n70376 & n70818) | (n70376 & n70819) | (n70818 & n70819);
  assign n70821 = (n70375 & n70818) | (n70375 & n70819) | (n70818 & n70819);
  assign n70822 = (n69736 & n70820) | (n69736 & n70821) | (n70820 & n70821);
  assign n33197 = x175 & x176;
  assign n33198 = x174 & x177;
  assign n33199 = n33197 & n33198;
  assign n33200 = n33197 | n33198;
  assign n33201 = ~n33199 & n33200;
  assign n57183 = n32706 & n33201;
  assign n57184 = (n33201 & n70695) | (n33201 & n57183) | (n70695 & n57183);
  assign n57185 = n32706 | n33201;
  assign n57186 = n70695 | n57185;
  assign n33204 = ~n57184 & n57186;
  assign n33205 = x173 & x178;
  assign n33206 = n33204 & n33205;
  assign n33207 = n33204 | n33205;
  assign n33208 = ~n33206 & n33207;
  assign n70823 = n32713 | n32715;
  assign n70824 = (n32713 & n70705) | (n32713 & n70823) | (n70705 & n70823);
  assign n57187 = n33208 & n70824;
  assign n70825 = (n32713 & n56910) | (n32713 & n70823) | (n56910 & n70823);
  assign n57188 = n33208 & n70825;
  assign n70826 = (n57187 & n57188) | (n57187 & n70398) | (n57188 & n70398);
  assign n70827 = (n57187 & n57188) | (n57187 & n70402) | (n57188 & n70402);
  assign n70828 = (n69887 & n70826) | (n69887 & n70827) | (n70826 & n70827);
  assign n57190 = n33208 | n70824;
  assign n57191 = n33208 | n70825;
  assign n70829 = (n57190 & n57191) | (n57190 & n70398) | (n57191 & n70398);
  assign n70830 = (n57190 & n57191) | (n57190 & n70402) | (n57191 & n70402);
  assign n70831 = (n69887 & n70829) | (n69887 & n70830) | (n70829 & n70830);
  assign n33211 = ~n70828 & n70831;
  assign n33212 = x172 & x179;
  assign n33213 = n33211 & n33212;
  assign n33214 = n33211 | n33212;
  assign n33215 = ~n33213 & n33214;
  assign n70832 = n32720 | n32722;
  assign n70833 = (n32720 & n56907) | (n32720 & n70832) | (n56907 & n70832);
  assign n57193 = n33215 & n70833;
  assign n70834 = n32235 | n32720;
  assign n70835 = (n32720 & n32722) | (n32720 & n70834) | (n32722 & n70834);
  assign n57194 = n33215 & n70835;
  assign n70836 = (n57193 & n57194) | (n57193 & n70524) | (n57194 & n70524);
  assign n70837 = (n57193 & n57194) | (n57193 & n70523) | (n57194 & n70523);
  assign n70838 = (n70013 & n70836) | (n70013 & n70837) | (n70836 & n70837);
  assign n57196 = n33215 | n70833;
  assign n57197 = n33215 | n70835;
  assign n70839 = (n57196 & n57197) | (n57196 & n70524) | (n57197 & n70524);
  assign n70840 = (n57196 & n57197) | (n57196 & n70523) | (n57197 & n70523);
  assign n70841 = (n70013 & n70839) | (n70013 & n70840) | (n70839 & n70840);
  assign n33218 = ~n70838 & n70841;
  assign n33219 = x171 & x180;
  assign n33220 = n33218 & n33219;
  assign n33221 = n33218 | n33219;
  assign n33222 = ~n33220 & n33221;
  assign n70842 = n32727 | n32729;
  assign n70843 = (n32727 & n56905) | (n32727 & n70842) | (n56905 & n70842);
  assign n57199 = n33222 & n70843;
  assign n70844 = n32242 | n32727;
  assign n70845 = (n32727 & n32729) | (n32727 & n70844) | (n32729 & n70844);
  assign n57200 = n33222 & n70845;
  assign n70846 = (n57199 & n57200) | (n57199 & n70520) | (n57200 & n70520);
  assign n70847 = (n57199 & n57200) | (n57199 & n70521) | (n57200 & n70521);
  assign n70848 = (n70133 & n70846) | (n70133 & n70847) | (n70846 & n70847);
  assign n57202 = n33222 | n70843;
  assign n57203 = n33222 | n70845;
  assign n70849 = (n57202 & n57203) | (n57202 & n70520) | (n57203 & n70520);
  assign n70850 = (n57202 & n57203) | (n57202 & n70521) | (n57203 & n70521);
  assign n70851 = (n70133 & n70849) | (n70133 & n70850) | (n70849 & n70850);
  assign n33225 = ~n70848 & n70851;
  assign n33226 = x170 & x181;
  assign n33227 = n33225 & n33226;
  assign n33228 = n33225 | n33226;
  assign n33229 = ~n33227 & n33228;
  assign n33230 = n70822 & n33229;
  assign n33231 = n70822 | n33229;
  assign n33232 = ~n33230 & n33231;
  assign n33233 = x169 & x182;
  assign n33234 = n33232 & n33233;
  assign n33235 = n33232 | n33233;
  assign n33236 = ~n33234 & n33235;
  assign n70852 = n32256 | n32741;
  assign n70853 = (n32741 & n32743) | (n32741 & n70852) | (n32743 & n70852);
  assign n57205 = n33236 & n70853;
  assign n57169 = n32741 | n32743;
  assign n57206 = n33236 & n57169;
  assign n57207 = (n70574 & n57205) | (n70574 & n57206) | (n57205 & n57206);
  assign n57208 = n33236 | n70853;
  assign n57209 = n33236 | n57169;
  assign n57210 = (n70574 & n57208) | (n70574 & n57209) | (n57208 & n57209);
  assign n33239 = ~n57207 & n57210;
  assign n33240 = x168 & x183;
  assign n33241 = n33239 & n33240;
  assign n33242 = n33239 | n33240;
  assign n33243 = ~n33241 & n33242;
  assign n57166 = n32748 | n56950;
  assign n70854 = n33243 & n57166;
  assign n57165 = n32748 | n56949;
  assign n70855 = n33243 & n57165;
  assign n70856 = (n70430 & n70854) | (n70430 & n70855) | (n70854 & n70855);
  assign n70857 = n33243 | n57166;
  assign n70858 = n33243 | n57165;
  assign n70859 = (n70430 & n70857) | (n70430 & n70858) | (n70857 & n70858);
  assign n33246 = ~n70856 & n70859;
  assign n33247 = x167 & x184;
  assign n33248 = n33246 & n33247;
  assign n33249 = n33246 | n33247;
  assign n33250 = ~n33248 & n33249;
  assign n33251 = n70816 & n33250;
  assign n33252 = n70816 | n33250;
  assign n33253 = ~n33251 & n33252;
  assign n33254 = x166 & x185;
  assign n33255 = n33253 & n33254;
  assign n33256 = n33253 | n33254;
  assign n33257 = ~n33255 & n33256;
  assign n57160 = n32762 | n32764;
  assign n57211 = n33257 & n57160;
  assign n57212 = n32762 & n33257;
  assign n57213 = (n70684 & n57211) | (n70684 & n57212) | (n57211 & n57212);
  assign n57214 = n33257 | n57160;
  assign n57215 = n32762 | n33257;
  assign n57216 = (n70684 & n57214) | (n70684 & n57215) | (n57214 & n57215);
  assign n33260 = ~n57213 & n57216;
  assign n33261 = x165 & x186;
  assign n33262 = n33260 & n33261;
  assign n33263 = n33260 | n33261;
  assign n33264 = ~n33262 & n33263;
  assign n57158 = n32769 | n56961;
  assign n70860 = n33264 & n57158;
  assign n70808 = n32284 | n32769;
  assign n70809 = (n32769 & n32771) | (n32769 & n70808) | (n32771 & n70808);
  assign n70861 = n33264 & n70809;
  assign n70862 = (n70514 & n70860) | (n70514 & n70861) | (n70860 & n70861);
  assign n70863 = n33264 | n57158;
  assign n70864 = n33264 | n70809;
  assign n70865 = (n70514 & n70863) | (n70514 & n70864) | (n70863 & n70864);
  assign n33267 = ~n70862 & n70865;
  assign n33268 = x164 & x187;
  assign n33269 = n33267 & n33268;
  assign n33270 = n33267 | n33268;
  assign n33271 = ~n33269 & n33270;
  assign n57155 = n32776 | n32778;
  assign n57217 = n33271 & n57155;
  assign n57218 = n32776 & n33271;
  assign n70866 = (n56890 & n57217) | (n56890 & n57218) | (n57217 & n57218);
  assign n70867 = (n57217 & n57218) | (n57217 & n70677) | (n57218 & n70677);
  assign n70868 = (n56401 & n70866) | (n56401 & n70867) | (n70866 & n70867);
  assign n57220 = n33271 | n57155;
  assign n57221 = n32776 | n33271;
  assign n70869 = (n56890 & n57220) | (n56890 & n57221) | (n57220 & n57221);
  assign n70870 = (n57220 & n57221) | (n57220 & n70677) | (n57221 & n70677);
  assign n70871 = (n56401 & n70869) | (n56401 & n70870) | (n70869 & n70870);
  assign n33274 = ~n70868 & n70871;
  assign n33275 = x163 & x188;
  assign n33276 = n33274 & n33275;
  assign n33277 = n33274 | n33275;
  assign n33278 = ~n33276 & n33277;
  assign n57153 = n32783 | n56967;
  assign n70872 = n33278 & n57153;
  assign n70806 = n32298 | n32783;
  assign n70807 = (n32783 & n32785) | (n32783 & n70806) | (n32785 & n70806);
  assign n70873 = n33278 & n70807;
  assign n70874 = (n56647 & n70872) | (n56647 & n70873) | (n70872 & n70873);
  assign n70875 = n33278 | n57153;
  assign n70876 = n33278 | n70807;
  assign n70877 = (n56647 & n70875) | (n56647 & n70876) | (n70875 & n70876);
  assign n33281 = ~n70874 & n70877;
  assign n33282 = x162 & x189;
  assign n33283 = n33281 & n33282;
  assign n33284 = n33281 | n33282;
  assign n33285 = ~n33283 & n33284;
  assign n57150 = n32790 | n32792;
  assign n70878 = n33285 & n57150;
  assign n70804 = n32305 | n32790;
  assign n70805 = (n32790 & n32792) | (n32790 & n70804) | (n32792 & n70804);
  assign n70879 = n33285 & n70805;
  assign n70880 = (n56712 & n70878) | (n56712 & n70879) | (n70878 & n70879);
  assign n70881 = n33285 | n57150;
  assign n70882 = n33285 | n70805;
  assign n70883 = (n56712 & n70881) | (n56712 & n70882) | (n70881 & n70882);
  assign n33288 = ~n70880 & n70883;
  assign n33289 = x161 & x190;
  assign n33290 = n33288 & n33289;
  assign n33291 = n33288 | n33289;
  assign n33292 = ~n33290 & n33291;
  assign n57147 = n32797 | n32799;
  assign n57223 = n33292 & n57147;
  assign n57224 = n32797 & n33292;
  assign n57225 = (n70675 & n57223) | (n70675 & n57224) | (n57223 & n57224);
  assign n57226 = n33292 | n57147;
  assign n57227 = n32797 | n33292;
  assign n57228 = (n70675 & n57226) | (n70675 & n57227) | (n57226 & n57227);
  assign n33295 = ~n57225 & n57228;
  assign n33296 = x160 & x191;
  assign n33297 = n33295 & n33296;
  assign n33298 = n33295 | n33296;
  assign n33299 = ~n33297 & n33298;
  assign n57229 = n32804 & n33299;
  assign n70884 = (n33299 & n56978) | (n33299 & n57229) | (n56978 & n57229);
  assign n70885 = (n33299 & n56977) | (n33299 & n57229) | (n56977 & n57229);
  assign n70886 = (n56642 & n70884) | (n56642 & n70885) | (n70884 & n70885);
  assign n57231 = n32804 | n33299;
  assign n70887 = n56978 | n57231;
  assign n70888 = n56977 | n57231;
  assign n70889 = (n56642 & n70887) | (n56642 & n70888) | (n70887 & n70888);
  assign n33302 = ~n70886 & n70889;
  assign n33303 = x159 & x192;
  assign n33304 = n33302 & n33303;
  assign n33305 = n33302 | n33303;
  assign n33306 = ~n33304 & n33305;
  assign n57145 = n32811 | n32813;
  assign n70890 = n33306 & n57145;
  assign n70802 = n32326 | n32811;
  assign n70803 = (n32811 & n32813) | (n32811 & n70802) | (n32813 & n70802);
  assign n70891 = n33306 & n70803;
  assign n70892 = (n56722 & n70890) | (n56722 & n70891) | (n70890 & n70891);
  assign n70893 = n33306 | n57145;
  assign n70894 = n33306 | n70803;
  assign n70895 = (n56722 & n70893) | (n56722 & n70894) | (n70893 & n70894);
  assign n33309 = ~n70892 & n70895;
  assign n33310 = x158 & x193;
  assign n33311 = n33309 & n33310;
  assign n33312 = n33309 | n33310;
  assign n33313 = ~n33311 & n33312;
  assign n57142 = n32818 | n32820;
  assign n57233 = n33313 & n57142;
  assign n57234 = n32818 & n33313;
  assign n57235 = (n70670 & n57233) | (n70670 & n57234) | (n57233 & n57234);
  assign n57236 = n33313 | n57142;
  assign n57237 = n32818 | n33313;
  assign n57238 = (n70670 & n57236) | (n70670 & n57237) | (n57236 & n57237);
  assign n33316 = ~n57235 & n57238;
  assign n33317 = x157 & x194;
  assign n33318 = n33316 & n33317;
  assign n33319 = n33316 | n33317;
  assign n33320 = ~n33318 & n33319;
  assign n57239 = n32825 & n33320;
  assign n70896 = (n33320 & n56988) | (n33320 & n57239) | (n56988 & n57239);
  assign n70897 = (n33320 & n56987) | (n33320 & n57239) | (n56987 & n57239);
  assign n70898 = (n56637 & n70896) | (n56637 & n70897) | (n70896 & n70897);
  assign n57241 = n32825 | n33320;
  assign n70899 = n56988 | n57241;
  assign n70900 = n56987 | n57241;
  assign n70901 = (n56637 & n70899) | (n56637 & n70900) | (n70899 & n70900);
  assign n33323 = ~n70898 & n70901;
  assign n33324 = x156 & x195;
  assign n33325 = n33323 & n33324;
  assign n33326 = n33323 | n33324;
  assign n33327 = ~n33325 & n33326;
  assign n57140 = n32832 | n32834;
  assign n70902 = n33327 & n57140;
  assign n70800 = n32347 | n32832;
  assign n70801 = (n32832 & n32834) | (n32832 & n70800) | (n32834 & n70800);
  assign n70903 = n33327 & n70801;
  assign n70904 = (n56732 & n70902) | (n56732 & n70903) | (n70902 & n70903);
  assign n70905 = n33327 | n57140;
  assign n70906 = n33327 | n70801;
  assign n70907 = (n56732 & n70905) | (n56732 & n70906) | (n70905 & n70906);
  assign n33330 = ~n70904 & n70907;
  assign n33331 = x155 & x196;
  assign n33332 = n33330 & n33331;
  assign n33333 = n33330 | n33331;
  assign n33334 = ~n33332 & n33333;
  assign n57137 = n32839 | n32841;
  assign n57243 = n33334 & n57137;
  assign n57244 = n32839 & n33334;
  assign n57245 = (n70665 & n57243) | (n70665 & n57244) | (n57243 & n57244);
  assign n57246 = n33334 | n57137;
  assign n57247 = n32839 | n33334;
  assign n57248 = (n70665 & n57246) | (n70665 & n57247) | (n57246 & n57247);
  assign n33337 = ~n57245 & n57248;
  assign n33338 = x154 & x197;
  assign n33339 = n33337 & n33338;
  assign n33340 = n33337 | n33338;
  assign n33341 = ~n33339 & n33340;
  assign n57249 = n32846 & n33341;
  assign n70908 = (n33341 & n56998) | (n33341 & n57249) | (n56998 & n57249);
  assign n70909 = (n33341 & n56997) | (n33341 & n57249) | (n56997 & n57249);
  assign n70910 = (n70501 & n70908) | (n70501 & n70909) | (n70908 & n70909);
  assign n57251 = n32846 | n33341;
  assign n70911 = n56998 | n57251;
  assign n70912 = n56997 | n57251;
  assign n70913 = (n70501 & n70911) | (n70501 & n70912) | (n70911 & n70912);
  assign n33344 = ~n70910 & n70913;
  assign n33345 = x153 & x198;
  assign n33346 = n33344 & n33345;
  assign n33347 = n33344 | n33345;
  assign n33348 = ~n33346 & n33347;
  assign n33349 = n70799 & n33348;
  assign n33350 = n70799 | n33348;
  assign n33351 = ~n33349 & n33350;
  assign n33352 = x152 & x199;
  assign n33353 = n33351 & n33352;
  assign n33354 = n33351 | n33352;
  assign n33355 = ~n33353 & n33354;
  assign n57132 = n32860 | n32862;
  assign n57253 = n33355 & n57132;
  assign n57254 = n32860 & n33355;
  assign n57255 = (n70660 & n57253) | (n70660 & n57254) | (n57253 & n57254);
  assign n57256 = n33355 | n57132;
  assign n57257 = n32860 | n33355;
  assign n57258 = (n70660 & n57256) | (n70660 & n57257) | (n57256 & n57257);
  assign n33358 = ~n57255 & n57258;
  assign n33359 = x151 & x200;
  assign n33360 = n33358 & n33359;
  assign n33361 = n33358 | n33359;
  assign n33362 = ~n33360 & n33361;
  assign n57259 = n32867 & n33362;
  assign n70914 = (n33362 & n57008) | (n33362 & n57259) | (n57008 & n57259);
  assign n70915 = (n33362 & n57007) | (n33362 & n57259) | (n57007 & n57259);
  assign n70916 = (n70496 & n70914) | (n70496 & n70915) | (n70914 & n70915);
  assign n57261 = n32867 | n33362;
  assign n70917 = n57008 | n57261;
  assign n70918 = n57007 | n57261;
  assign n70919 = (n70496 & n70917) | (n70496 & n70918) | (n70917 & n70918);
  assign n33365 = ~n70916 & n70919;
  assign n33366 = x150 & x201;
  assign n33367 = n33365 & n33366;
  assign n33368 = n33365 | n33366;
  assign n33369 = ~n33367 & n33368;
  assign n33370 = n70794 & n33369;
  assign n33371 = n70794 | n33369;
  assign n33372 = ~n33370 & n33371;
  assign n33373 = x149 & x202;
  assign n33374 = n33372 & n33373;
  assign n33375 = n33372 | n33373;
  assign n33376 = ~n33374 & n33375;
  assign n57127 = n32881 | n32883;
  assign n57263 = n33376 & n57127;
  assign n57264 = n32881 & n33376;
  assign n57265 = (n56866 & n57263) | (n56866 & n57264) | (n57263 & n57264);
  assign n57266 = n33376 | n57127;
  assign n57267 = n32881 | n33376;
  assign n57268 = (n56866 & n57266) | (n56866 & n57267) | (n57266 & n57267);
  assign n33379 = ~n57265 & n57268;
  assign n33380 = x148 & x203;
  assign n33381 = n33379 & n33380;
  assign n33382 = n33379 | n33380;
  assign n33383 = ~n33381 & n33382;
  assign n57269 = n32888 & n33383;
  assign n57270 = (n33383 & n70774) | (n33383 & n57269) | (n70774 & n57269);
  assign n57271 = n32888 | n33383;
  assign n57272 = n70774 | n57271;
  assign n33386 = ~n57270 & n57272;
  assign n33387 = x147 & x204;
  assign n33388 = n33386 & n33387;
  assign n33389 = n33386 | n33387;
  assign n33390 = ~n33388 & n33389;
  assign n57273 = n32895 & n33390;
  assign n57274 = (n33390 & n57022) | (n33390 & n57273) | (n57022 & n57273);
  assign n57275 = n32895 | n33390;
  assign n57276 = n57022 | n57275;
  assign n33393 = ~n57274 & n57276;
  assign n33394 = x146 & x205;
  assign n33395 = n33393 & n33394;
  assign n33396 = n33393 | n33394;
  assign n33397 = ~n33395 & n33396;
  assign n57277 = n32902 & n33397;
  assign n57278 = (n33397 & n57026) | (n33397 & n57277) | (n57026 & n57277);
  assign n57279 = n32902 | n33397;
  assign n57280 = n57026 | n57279;
  assign n33400 = ~n57278 & n57280;
  assign n33401 = x145 & x206;
  assign n33402 = n33400 & n33401;
  assign n33403 = n33400 | n33401;
  assign n33404 = ~n33402 & n33403;
  assign n57281 = n32909 & n33404;
  assign n57282 = (n33404 & n57030) | (n33404 & n57281) | (n57030 & n57281);
  assign n57283 = n32909 | n33404;
  assign n57284 = n57030 | n57283;
  assign n33407 = ~n57282 & n57284;
  assign n33408 = x144 & x207;
  assign n33409 = n33407 & n33408;
  assign n33410 = n33407 | n33408;
  assign n33411 = ~n33409 & n33410;
  assign n57285 = n32916 & n33411;
  assign n57286 = (n33411 & n57034) | (n33411 & n57285) | (n57034 & n57285);
  assign n57287 = n32916 | n33411;
  assign n57288 = n57034 | n57287;
  assign n33414 = ~n57286 & n57288;
  assign n33415 = x143 & x208;
  assign n33416 = n33414 & n33415;
  assign n33417 = n33414 | n33415;
  assign n33418 = ~n33416 & n33417;
  assign n57289 = n32923 & n33418;
  assign n57290 = (n33418 & n57038) | (n33418 & n57289) | (n57038 & n57289);
  assign n57291 = n32923 | n33418;
  assign n57292 = n57038 | n57291;
  assign n33421 = ~n57290 & n57292;
  assign n33422 = x142 & x209;
  assign n33423 = n33421 & n33422;
  assign n33424 = n33421 | n33422;
  assign n33425 = ~n33423 & n33424;
  assign n57293 = n32930 & n33425;
  assign n57294 = (n33425 & n57042) | (n33425 & n57293) | (n57042 & n57293);
  assign n57295 = n32930 | n33425;
  assign n57296 = n57042 | n57295;
  assign n33428 = ~n57294 & n57296;
  assign n33429 = x141 & x210;
  assign n33430 = n33428 & n33429;
  assign n33431 = n33428 | n33429;
  assign n33432 = ~n33430 & n33431;
  assign n57297 = n32937 & n33432;
  assign n57298 = (n33432 & n57046) | (n33432 & n57297) | (n57046 & n57297);
  assign n57299 = n32937 | n33432;
  assign n57300 = n57046 | n57299;
  assign n33435 = ~n57298 & n57300;
  assign n33436 = x140 & x211;
  assign n33437 = n33435 & n33436;
  assign n33438 = n33435 | n33436;
  assign n33439 = ~n33437 & n33438;
  assign n57301 = n32944 & n33439;
  assign n57302 = (n33439 & n57050) | (n33439 & n57301) | (n57050 & n57301);
  assign n57303 = n32944 | n33439;
  assign n57304 = n57050 | n57303;
  assign n33442 = ~n57302 & n57304;
  assign n33443 = x139 & x212;
  assign n33444 = n33442 & n33443;
  assign n33445 = n33442 | n33443;
  assign n33446 = ~n33444 & n33445;
  assign n57305 = n32951 & n33446;
  assign n57306 = (n33446 & n57054) | (n33446 & n57305) | (n57054 & n57305);
  assign n57307 = n32951 | n33446;
  assign n57308 = n57054 | n57307;
  assign n33449 = ~n57306 & n57308;
  assign n33450 = x138 & x213;
  assign n33451 = n33449 & n33450;
  assign n33452 = n33449 | n33450;
  assign n33453 = ~n33451 & n33452;
  assign n57309 = n32958 & n33453;
  assign n57310 = (n33453 & n57058) | (n33453 & n57309) | (n57058 & n57309);
  assign n57311 = n32958 | n33453;
  assign n57312 = n57058 | n57311;
  assign n33456 = ~n57310 & n57312;
  assign n33457 = x137 & x214;
  assign n33458 = n33456 & n33457;
  assign n33459 = n33456 | n33457;
  assign n33460 = ~n33458 & n33459;
  assign n57313 = n32965 & n33460;
  assign n57314 = (n33460 & n57062) | (n33460 & n57313) | (n57062 & n57313);
  assign n57315 = n32965 | n33460;
  assign n57316 = n57062 | n57315;
  assign n33463 = ~n57314 & n57316;
  assign n33464 = x136 & x215;
  assign n33465 = n33463 & n33464;
  assign n33466 = n33463 | n33464;
  assign n33467 = ~n33465 & n33466;
  assign n57317 = n32972 & n33467;
  assign n57318 = (n33467 & n57066) | (n33467 & n57317) | (n57066 & n57317);
  assign n57319 = n32972 | n33467;
  assign n57320 = n57066 | n57319;
  assign n33470 = ~n57318 & n57320;
  assign n33471 = x135 & x216;
  assign n33472 = n33470 & n33471;
  assign n33473 = n33470 | n33471;
  assign n33474 = ~n33472 & n33473;
  assign n57321 = n32979 & n33474;
  assign n57322 = (n33474 & n57070) | (n33474 & n57321) | (n57070 & n57321);
  assign n57323 = n32979 | n33474;
  assign n57324 = n57070 | n57323;
  assign n33477 = ~n57322 & n57324;
  assign n33478 = x134 & x217;
  assign n33479 = n33477 & n33478;
  assign n33480 = n33477 | n33478;
  assign n33481 = ~n33479 & n33480;
  assign n57325 = n32986 & n33481;
  assign n57326 = (n33481 & n57074) | (n33481 & n57325) | (n57074 & n57325);
  assign n57327 = n32986 | n33481;
  assign n57328 = n57074 | n57327;
  assign n33484 = ~n57326 & n57328;
  assign n33485 = x133 & x218;
  assign n33486 = n33484 & n33485;
  assign n33487 = n33484 | n33485;
  assign n33488 = ~n33486 & n33487;
  assign n57329 = n32993 & n33488;
  assign n57330 = (n33488 & n57078) | (n33488 & n57329) | (n57078 & n57329);
  assign n57331 = n32993 | n33488;
  assign n57332 = n57078 | n57331;
  assign n33491 = ~n57330 & n57332;
  assign n33492 = x132 & x219;
  assign n33493 = n33491 & n33492;
  assign n33494 = n33491 | n33492;
  assign n33495 = ~n33493 & n33494;
  assign n57333 = n33000 & n33495;
  assign n57334 = (n33495 & n57082) | (n33495 & n57333) | (n57082 & n57333);
  assign n57335 = n33000 | n33495;
  assign n57336 = n57082 | n57335;
  assign n33498 = ~n57334 & n57336;
  assign n33499 = x131 & x220;
  assign n33500 = n33498 & n33499;
  assign n33501 = n33498 | n33499;
  assign n33502 = ~n33500 & n33501;
  assign n57337 = n33007 & n33502;
  assign n57338 = (n33502 & n57086) | (n33502 & n57337) | (n57086 & n57337);
  assign n57339 = n33007 | n33502;
  assign n57340 = n57086 | n57339;
  assign n33505 = ~n57338 & n57340;
  assign n33506 = x130 & x221;
  assign n33507 = n33505 & n33506;
  assign n33508 = n33505 | n33506;
  assign n33509 = ~n33507 & n33508;
  assign n57341 = n33014 & n33509;
  assign n57342 = (n33509 & n57091) | (n33509 & n57341) | (n57091 & n57341);
  assign n57343 = n33014 | n33509;
  assign n57344 = n57091 | n57343;
  assign n33512 = ~n57342 & n57344;
  assign n33513 = x129 & x222;
  assign n33514 = n33512 & n33513;
  assign n33515 = n33512 | n33513;
  assign n33516 = ~n33514 & n33515;
  assign n57125 = n33021 | n33023;
  assign n57345 = n33516 & n57125;
  assign n57346 = n33021 & n33516;
  assign n57347 = (n56861 & n57345) | (n56861 & n57346) | (n57345 & n57346);
  assign n57348 = n33516 | n57125;
  assign n57349 = n33021 | n33516;
  assign n57350 = (n56861 & n57348) | (n56861 & n57349) | (n57348 & n57349);
  assign n33519 = ~n57347 & n57350;
  assign n33520 = x128 & x223;
  assign n33521 = n33519 & n33520;
  assign n33522 = n33519 | n33520;
  assign n33523 = ~n33521 & n33522;
  assign n57123 = n33028 | n33030;
  assign n70920 = n33523 & n57123;
  assign n70921 = n33028 & n33523;
  assign n70922 = (n56859 & n70920) | (n56859 & n70921) | (n70920 & n70921);
  assign n70923 = n33523 | n57123;
  assign n70924 = n33028 | n33523;
  assign n70925 = (n56859 & n70923) | (n56859 & n70924) | (n70923 & n70924);
  assign n33526 = ~n70922 & n70925;
  assign n33527 = x127 & x224;
  assign n33528 = n33526 & n33527;
  assign n33529 = n33526 | n33527;
  assign n33530 = ~n33528 & n33529;
  assign n57121 = n33035 | n33037;
  assign n70926 = n33530 & n57121;
  assign n70927 = n33035 & n33530;
  assign n70928 = (n56857 & n70926) | (n56857 & n70927) | (n70926 & n70927);
  assign n70929 = n33530 | n57121;
  assign n70930 = n33035 | n33530;
  assign n70931 = (n56857 & n70929) | (n56857 & n70930) | (n70929 & n70930);
  assign n33533 = ~n70928 & n70931;
  assign n33534 = x126 & x225;
  assign n33535 = n33533 & n33534;
  assign n33536 = n33533 | n33534;
  assign n33537 = ~n33535 & n33536;
  assign n33538 = n57120 & n33537;
  assign n33539 = n57120 | n33537;
  assign n33540 = ~n33538 & n33539;
  assign n33541 = x125 & x226;
  assign n33542 = n33540 & n33541;
  assign n33543 = n33540 | n33541;
  assign n33544 = ~n33542 & n33543;
  assign n33545 = n57118 & n33544;
  assign n33546 = n57118 | n33544;
  assign n33547 = ~n33545 & n33546;
  assign n33548 = x124 & x227;
  assign n33549 = n33547 & n33548;
  assign n33550 = n33547 | n33548;
  assign n33551 = ~n33549 & n33550;
  assign n33552 = n57116 & n33551;
  assign n33553 = n57116 | n33551;
  assign n33554 = ~n33552 & n33553;
  assign n33555 = x123 & x228;
  assign n33556 = n33554 & n33555;
  assign n33557 = n33554 | n33555;
  assign n33558 = ~n33556 & n33557;
  assign n33559 = n57114 & n33558;
  assign n33560 = n57114 | n33558;
  assign n33561 = ~n33559 & n33560;
  assign n33562 = x122 & x229;
  assign n33563 = n33561 & n33562;
  assign n33564 = n33561 | n33562;
  assign n33565 = ~n33563 & n33564;
  assign n33566 = n57112 & n33565;
  assign n33567 = n57112 | n33565;
  assign n33568 = ~n33566 & n33567;
  assign n33569 = x121 & x230;
  assign n33570 = n33568 & n33569;
  assign n33571 = n33568 | n33569;
  assign n33572 = ~n33570 & n33571;
  assign n33573 = n57110 & n33572;
  assign n33574 = n57110 | n33572;
  assign n33575 = ~n33573 & n33574;
  assign n33576 = x120 & x231;
  assign n33577 = n33575 & n33576;
  assign n33578 = n33575 | n33576;
  assign n33579 = ~n33577 & n33578;
  assign n33580 = n57108 & n33579;
  assign n33581 = n57108 | n33579;
  assign n33582 = ~n33580 & n33581;
  assign n33583 = x119 & x232;
  assign n33584 = n33582 & n33583;
  assign n33585 = n33582 | n33583;
  assign n33586 = ~n33584 & n33585;
  assign n33587 = n57106 & n33586;
  assign n33588 = n57106 | n33586;
  assign n33589 = ~n33587 & n33588;
  assign n33590 = x118 & x233;
  assign n33591 = n33589 & n33590;
  assign n33592 = n33589 | n33590;
  assign n33593 = ~n33591 & n33592;
  assign n33594 = n57104 & n33593;
  assign n33595 = n57104 | n33593;
  assign n33596 = ~n33594 & n33595;
  assign n33597 = x117 & x234;
  assign n33598 = n33596 & n33597;
  assign n33599 = n33596 | n33597;
  assign n33600 = ~n33598 & n33599;
  assign n33601 = n57102 & n33600;
  assign n33602 = n57102 | n33600;
  assign n33603 = ~n33601 & n33602;
  assign n33604 = x116 & x235;
  assign n33605 = n33603 & n33604;
  assign n33606 = n33603 | n33604;
  assign n33607 = ~n33605 & n33606;
  assign n33608 = n57100 & n33607;
  assign n33609 = n57100 | n33607;
  assign n33610 = ~n33608 & n33609;
  assign n33611 = x115 & x236;
  assign n33612 = n33610 & n33611;
  assign n33613 = n33610 | n33611;
  assign n33614 = ~n33612 & n33613;
  assign n33615 = n57098 & n33614;
  assign n33616 = n57098 | n33614;
  assign n33617 = ~n33615 & n33616;
  assign n33618 = x114 & x237;
  assign n33619 = n33617 & n33618;
  assign n33620 = n33617 | n33618;
  assign n33621 = ~n33619 & n33620;
  assign n33622 = n57096 & n33621;
  assign n33623 = n57096 | n33621;
  assign n33624 = ~n33622 & n33623;
  assign n33625 = x113 & x238;
  assign n33626 = n33624 & n33625;
  assign n33627 = n33624 | n33625;
  assign n33628 = ~n33626 & n33627;
  assign n33629 = n33133 & n33628;
  assign n33630 = n33133 | n33628;
  assign n33631 = ~n33629 & n33630;
  assign n33632 = x112 & x239;
  assign n33633 = n33631 & n33632;
  assign n33634 = n33631 | n33632;
  assign n33635 = ~n33633 & n33634;
  assign n70932 = n33133 | n33625;
  assign n70933 = (n33133 & n33624) | (n33133 & n70932) | (n33624 & n70932);
  assign n57352 = (n33626 & n33628) | (n33626 & n70933) | (n33628 & n70933);
  assign n70934 = n33619 | n57096;
  assign n70935 = (n33619 & n33621) | (n33619 & n70934) | (n33621 & n70934);
  assign n33638 = n33612 | n33615;
  assign n33639 = n33605 | n33608;
  assign n33640 = n33598 | n33601;
  assign n33641 = n33591 | n33594;
  assign n33642 = n33584 | n33587;
  assign n33643 = n33577 | n33580;
  assign n33644 = n33570 | n33573;
  assign n33645 = n33563 | n33566;
  assign n33646 = n33556 | n33559;
  assign n57353 = n33549 | n33551;
  assign n57354 = (n33549 & n57116) | (n33549 & n57353) | (n57116 & n57353);
  assign n57355 = n33542 | n33544;
  assign n57356 = (n33542 & n57118) | (n33542 & n57355) | (n57118 & n57355);
  assign n57122 = (n33035 & n56857) | (n33035 & n57121) | (n56857 & n57121);
  assign n57124 = (n33028 & n56859) | (n33028 & n57123) | (n56859 & n57123);
  assign n57369 = n33360 | n33362;
  assign n70938 = n32867 | n33360;
  assign n70939 = (n33360 & n33362) | (n33360 & n70938) | (n33362 & n70938);
  assign n70940 = (n57008 & n57369) | (n57008 & n70939) | (n57369 & n70939);
  assign n70941 = (n57007 & n57369) | (n57007 & n70939) | (n57369 & n70939);
  assign n70942 = (n70496 & n70940) | (n70496 & n70941) | (n70940 & n70941);
  assign n57374 = n33339 | n33341;
  assign n70943 = n32846 | n33339;
  assign n70944 = (n33339 & n33341) | (n33339 & n70943) | (n33341 & n70943);
  assign n70945 = (n56998 & n57374) | (n56998 & n70944) | (n57374 & n70944);
  assign n70946 = (n56997 & n57374) | (n56997 & n70944) | (n57374 & n70944);
  assign n70947 = (n70501 & n70945) | (n70501 & n70946) | (n70945 & n70946);
  assign n57141 = (n56732 & n70801) | (n56732 & n57140) | (n70801 & n57140);
  assign n57379 = n33318 | n33320;
  assign n70948 = n32825 | n33318;
  assign n70949 = (n33318 & n33320) | (n33318 & n70948) | (n33320 & n70948);
  assign n70950 = (n56988 & n57379) | (n56988 & n70949) | (n57379 & n70949);
  assign n70951 = (n56987 & n57379) | (n56987 & n70949) | (n57379 & n70949);
  assign n70952 = (n56637 & n70950) | (n56637 & n70951) | (n70950 & n70951);
  assign n57146 = (n56722 & n70803) | (n56722 & n57145) | (n70803 & n57145);
  assign n57384 = n33297 | n33299;
  assign n70953 = n32804 | n33297;
  assign n70954 = (n33297 & n33299) | (n33297 & n70953) | (n33299 & n70953);
  assign n70955 = (n56978 & n57384) | (n56978 & n70954) | (n57384 & n70954);
  assign n70956 = (n56977 & n57384) | (n56977 & n70954) | (n57384 & n70954);
  assign n70957 = (n56642 & n70955) | (n56642 & n70956) | (n70955 & n70956);
  assign n57151 = (n56712 & n70805) | (n56712 & n57150) | (n70805 & n57150);
  assign n70958 = n32776 | n33269;
  assign n70959 = (n33269 & n33271) | (n33269 & n70958) | (n33271 & n70958);
  assign n70960 = n33269 | n33271;
  assign n70961 = (n33269 & n57155) | (n33269 & n70960) | (n57155 & n70960);
  assign n70962 = (n56890 & n70959) | (n56890 & n70961) | (n70959 & n70961);
  assign n70963 = (n70677 & n70959) | (n70677 & n70961) | (n70959 & n70961);
  assign n70964 = (n56401 & n70962) | (n56401 & n70963) | (n70962 & n70963);
  assign n33698 = x175 & x177;
  assign n70973 = n32706 | n33199;
  assign n70974 = (n33199 & n33201) | (n33199 & n70973) | (n33201 & n70973);
  assign n57419 = n33698 & n70974;
  assign n70975 = n33199 & n33698;
  assign n70976 = (n33201 & n33698) | (n33201 & n70975) | (n33698 & n70975);
  assign n57421 = (n70695 & n57419) | (n70695 & n70976) | (n57419 & n70976);
  assign n57422 = n33698 | n70974;
  assign n70977 = n33199 | n33698;
  assign n70978 = n33201 | n70977;
  assign n57424 = (n70695 & n57422) | (n70695 & n70978) | (n57422 & n70978);
  assign n33701 = ~n57421 & n57424;
  assign n33702 = x174 & x178;
  assign n33703 = n33701 & n33702;
  assign n33704 = n33701 | n33702;
  assign n33705 = ~n33703 & n33704;
  assign n70979 = n33206 | n33208;
  assign n70980 = (n33206 & n70824) | (n33206 & n70979) | (n70824 & n70979);
  assign n57425 = n33705 & n70980;
  assign n70981 = (n33206 & n70825) | (n33206 & n70979) | (n70825 & n70979);
  assign n57426 = n33705 & n70981;
  assign n70982 = (n57425 & n57426) | (n57425 & n70398) | (n57426 & n70398);
  assign n70983 = (n57425 & n57426) | (n57425 & n70402) | (n57426 & n70402);
  assign n70984 = (n69887 & n70982) | (n69887 & n70983) | (n70982 & n70983);
  assign n57428 = n33705 | n70980;
  assign n57429 = n33705 | n70981;
  assign n70985 = (n57428 & n57429) | (n57428 & n70398) | (n57429 & n70398);
  assign n70986 = (n57428 & n57429) | (n57428 & n70402) | (n57429 & n70402);
  assign n70987 = (n69887 & n70985) | (n69887 & n70986) | (n70985 & n70986);
  assign n33708 = ~n70984 & n70987;
  assign n33709 = x173 & x179;
  assign n33710 = n33708 & n33709;
  assign n33711 = n33708 | n33709;
  assign n33712 = ~n33710 & n33711;
  assign n70988 = n33213 | n33215;
  assign n70993 = (n33213 & n70835) | (n33213 & n70988) | (n70835 & n70988);
  assign n57432 = n33712 & n70993;
  assign n70990 = n33712 & n70988;
  assign n70991 = n33213 & n33712;
  assign n70992 = (n70833 & n70990) | (n70833 & n70991) | (n70990 & n70991);
  assign n70994 = (n57432 & n70524) | (n57432 & n70992) | (n70524 & n70992);
  assign n70995 = (n57432 & n70523) | (n57432 & n70992) | (n70523 & n70992);
  assign n70996 = (n70013 & n70994) | (n70013 & n70995) | (n70994 & n70995);
  assign n57435 = n33712 | n70993;
  assign n70997 = n33712 | n70988;
  assign n70998 = n33213 | n33712;
  assign n70999 = (n70833 & n70997) | (n70833 & n70998) | (n70997 & n70998);
  assign n71000 = (n57435 & n70524) | (n57435 & n70999) | (n70524 & n70999);
  assign n71001 = (n57435 & n70523) | (n57435 & n70999) | (n70523 & n70999);
  assign n71002 = (n70013 & n71000) | (n70013 & n71001) | (n71000 & n71001);
  assign n33715 = ~n70996 & n71002;
  assign n33716 = x172 & x180;
  assign n33717 = n33715 & n33716;
  assign n33718 = n33715 | n33716;
  assign n33719 = ~n33717 & n33718;
  assign n70967 = n33220 | n33222;
  assign n70968 = (n33220 & n70843) | (n33220 & n70967) | (n70843 & n70967);
  assign n70969 = (n33220 & n70845) | (n33220 & n70967) | (n70845 & n70967);
  assign n70971 = (n70521 & n70968) | (n70521 & n70969) | (n70968 & n70969);
  assign n71003 = n33719 & n70971;
  assign n70970 = (n70520 & n70968) | (n70520 & n70969) | (n70968 & n70969);
  assign n71004 = n33719 & n70970;
  assign n71005 = (n70133 & n71003) | (n70133 & n71004) | (n71003 & n71004);
  assign n71006 = n33719 | n70971;
  assign n71007 = n33719 | n70970;
  assign n71008 = (n70133 & n71006) | (n70133 & n71007) | (n71006 & n71007);
  assign n33722 = ~n71005 & n71008;
  assign n33723 = x171 & x181;
  assign n33724 = n33722 & n33723;
  assign n33725 = n33722 | n33723;
  assign n33726 = ~n33724 & n33725;
  assign n57405 = n33227 | n33229;
  assign n57437 = n33726 & n57405;
  assign n57438 = n33227 & n33726;
  assign n57439 = (n70822 & n57437) | (n70822 & n57438) | (n57437 & n57438);
  assign n57440 = n33726 | n57405;
  assign n57441 = n33227 | n33726;
  assign n57442 = (n70822 & n57440) | (n70822 & n57441) | (n57440 & n57441);
  assign n33729 = ~n57439 & n57442;
  assign n33730 = x170 & x182;
  assign n33731 = n33729 & n33730;
  assign n33732 = n33729 | n33730;
  assign n33733 = ~n33731 & n33732;
  assign n57403 = n33234 | n57206;
  assign n71009 = n33733 & n57403;
  assign n57402 = n33234 | n57205;
  assign n71010 = n33733 & n57402;
  assign n71011 = (n70574 & n71009) | (n70574 & n71010) | (n71009 & n71010);
  assign n71012 = n33733 | n57403;
  assign n71013 = n33733 | n57402;
  assign n71014 = (n70574 & n71012) | (n70574 & n71013) | (n71012 & n71013);
  assign n33736 = ~n71011 & n71014;
  assign n33737 = x169 & x183;
  assign n33738 = n33736 & n33737;
  assign n33739 = n33736 | n33737;
  assign n33740 = ~n33738 & n33739;
  assign n57400 = n33241 | n33243;
  assign n57443 = n33740 & n57400;
  assign n57444 = n33241 & n33740;
  assign n71015 = (n57166 & n57443) | (n57166 & n57444) | (n57443 & n57444);
  assign n71016 = (n57165 & n57443) | (n57165 & n57444) | (n57443 & n57444);
  assign n71017 = (n70430 & n71015) | (n70430 & n71016) | (n71015 & n71016);
  assign n57446 = n33740 | n57400;
  assign n57447 = n33241 | n33740;
  assign n71018 = (n57166 & n57446) | (n57166 & n57447) | (n57446 & n57447);
  assign n71019 = (n57165 & n57446) | (n57165 & n57447) | (n57446 & n57447);
  assign n71020 = (n70430 & n71018) | (n70430 & n71019) | (n71018 & n71019);
  assign n33743 = ~n71017 & n71020;
  assign n33744 = x168 & x184;
  assign n33745 = n33743 & n33744;
  assign n33746 = n33743 | n33744;
  assign n33747 = ~n33745 & n33746;
  assign n57398 = n33248 | n33250;
  assign n57449 = n33747 & n57398;
  assign n57450 = n33248 & n33747;
  assign n57451 = (n70816 & n57449) | (n70816 & n57450) | (n57449 & n57450);
  assign n57452 = n33747 | n57398;
  assign n57453 = n33248 | n33747;
  assign n57454 = (n70816 & n57452) | (n70816 & n57453) | (n57452 & n57453);
  assign n33750 = ~n57451 & n57454;
  assign n33751 = x167 & x185;
  assign n33752 = n33750 & n33751;
  assign n33753 = n33750 | n33751;
  assign n33754 = ~n33752 & n33753;
  assign n57396 = n33255 | n57211;
  assign n71021 = n33754 & n57396;
  assign n70965 = n32762 | n33255;
  assign n70966 = (n33255 & n33257) | (n33255 & n70965) | (n33257 & n70965);
  assign n71022 = n33754 & n70966;
  assign n71023 = (n70684 & n71021) | (n70684 & n71022) | (n71021 & n71022);
  assign n71024 = n33754 | n57396;
  assign n71025 = n33754 | n70966;
  assign n71026 = (n70684 & n71024) | (n70684 & n71025) | (n71024 & n71025);
  assign n33757 = ~n71023 & n71026;
  assign n33758 = x166 & x186;
  assign n33759 = n33757 & n33758;
  assign n33760 = n33757 | n33758;
  assign n33761 = ~n33759 & n33760;
  assign n57393 = n33262 | n33264;
  assign n57455 = n33761 & n57393;
  assign n57456 = n33262 & n33761;
  assign n71027 = (n57158 & n57455) | (n57158 & n57456) | (n57455 & n57456);
  assign n71028 = (n57455 & n57456) | (n57455 & n70809) | (n57456 & n70809);
  assign n71029 = (n70514 & n71027) | (n70514 & n71028) | (n71027 & n71028);
  assign n57458 = n33761 | n57393;
  assign n57459 = n33262 | n33761;
  assign n71030 = (n57158 & n57458) | (n57158 & n57459) | (n57458 & n57459);
  assign n71031 = (n57458 & n57459) | (n57458 & n70809) | (n57459 & n70809);
  assign n71032 = (n70514 & n71030) | (n70514 & n71031) | (n71030 & n71031);
  assign n33764 = ~n71029 & n71032;
  assign n33765 = x165 & x187;
  assign n33766 = n33764 & n33765;
  assign n33767 = n33764 | n33765;
  assign n33768 = ~n33766 & n33767;
  assign n33769 = n70964 & n33768;
  assign n33770 = n70964 | n33768;
  assign n33771 = ~n33769 & n33770;
  assign n33772 = x164 & x188;
  assign n33773 = n33771 & n33772;
  assign n33774 = n33771 | n33772;
  assign n33775 = ~n33773 & n33774;
  assign n57388 = n33276 | n33278;
  assign n57461 = n33775 & n57388;
  assign n57462 = n33276 & n33775;
  assign n71033 = (n57153 & n57461) | (n57153 & n57462) | (n57461 & n57462);
  assign n71034 = (n57461 & n57462) | (n57461 & n70807) | (n57462 & n70807);
  assign n71035 = (n56647 & n71033) | (n56647 & n71034) | (n71033 & n71034);
  assign n57464 = n33775 | n57388;
  assign n57465 = n33276 | n33775;
  assign n71036 = (n57153 & n57464) | (n57153 & n57465) | (n57464 & n57465);
  assign n71037 = (n57464 & n57465) | (n57464 & n70807) | (n57465 & n70807);
  assign n71038 = (n56647 & n71036) | (n56647 & n71037) | (n71036 & n71037);
  assign n33778 = ~n71035 & n71038;
  assign n33779 = x163 & x189;
  assign n33780 = n33778 & n33779;
  assign n33781 = n33778 | n33779;
  assign n33782 = ~n33780 & n33781;
  assign n57386 = n33283 | n33285;
  assign n57467 = n33782 & n57386;
  assign n57468 = n33283 & n33782;
  assign n57469 = (n57151 & n57467) | (n57151 & n57468) | (n57467 & n57468);
  assign n57470 = n33782 | n57386;
  assign n57471 = n33283 | n33782;
  assign n57472 = (n57151 & n57470) | (n57151 & n57471) | (n57470 & n57471);
  assign n33785 = ~n57469 & n57472;
  assign n33786 = x162 & x190;
  assign n33787 = n33785 & n33786;
  assign n33788 = n33785 | n33786;
  assign n33789 = ~n33787 & n33788;
  assign n57473 = n33290 & n33789;
  assign n57474 = (n33789 & n57225) | (n33789 & n57473) | (n57225 & n57473);
  assign n57475 = n33290 | n33789;
  assign n57476 = n57225 | n57475;
  assign n33792 = ~n57474 & n57476;
  assign n33793 = x161 & x191;
  assign n33794 = n33792 & n33793;
  assign n33795 = n33792 | n33793;
  assign n33796 = ~n33794 & n33795;
  assign n33797 = n70957 & n33796;
  assign n33798 = n70957 | n33796;
  assign n33799 = ~n33797 & n33798;
  assign n33800 = x160 & x192;
  assign n33801 = n33799 & n33800;
  assign n33802 = n33799 | n33800;
  assign n33803 = ~n33801 & n33802;
  assign n57381 = n33304 | n33306;
  assign n57477 = n33803 & n57381;
  assign n57478 = n33304 & n33803;
  assign n57479 = (n57146 & n57477) | (n57146 & n57478) | (n57477 & n57478);
  assign n57480 = n33803 | n57381;
  assign n57481 = n33304 | n33803;
  assign n57482 = (n57146 & n57480) | (n57146 & n57481) | (n57480 & n57481);
  assign n33806 = ~n57479 & n57482;
  assign n33807 = x159 & x193;
  assign n33808 = n33806 & n33807;
  assign n33809 = n33806 | n33807;
  assign n33810 = ~n33808 & n33809;
  assign n57483 = n33311 & n33810;
  assign n57484 = (n33810 & n57235) | (n33810 & n57483) | (n57235 & n57483);
  assign n57485 = n33311 | n33810;
  assign n57486 = n57235 | n57485;
  assign n33813 = ~n57484 & n57486;
  assign n33814 = x158 & x194;
  assign n33815 = n33813 & n33814;
  assign n33816 = n33813 | n33814;
  assign n33817 = ~n33815 & n33816;
  assign n33818 = n70952 & n33817;
  assign n33819 = n70952 | n33817;
  assign n33820 = ~n33818 & n33819;
  assign n33821 = x157 & x195;
  assign n33822 = n33820 & n33821;
  assign n33823 = n33820 | n33821;
  assign n33824 = ~n33822 & n33823;
  assign n57376 = n33325 | n33327;
  assign n57487 = n33824 & n57376;
  assign n57488 = n33325 & n33824;
  assign n57489 = (n57141 & n57487) | (n57141 & n57488) | (n57487 & n57488);
  assign n57490 = n33824 | n57376;
  assign n57491 = n33325 | n33824;
  assign n57492 = (n57141 & n57490) | (n57141 & n57491) | (n57490 & n57491);
  assign n33827 = ~n57489 & n57492;
  assign n33828 = x156 & x196;
  assign n33829 = n33827 & n33828;
  assign n33830 = n33827 | n33828;
  assign n33831 = ~n33829 & n33830;
  assign n57493 = n33332 & n33831;
  assign n57494 = (n33831 & n57245) | (n33831 & n57493) | (n57245 & n57493);
  assign n57495 = n33332 | n33831;
  assign n57496 = n57245 | n57495;
  assign n33834 = ~n57494 & n57496;
  assign n33835 = x155 & x197;
  assign n33836 = n33834 & n33835;
  assign n33837 = n33834 | n33835;
  assign n33838 = ~n33836 & n33837;
  assign n33839 = n70947 & n33838;
  assign n33840 = n70947 | n33838;
  assign n33841 = ~n33839 & n33840;
  assign n33842 = x154 & x198;
  assign n33843 = n33841 & n33842;
  assign n33844 = n33841 | n33842;
  assign n33845 = ~n33843 & n33844;
  assign n57371 = n33346 | n33348;
  assign n57497 = n33845 & n57371;
  assign n57498 = n33346 & n33845;
  assign n57499 = (n70799 & n57497) | (n70799 & n57498) | (n57497 & n57498);
  assign n57500 = n33845 | n57371;
  assign n57501 = n33346 | n33845;
  assign n57502 = (n70799 & n57500) | (n70799 & n57501) | (n57500 & n57501);
  assign n33848 = ~n57499 & n57502;
  assign n33849 = x153 & x199;
  assign n33850 = n33848 & n33849;
  assign n33851 = n33848 | n33849;
  assign n33852 = ~n33850 & n33851;
  assign n57503 = n33353 & n33852;
  assign n71039 = (n33852 & n57254) | (n33852 & n57503) | (n57254 & n57503);
  assign n71040 = (n33852 & n57253) | (n33852 & n57503) | (n57253 & n57503);
  assign n71041 = (n70660 & n71039) | (n70660 & n71040) | (n71039 & n71040);
  assign n57505 = n33353 | n33852;
  assign n71042 = n57254 | n57505;
  assign n71043 = n57253 | n57505;
  assign n71044 = (n70660 & n71042) | (n70660 & n71043) | (n71042 & n71043);
  assign n33855 = ~n71041 & n71044;
  assign n33856 = x152 & x200;
  assign n33857 = n33855 & n33856;
  assign n33858 = n33855 | n33856;
  assign n33859 = ~n33857 & n33858;
  assign n33860 = n70942 & n33859;
  assign n33861 = n70942 | n33859;
  assign n33862 = ~n33860 & n33861;
  assign n33863 = x151 & x201;
  assign n33864 = n33862 & n33863;
  assign n33865 = n33862 | n33863;
  assign n33866 = ~n33864 & n33865;
  assign n57366 = n33367 | n33369;
  assign n57507 = n33866 & n57366;
  assign n57508 = n33367 & n33866;
  assign n57509 = (n70794 & n57507) | (n70794 & n57508) | (n57507 & n57508);
  assign n57510 = n33866 | n57366;
  assign n57511 = n33367 | n33866;
  assign n57512 = (n70794 & n57510) | (n70794 & n57511) | (n57510 & n57511);
  assign n33869 = ~n57509 & n57512;
  assign n33870 = x150 & x202;
  assign n33871 = n33869 & n33870;
  assign n33872 = n33869 | n33870;
  assign n33873 = ~n33871 & n33872;
  assign n57513 = n33374 & n33873;
  assign n71045 = (n33873 & n57264) | (n33873 & n57513) | (n57264 & n57513);
  assign n71046 = (n33873 & n57263) | (n33873 & n57513) | (n57263 & n57513);
  assign n71047 = (n56866 & n71045) | (n56866 & n71046) | (n71045 & n71046);
  assign n57515 = n33374 | n33873;
  assign n71048 = n57264 | n57515;
  assign n71049 = n57263 | n57515;
  assign n71050 = (n56866 & n71048) | (n56866 & n71049) | (n71048 & n71049);
  assign n33876 = ~n71047 & n71050;
  assign n33877 = x149 & x203;
  assign n33878 = n33876 & n33877;
  assign n33879 = n33876 | n33877;
  assign n33880 = ~n33878 & n33879;
  assign n57364 = n33381 | n33383;
  assign n71051 = n33880 & n57364;
  assign n70936 = n32888 | n33381;
  assign n70937 = (n33381 & n33383) | (n33381 & n70936) | (n33383 & n70936);
  assign n71052 = n33880 & n70937;
  assign n71053 = (n70774 & n71051) | (n70774 & n71052) | (n71051 & n71052);
  assign n71054 = n33880 | n57364;
  assign n71055 = n33880 | n70937;
  assign n71056 = (n70774 & n71054) | (n70774 & n71055) | (n71054 & n71055);
  assign n33883 = ~n71053 & n71056;
  assign n33884 = x148 & x204;
  assign n33885 = n33883 & n33884;
  assign n33886 = n33883 | n33884;
  assign n33887 = ~n33885 & n33886;
  assign n57517 = n33388 & n33887;
  assign n71057 = (n33887 & n57273) | (n33887 & n57517) | (n57273 & n57517);
  assign n71058 = (n33390 & n33887) | (n33390 & n57517) | (n33887 & n57517);
  assign n71059 = (n57022 & n71057) | (n57022 & n71058) | (n71057 & n71058);
  assign n57519 = n33388 | n33887;
  assign n71060 = n57273 | n57519;
  assign n71061 = n33390 | n57519;
  assign n71062 = (n57022 & n71060) | (n57022 & n71061) | (n71060 & n71061);
  assign n33890 = ~n71059 & n71062;
  assign n33891 = x147 & x205;
  assign n33892 = n33890 & n33891;
  assign n33893 = n33890 | n33891;
  assign n33894 = ~n33892 & n33893;
  assign n57521 = n33395 & n33894;
  assign n57522 = (n33894 & n57278) | (n33894 & n57521) | (n57278 & n57521);
  assign n57523 = n33395 | n33894;
  assign n57524 = n57278 | n57523;
  assign n33897 = ~n57522 & n57524;
  assign n33898 = x146 & x206;
  assign n33899 = n33897 & n33898;
  assign n33900 = n33897 | n33898;
  assign n33901 = ~n33899 & n33900;
  assign n57525 = n33402 & n33901;
  assign n57526 = (n33901 & n57282) | (n33901 & n57525) | (n57282 & n57525);
  assign n57527 = n33402 | n33901;
  assign n57528 = n57282 | n57527;
  assign n33904 = ~n57526 & n57528;
  assign n33905 = x145 & x207;
  assign n33906 = n33904 & n33905;
  assign n33907 = n33904 | n33905;
  assign n33908 = ~n33906 & n33907;
  assign n57529 = n33409 & n33908;
  assign n57530 = (n33908 & n57286) | (n33908 & n57529) | (n57286 & n57529);
  assign n57531 = n33409 | n33908;
  assign n57532 = n57286 | n57531;
  assign n33911 = ~n57530 & n57532;
  assign n33912 = x144 & x208;
  assign n33913 = n33911 & n33912;
  assign n33914 = n33911 | n33912;
  assign n33915 = ~n33913 & n33914;
  assign n57533 = n33416 & n33915;
  assign n57534 = (n33915 & n57290) | (n33915 & n57533) | (n57290 & n57533);
  assign n57535 = n33416 | n33915;
  assign n57536 = n57290 | n57535;
  assign n33918 = ~n57534 & n57536;
  assign n33919 = x143 & x209;
  assign n33920 = n33918 & n33919;
  assign n33921 = n33918 | n33919;
  assign n33922 = ~n33920 & n33921;
  assign n57537 = n33423 & n33922;
  assign n57538 = (n33922 & n57294) | (n33922 & n57537) | (n57294 & n57537);
  assign n57539 = n33423 | n33922;
  assign n57540 = n57294 | n57539;
  assign n33925 = ~n57538 & n57540;
  assign n33926 = x142 & x210;
  assign n33927 = n33925 & n33926;
  assign n33928 = n33925 | n33926;
  assign n33929 = ~n33927 & n33928;
  assign n57541 = n33430 & n33929;
  assign n57542 = (n33929 & n57298) | (n33929 & n57541) | (n57298 & n57541);
  assign n57543 = n33430 | n33929;
  assign n57544 = n57298 | n57543;
  assign n33932 = ~n57542 & n57544;
  assign n33933 = x141 & x211;
  assign n33934 = n33932 & n33933;
  assign n33935 = n33932 | n33933;
  assign n33936 = ~n33934 & n33935;
  assign n57545 = n33437 & n33936;
  assign n57546 = (n33936 & n57302) | (n33936 & n57545) | (n57302 & n57545);
  assign n57547 = n33437 | n33936;
  assign n57548 = n57302 | n57547;
  assign n33939 = ~n57546 & n57548;
  assign n33940 = x140 & x212;
  assign n33941 = n33939 & n33940;
  assign n33942 = n33939 | n33940;
  assign n33943 = ~n33941 & n33942;
  assign n57549 = n33444 & n33943;
  assign n57550 = (n33943 & n57306) | (n33943 & n57549) | (n57306 & n57549);
  assign n57551 = n33444 | n33943;
  assign n57552 = n57306 | n57551;
  assign n33946 = ~n57550 & n57552;
  assign n33947 = x139 & x213;
  assign n33948 = n33946 & n33947;
  assign n33949 = n33946 | n33947;
  assign n33950 = ~n33948 & n33949;
  assign n57553 = n33451 & n33950;
  assign n57554 = (n33950 & n57310) | (n33950 & n57553) | (n57310 & n57553);
  assign n57555 = n33451 | n33950;
  assign n57556 = n57310 | n57555;
  assign n33953 = ~n57554 & n57556;
  assign n33954 = x138 & x214;
  assign n33955 = n33953 & n33954;
  assign n33956 = n33953 | n33954;
  assign n33957 = ~n33955 & n33956;
  assign n57557 = n33458 & n33957;
  assign n57558 = (n33957 & n57314) | (n33957 & n57557) | (n57314 & n57557);
  assign n57559 = n33458 | n33957;
  assign n57560 = n57314 | n57559;
  assign n33960 = ~n57558 & n57560;
  assign n33961 = x137 & x215;
  assign n33962 = n33960 & n33961;
  assign n33963 = n33960 | n33961;
  assign n33964 = ~n33962 & n33963;
  assign n57561 = n33465 & n33964;
  assign n57562 = (n33964 & n57318) | (n33964 & n57561) | (n57318 & n57561);
  assign n57563 = n33465 | n33964;
  assign n57564 = n57318 | n57563;
  assign n33967 = ~n57562 & n57564;
  assign n33968 = x136 & x216;
  assign n33969 = n33967 & n33968;
  assign n33970 = n33967 | n33968;
  assign n33971 = ~n33969 & n33970;
  assign n57565 = n33472 & n33971;
  assign n57566 = (n33971 & n57322) | (n33971 & n57565) | (n57322 & n57565);
  assign n57567 = n33472 | n33971;
  assign n57568 = n57322 | n57567;
  assign n33974 = ~n57566 & n57568;
  assign n33975 = x135 & x217;
  assign n33976 = n33974 & n33975;
  assign n33977 = n33974 | n33975;
  assign n33978 = ~n33976 & n33977;
  assign n57569 = n33479 & n33978;
  assign n57570 = (n33978 & n57326) | (n33978 & n57569) | (n57326 & n57569);
  assign n57571 = n33479 | n33978;
  assign n57572 = n57326 | n57571;
  assign n33981 = ~n57570 & n57572;
  assign n33982 = x134 & x218;
  assign n33983 = n33981 & n33982;
  assign n33984 = n33981 | n33982;
  assign n33985 = ~n33983 & n33984;
  assign n57573 = n33486 & n33985;
  assign n57574 = (n33985 & n57330) | (n33985 & n57573) | (n57330 & n57573);
  assign n57575 = n33486 | n33985;
  assign n57576 = n57330 | n57575;
  assign n33988 = ~n57574 & n57576;
  assign n33989 = x133 & x219;
  assign n33990 = n33988 & n33989;
  assign n33991 = n33988 | n33989;
  assign n33992 = ~n33990 & n33991;
  assign n57577 = n33493 & n33992;
  assign n57578 = (n33992 & n57334) | (n33992 & n57577) | (n57334 & n57577);
  assign n57579 = n33493 | n33992;
  assign n57580 = n57334 | n57579;
  assign n33995 = ~n57578 & n57580;
  assign n33996 = x132 & x220;
  assign n33997 = n33995 & n33996;
  assign n33998 = n33995 | n33996;
  assign n33999 = ~n33997 & n33998;
  assign n57581 = n33500 & n33999;
  assign n57582 = (n33999 & n57338) | (n33999 & n57581) | (n57338 & n57581);
  assign n57583 = n33500 | n33999;
  assign n57584 = n57338 | n57583;
  assign n34002 = ~n57582 & n57584;
  assign n34003 = x131 & x221;
  assign n34004 = n34002 & n34003;
  assign n34005 = n34002 | n34003;
  assign n34006 = ~n34004 & n34005;
  assign n57585 = n33507 & n34006;
  assign n57586 = (n34006 & n57342) | (n34006 & n57585) | (n57342 & n57585);
  assign n57587 = n33507 | n34006;
  assign n57588 = n57342 | n57587;
  assign n34009 = ~n57586 & n57588;
  assign n34010 = x130 & x222;
  assign n34011 = n34009 & n34010;
  assign n34012 = n34009 | n34010;
  assign n34013 = ~n34011 & n34012;
  assign n57589 = n33514 & n34013;
  assign n57590 = (n34013 & n57347) | (n34013 & n57589) | (n57347 & n57589);
  assign n57591 = n33514 | n34013;
  assign n57592 = n57347 | n57591;
  assign n34016 = ~n57590 & n57592;
  assign n34017 = x129 & x223;
  assign n34018 = n34016 & n34017;
  assign n34019 = n34016 | n34017;
  assign n34020 = ~n34018 & n34019;
  assign n57361 = n33521 | n33523;
  assign n57593 = n34020 & n57361;
  assign n57594 = n33521 & n34020;
  assign n57595 = (n57124 & n57593) | (n57124 & n57594) | (n57593 & n57594);
  assign n57596 = n34020 | n57361;
  assign n57597 = n33521 | n34020;
  assign n57598 = (n57124 & n57596) | (n57124 & n57597) | (n57596 & n57597);
  assign n34023 = ~n57595 & n57598;
  assign n34024 = x128 & x224;
  assign n34025 = n34023 & n34024;
  assign n34026 = n34023 | n34024;
  assign n34027 = ~n34025 & n34026;
  assign n57359 = n33528 | n33530;
  assign n71063 = n34027 & n57359;
  assign n71064 = n33528 & n34027;
  assign n71065 = (n57122 & n71063) | (n57122 & n71064) | (n71063 & n71064);
  assign n71066 = n34027 | n57359;
  assign n71067 = n33528 | n34027;
  assign n71068 = (n57122 & n71066) | (n57122 & n71067) | (n71066 & n71067);
  assign n34030 = ~n71065 & n71068;
  assign n34031 = x127 & x225;
  assign n34032 = n34030 & n34031;
  assign n34033 = n34030 | n34031;
  assign n34034 = ~n34032 & n34033;
  assign n57357 = n33535 | n33537;
  assign n71069 = n34034 & n57357;
  assign n71070 = n33535 & n34034;
  assign n71071 = (n57120 & n71069) | (n57120 & n71070) | (n71069 & n71070);
  assign n71072 = n34034 | n57357;
  assign n71073 = n33535 | n34034;
  assign n71074 = (n57120 & n71072) | (n57120 & n71073) | (n71072 & n71073);
  assign n34037 = ~n71071 & n71074;
  assign n34038 = x126 & x226;
  assign n34039 = n34037 & n34038;
  assign n34040 = n34037 | n34038;
  assign n34041 = ~n34039 & n34040;
  assign n34042 = n57356 & n34041;
  assign n34043 = n57356 | n34041;
  assign n34044 = ~n34042 & n34043;
  assign n34045 = x125 & x227;
  assign n34046 = n34044 & n34045;
  assign n34047 = n34044 | n34045;
  assign n34048 = ~n34046 & n34047;
  assign n34049 = n57354 & n34048;
  assign n34050 = n57354 | n34048;
  assign n34051 = ~n34049 & n34050;
  assign n34052 = x124 & x228;
  assign n34053 = n34051 & n34052;
  assign n34054 = n34051 | n34052;
  assign n34055 = ~n34053 & n34054;
  assign n34056 = n33646 & n34055;
  assign n34057 = n33646 | n34055;
  assign n34058 = ~n34056 & n34057;
  assign n34059 = x123 & x229;
  assign n34060 = n34058 & n34059;
  assign n34061 = n34058 | n34059;
  assign n34062 = ~n34060 & n34061;
  assign n34063 = n33645 & n34062;
  assign n34064 = n33645 | n34062;
  assign n34065 = ~n34063 & n34064;
  assign n34066 = x122 & x230;
  assign n34067 = n34065 & n34066;
  assign n34068 = n34065 | n34066;
  assign n34069 = ~n34067 & n34068;
  assign n34070 = n33644 & n34069;
  assign n34071 = n33644 | n34069;
  assign n34072 = ~n34070 & n34071;
  assign n34073 = x121 & x231;
  assign n34074 = n34072 & n34073;
  assign n34075 = n34072 | n34073;
  assign n34076 = ~n34074 & n34075;
  assign n34077 = n33643 & n34076;
  assign n34078 = n33643 | n34076;
  assign n34079 = ~n34077 & n34078;
  assign n34080 = x120 & x232;
  assign n34081 = n34079 & n34080;
  assign n34082 = n34079 | n34080;
  assign n34083 = ~n34081 & n34082;
  assign n34084 = n33642 & n34083;
  assign n34085 = n33642 | n34083;
  assign n34086 = ~n34084 & n34085;
  assign n34087 = x119 & x233;
  assign n34088 = n34086 & n34087;
  assign n34089 = n34086 | n34087;
  assign n34090 = ~n34088 & n34089;
  assign n34091 = n33641 & n34090;
  assign n34092 = n33641 | n34090;
  assign n34093 = ~n34091 & n34092;
  assign n34094 = x118 & x234;
  assign n34095 = n34093 & n34094;
  assign n34096 = n34093 | n34094;
  assign n34097 = ~n34095 & n34096;
  assign n34098 = n33640 & n34097;
  assign n34099 = n33640 | n34097;
  assign n34100 = ~n34098 & n34099;
  assign n34101 = x117 & x235;
  assign n34102 = n34100 & n34101;
  assign n34103 = n34100 | n34101;
  assign n34104 = ~n34102 & n34103;
  assign n34105 = n33639 & n34104;
  assign n34106 = n33639 | n34104;
  assign n34107 = ~n34105 & n34106;
  assign n34108 = x116 & x236;
  assign n34109 = n34107 & n34108;
  assign n34110 = n34107 | n34108;
  assign n34111 = ~n34109 & n34110;
  assign n34112 = n33638 & n34111;
  assign n34113 = n33638 | n34111;
  assign n34114 = ~n34112 & n34113;
  assign n34115 = x115 & x237;
  assign n34116 = n34114 & n34115;
  assign n34117 = n34114 | n34115;
  assign n34118 = ~n34116 & n34117;
  assign n34119 = n70935 & n34118;
  assign n34120 = n70935 | n34118;
  assign n34121 = ~n34119 & n34120;
  assign n34122 = x114 & x238;
  assign n34123 = n34121 & n34122;
  assign n34124 = n34121 | n34122;
  assign n34125 = ~n34123 & n34124;
  assign n34126 = n57352 & n34125;
  assign n34127 = n57352 | n34125;
  assign n34128 = ~n34126 & n34127;
  assign n34129 = x113 & x239;
  assign n34130 = n34128 & n34129;
  assign n34131 = n34128 | n34129;
  assign n34132 = ~n34130 & n34131;
  assign n34133 = n33633 & n34132;
  assign n34134 = n33633 | n34132;
  assign n34135 = ~n34133 & n34134;
  assign n71075 = n33633 | n34129;
  assign n71076 = (n33633 & n34128) | (n33633 & n71075) | (n34128 & n71075);
  assign n57600 = (n34130 & n34132) | (n34130 & n71076) | (n34132 & n71076);
  assign n57601 = n34123 | n57352;
  assign n57602 = (n34123 & n34125) | (n34123 & n57601) | (n34125 & n57601);
  assign n71077 = n34116 | n70935;
  assign n71078 = (n34116 & n34118) | (n34116 & n71077) | (n34118 & n71077);
  assign n34139 = n34109 | n34112;
  assign n34140 = n34102 | n34105;
  assign n34141 = n34095 | n34098;
  assign n34142 = n34088 | n34091;
  assign n34143 = n34081 | n34084;
  assign n34144 = n34074 | n34077;
  assign n34145 = n34067 | n34070;
  assign n34146 = n34060 | n34063;
  assign n57603 = n34053 | n34055;
  assign n57604 = (n33646 & n34053) | (n33646 & n57603) | (n34053 & n57603);
  assign n57605 = n34046 | n34048;
  assign n57606 = (n34046 & n57354) | (n34046 & n57605) | (n57354 & n57605);
  assign n57358 = (n33535 & n57120) | (n33535 & n57357) | (n57120 & n57357);
  assign n57360 = (n33528 & n57122) | (n33528 & n57359) | (n57122 & n57359);
  assign n57365 = (n70774 & n70937) | (n70774 & n57364) | (n70937 & n57364);
  assign n57616 = n33871 | n33873;
  assign n71079 = n33374 | n33871;
  assign n71080 = (n33871 & n33873) | (n33871 & n71079) | (n33873 & n71079);
  assign n71081 = (n57264 & n57616) | (n57264 & n71080) | (n57616 & n71080);
  assign n71082 = (n57263 & n57616) | (n57263 & n71080) | (n57616 & n71080);
  assign n71083 = (n56866 & n71081) | (n56866 & n71082) | (n71081 & n71082);
  assign n57621 = n33850 | n33852;
  assign n71084 = n33353 | n33850;
  assign n71085 = (n33850 & n33852) | (n33850 & n71084) | (n33852 & n71084);
  assign n71086 = (n57254 & n57621) | (n57254 & n71085) | (n57621 & n71085);
  assign n71087 = (n57253 & n57621) | (n57253 & n71085) | (n57621 & n71085);
  assign n71088 = (n70660 & n71086) | (n70660 & n71087) | (n71086 & n71087);
  assign n57154 = (n56647 & n70807) | (n56647 & n57153) | (n70807 & n57153);
  assign n71097 = n33262 | n33759;
  assign n71098 = (n33759 & n33761) | (n33759 & n71097) | (n33761 & n71097);
  assign n71099 = n33759 | n33761;
  assign n71100 = (n33759 & n57393) | (n33759 & n71099) | (n57393 & n71099);
  assign n71101 = (n57158 & n71098) | (n57158 & n71100) | (n71098 & n71100);
  assign n71102 = (n70809 & n71098) | (n70809 & n71100) | (n71098 & n71100);
  assign n71103 = (n70514 & n71101) | (n70514 & n71102) | (n71101 & n71102);
  assign n57167 = (n70430 & n57165) | (n70430 & n57166) | (n57165 & n57166);
  assign n34198 = x175 & x178;
  assign n71108 = n33698 & n34198;
  assign n71109 = n70974 & n71108;
  assign n57665 = n34198 & n70976;
  assign n57666 = (n70695 & n71109) | (n70695 & n57665) | (n71109 & n57665);
  assign n71110 = n33698 | n34198;
  assign n71111 = (n34198 & n70974) | (n34198 & n71110) | (n70974 & n71110);
  assign n57668 = n34198 | n70976;
  assign n57669 = (n70695 & n71111) | (n70695 & n57668) | (n71111 & n57668);
  assign n34201 = ~n57666 & n57669;
  assign n71112 = n33703 | n33705;
  assign n71114 = n34201 & n71112;
  assign n71115 = n33703 & n34201;
  assign n71116 = (n70980 & n71114) | (n70980 & n71115) | (n71114 & n71115);
  assign n71118 = (n70981 & n71114) | (n70981 & n71115) | (n71114 & n71115);
  assign n71119 = (n70398 & n71116) | (n70398 & n71118) | (n71116 & n71118);
  assign n71120 = (n70402 & n71116) | (n70402 & n71118) | (n71116 & n71118);
  assign n71121 = (n69887 & n71119) | (n69887 & n71120) | (n71119 & n71120);
  assign n71122 = n34201 | n71112;
  assign n71123 = n33703 | n34201;
  assign n71124 = (n70980 & n71122) | (n70980 & n71123) | (n71122 & n71123);
  assign n71125 = (n70981 & n71122) | (n70981 & n71123) | (n71122 & n71123);
  assign n71126 = (n70398 & n71124) | (n70398 & n71125) | (n71124 & n71125);
  assign n71127 = (n70402 & n71124) | (n70402 & n71125) | (n71124 & n71125);
  assign n71128 = (n69887 & n71126) | (n69887 & n71127) | (n71126 & n71127);
  assign n34204 = ~n71121 & n71128;
  assign n34205 = x174 & x179;
  assign n34206 = n34204 & n34205;
  assign n34207 = n34204 | n34205;
  assign n34208 = ~n34206 & n34207;
  assign n57676 = n33710 & n34208;
  assign n71129 = (n34208 & n57676) | (n34208 & n70995) | (n57676 & n70995);
  assign n71130 = (n34208 & n57676) | (n34208 & n70994) | (n57676 & n70994);
  assign n71131 = (n70013 & n71129) | (n70013 & n71130) | (n71129 & n71130);
  assign n57678 = n33710 | n34208;
  assign n71132 = n57678 | n70995;
  assign n71133 = n57678 | n70994;
  assign n71134 = (n70013 & n71132) | (n70013 & n71133) | (n71132 & n71133);
  assign n34211 = ~n71131 & n71134;
  assign n34212 = x173 & x180;
  assign n34213 = n34211 & n34212;
  assign n34214 = n34211 | n34212;
  assign n34215 = ~n34213 & n34214;
  assign n57659 = n33717 | n33719;
  assign n57680 = n34215 & n57659;
  assign n57681 = n33717 & n34215;
  assign n71135 = (n57680 & n57681) | (n57680 & n70971) | (n57681 & n70971);
  assign n71136 = (n57680 & n57681) | (n57680 & n70970) | (n57681 & n70970);
  assign n71137 = (n70133 & n71135) | (n70133 & n71136) | (n71135 & n71136);
  assign n57683 = n34215 | n57659;
  assign n57684 = n33717 | n34215;
  assign n71138 = (n57683 & n57684) | (n57683 & n70971) | (n57684 & n70971);
  assign n71139 = (n57683 & n57684) | (n57683 & n70970) | (n57684 & n70970);
  assign n71140 = (n70133 & n71138) | (n70133 & n71139) | (n71138 & n71139);
  assign n34218 = ~n71137 & n71140;
  assign n34219 = x172 & x181;
  assign n34220 = n34218 & n34219;
  assign n34221 = n34218 | n34219;
  assign n34222 = ~n34220 & n34221;
  assign n71141 = n33724 | n33726;
  assign n71142 = (n33724 & n57405) | (n33724 & n71141) | (n57405 & n71141);
  assign n57686 = n34222 & n71142;
  assign n71143 = n33227 | n33724;
  assign n71144 = (n33724 & n33726) | (n33724 & n71143) | (n33726 & n71143);
  assign n57687 = n34222 & n71144;
  assign n57688 = (n70822 & n57686) | (n70822 & n57687) | (n57686 & n57687);
  assign n57689 = n34222 | n71142;
  assign n57690 = n34222 | n71144;
  assign n57691 = (n70822 & n57689) | (n70822 & n57690) | (n57689 & n57690);
  assign n34225 = ~n57688 & n57691;
  assign n34226 = x171 & x182;
  assign n34227 = n34225 & n34226;
  assign n34228 = n34225 | n34226;
  assign n34229 = ~n34227 & n34228;
  assign n57654 = n33731 | n33733;
  assign n57692 = n34229 & n57654;
  assign n57693 = n33731 & n34229;
  assign n71145 = (n57403 & n57692) | (n57403 & n57693) | (n57692 & n57693);
  assign n71146 = (n57402 & n57692) | (n57402 & n57693) | (n57692 & n57693);
  assign n71147 = (n70574 & n71145) | (n70574 & n71146) | (n71145 & n71146);
  assign n57695 = n34229 | n57654;
  assign n57696 = n33731 | n34229;
  assign n71148 = (n57403 & n57695) | (n57403 & n57696) | (n57695 & n57696);
  assign n71149 = (n57402 & n57695) | (n57402 & n57696) | (n57695 & n57696);
  assign n71150 = (n70574 & n71148) | (n70574 & n71149) | (n71148 & n71149);
  assign n34232 = ~n71147 & n71150;
  assign n34233 = x170 & x183;
  assign n34234 = n34232 & n34233;
  assign n34235 = n34232 | n34233;
  assign n34236 = ~n34234 & n34235;
  assign n71151 = n33738 | n33740;
  assign n71152 = (n33738 & n57400) | (n33738 & n71151) | (n57400 & n71151);
  assign n57698 = n34236 & n71152;
  assign n71153 = n33241 | n33738;
  assign n71154 = (n33738 & n33740) | (n33738 & n71153) | (n33740 & n71153);
  assign n57699 = n34236 & n71154;
  assign n57700 = (n57167 & n57698) | (n57167 & n57699) | (n57698 & n57699);
  assign n57701 = n34236 | n71152;
  assign n57702 = n34236 | n71154;
  assign n57703 = (n57167 & n57701) | (n57167 & n57702) | (n57701 & n57702);
  assign n34239 = ~n57700 & n57703;
  assign n34240 = x169 & x184;
  assign n34241 = n34239 & n34240;
  assign n34242 = n34239 | n34240;
  assign n34243 = ~n34241 & n34242;
  assign n71104 = n33745 | n33747;
  assign n71105 = (n33745 & n57398) | (n33745 & n71104) | (n57398 & n71104);
  assign n71155 = n34243 & n71105;
  assign n71106 = n33248 | n33745;
  assign n71107 = (n33745 & n33747) | (n33745 & n71106) | (n33747 & n71106);
  assign n71156 = n34243 & n71107;
  assign n71157 = (n70816 & n71155) | (n70816 & n71156) | (n71155 & n71156);
  assign n71158 = n34243 | n71105;
  assign n71159 = n34243 | n71107;
  assign n71160 = (n70816 & n71158) | (n70816 & n71159) | (n71158 & n71159);
  assign n34246 = ~n71157 & n71160;
  assign n34247 = x168 & x185;
  assign n34248 = n34246 & n34247;
  assign n34249 = n34246 | n34247;
  assign n34250 = ~n34248 & n34249;
  assign n57646 = n33752 | n33754;
  assign n57704 = n34250 & n57646;
  assign n57705 = n33752 & n34250;
  assign n71161 = (n57396 & n57704) | (n57396 & n57705) | (n57704 & n57705);
  assign n71162 = (n57704 & n57705) | (n57704 & n70966) | (n57705 & n70966);
  assign n71163 = (n70684 & n71161) | (n70684 & n71162) | (n71161 & n71162);
  assign n57707 = n34250 | n57646;
  assign n57708 = n33752 | n34250;
  assign n71164 = (n57396 & n57707) | (n57396 & n57708) | (n57707 & n57708);
  assign n71165 = (n57707 & n57708) | (n57707 & n70966) | (n57708 & n70966);
  assign n71166 = (n70684 & n71164) | (n70684 & n71165) | (n71164 & n71165);
  assign n34253 = ~n71163 & n71166;
  assign n34254 = x167 & x186;
  assign n34255 = n34253 & n34254;
  assign n34256 = n34253 | n34254;
  assign n34257 = ~n34255 & n34256;
  assign n34258 = n71103 & n34257;
  assign n34259 = n71103 | n34257;
  assign n34260 = ~n34258 & n34259;
  assign n34261 = x166 & x187;
  assign n34262 = n34260 & n34261;
  assign n34263 = n34260 | n34261;
  assign n34264 = ~n34262 & n34263;
  assign n57641 = n33766 | n33768;
  assign n57710 = n34264 & n57641;
  assign n57711 = n33766 & n34264;
  assign n57712 = (n70964 & n57710) | (n70964 & n57711) | (n57710 & n57711);
  assign n57713 = n34264 | n57641;
  assign n57714 = n33766 | n34264;
  assign n57715 = (n70964 & n57713) | (n70964 & n57714) | (n57713 & n57714);
  assign n34267 = ~n57712 & n57715;
  assign n34268 = x165 & x188;
  assign n34269 = n34267 & n34268;
  assign n34270 = n34267 | n34268;
  assign n34271 = ~n34269 & n34270;
  assign n57639 = n33773 | n57461;
  assign n71167 = n34271 & n57639;
  assign n71095 = n33276 | n33773;
  assign n71096 = (n33773 & n33775) | (n33773 & n71095) | (n33775 & n71095);
  assign n71168 = n34271 & n71096;
  assign n71169 = (n57154 & n71167) | (n57154 & n71168) | (n71167 & n71168);
  assign n71170 = n34271 | n57639;
  assign n71171 = n34271 | n71096;
  assign n71172 = (n57154 & n71170) | (n57154 & n71171) | (n71170 & n71171);
  assign n34274 = ~n71169 & n71172;
  assign n34275 = x164 & x189;
  assign n34276 = n34274 & n34275;
  assign n34277 = n34274 | n34275;
  assign n34278 = ~n34276 & n34277;
  assign n57716 = n33780 & n34278;
  assign n71173 = (n34278 & n57467) | (n34278 & n57716) | (n57467 & n57716);
  assign n71174 = (n34278 & n57468) | (n34278 & n57716) | (n57468 & n57716);
  assign n71175 = (n57151 & n71173) | (n57151 & n71174) | (n71173 & n71174);
  assign n57718 = n33780 | n34278;
  assign n71176 = n57467 | n57718;
  assign n71177 = n57468 | n57718;
  assign n71178 = (n57151 & n71176) | (n57151 & n71177) | (n71176 & n71177);
  assign n34281 = ~n71175 & n71178;
  assign n34282 = x163 & x190;
  assign n34283 = n34281 & n34282;
  assign n34284 = n34281 | n34282;
  assign n34285 = ~n34283 & n34284;
  assign n57636 = n33787 | n33789;
  assign n71179 = n34285 & n57636;
  assign n71093 = n33290 | n33787;
  assign n71094 = (n33787 & n33789) | (n33787 & n71093) | (n33789 & n71093);
  assign n71180 = n34285 & n71094;
  assign n71181 = (n57225 & n71179) | (n57225 & n71180) | (n71179 & n71180);
  assign n71182 = n34285 | n57636;
  assign n71183 = n34285 | n71094;
  assign n71184 = (n57225 & n71182) | (n57225 & n71183) | (n71182 & n71183);
  assign n34288 = ~n71181 & n71184;
  assign n34289 = x162 & x191;
  assign n34290 = n34288 & n34289;
  assign n34291 = n34288 | n34289;
  assign n34292 = ~n34290 & n34291;
  assign n57633 = n33794 | n33796;
  assign n57720 = n34292 & n57633;
  assign n57721 = n33794 & n34292;
  assign n57722 = (n70957 & n57720) | (n70957 & n57721) | (n57720 & n57721);
  assign n57723 = n34292 | n57633;
  assign n57724 = n33794 | n34292;
  assign n57725 = (n70957 & n57723) | (n70957 & n57724) | (n57723 & n57724);
  assign n34295 = ~n57722 & n57725;
  assign n34296 = x161 & x192;
  assign n34297 = n34295 & n34296;
  assign n34298 = n34295 | n34296;
  assign n34299 = ~n34297 & n34298;
  assign n57726 = n33801 & n34299;
  assign n71185 = (n34299 & n57478) | (n34299 & n57726) | (n57478 & n57726);
  assign n71186 = (n34299 & n57477) | (n34299 & n57726) | (n57477 & n57726);
  assign n71187 = (n57146 & n71185) | (n57146 & n71186) | (n71185 & n71186);
  assign n57728 = n33801 | n34299;
  assign n71188 = n57478 | n57728;
  assign n71189 = n57477 | n57728;
  assign n71190 = (n57146 & n71188) | (n57146 & n71189) | (n71188 & n71189);
  assign n34302 = ~n71187 & n71190;
  assign n34303 = x160 & x193;
  assign n34304 = n34302 & n34303;
  assign n34305 = n34302 | n34303;
  assign n34306 = ~n34304 & n34305;
  assign n57631 = n33808 | n33810;
  assign n71191 = n34306 & n57631;
  assign n71091 = n33311 | n33808;
  assign n71092 = (n33808 & n33810) | (n33808 & n71091) | (n33810 & n71091);
  assign n71192 = n34306 & n71092;
  assign n71193 = (n57235 & n71191) | (n57235 & n71192) | (n71191 & n71192);
  assign n71194 = n34306 | n57631;
  assign n71195 = n34306 | n71092;
  assign n71196 = (n57235 & n71194) | (n57235 & n71195) | (n71194 & n71195);
  assign n34309 = ~n71193 & n71196;
  assign n34310 = x159 & x194;
  assign n34311 = n34309 & n34310;
  assign n34312 = n34309 | n34310;
  assign n34313 = ~n34311 & n34312;
  assign n57628 = n33815 | n33817;
  assign n57730 = n34313 & n57628;
  assign n57731 = n33815 & n34313;
  assign n57732 = (n70952 & n57730) | (n70952 & n57731) | (n57730 & n57731);
  assign n57733 = n34313 | n57628;
  assign n57734 = n33815 | n34313;
  assign n57735 = (n70952 & n57733) | (n70952 & n57734) | (n57733 & n57734);
  assign n34316 = ~n57732 & n57735;
  assign n34317 = x158 & x195;
  assign n34318 = n34316 & n34317;
  assign n34319 = n34316 | n34317;
  assign n34320 = ~n34318 & n34319;
  assign n57736 = n33822 & n34320;
  assign n71197 = (n34320 & n57488) | (n34320 & n57736) | (n57488 & n57736);
  assign n71198 = (n34320 & n57487) | (n34320 & n57736) | (n57487 & n57736);
  assign n71199 = (n57141 & n71197) | (n57141 & n71198) | (n71197 & n71198);
  assign n57738 = n33822 | n34320;
  assign n71200 = n57488 | n57738;
  assign n71201 = n57487 | n57738;
  assign n71202 = (n57141 & n71200) | (n57141 & n71201) | (n71200 & n71201);
  assign n34323 = ~n71199 & n71202;
  assign n34324 = x157 & x196;
  assign n34325 = n34323 & n34324;
  assign n34326 = n34323 | n34324;
  assign n34327 = ~n34325 & n34326;
  assign n57626 = n33829 | n33831;
  assign n71203 = n34327 & n57626;
  assign n71089 = n33332 | n33829;
  assign n71090 = (n33829 & n33831) | (n33829 & n71089) | (n33831 & n71089);
  assign n71204 = n34327 & n71090;
  assign n71205 = (n57245 & n71203) | (n57245 & n71204) | (n71203 & n71204);
  assign n71206 = n34327 | n57626;
  assign n71207 = n34327 | n71090;
  assign n71208 = (n57245 & n71206) | (n57245 & n71207) | (n71206 & n71207);
  assign n34330 = ~n71205 & n71208;
  assign n34331 = x156 & x197;
  assign n34332 = n34330 & n34331;
  assign n34333 = n34330 | n34331;
  assign n34334 = ~n34332 & n34333;
  assign n57623 = n33836 | n33838;
  assign n57740 = n34334 & n57623;
  assign n57741 = n33836 & n34334;
  assign n57742 = (n70947 & n57740) | (n70947 & n57741) | (n57740 & n57741);
  assign n57743 = n34334 | n57623;
  assign n57744 = n33836 | n34334;
  assign n57745 = (n70947 & n57743) | (n70947 & n57744) | (n57743 & n57744);
  assign n34337 = ~n57742 & n57745;
  assign n34338 = x155 & x198;
  assign n34339 = n34337 & n34338;
  assign n34340 = n34337 | n34338;
  assign n34341 = ~n34339 & n34340;
  assign n57746 = n33843 & n34341;
  assign n71209 = (n34341 & n57498) | (n34341 & n57746) | (n57498 & n57746);
  assign n71210 = (n34341 & n57497) | (n34341 & n57746) | (n57497 & n57746);
  assign n71211 = (n70799 & n71209) | (n70799 & n71210) | (n71209 & n71210);
  assign n57748 = n33843 | n34341;
  assign n71212 = n57498 | n57748;
  assign n71213 = n57497 | n57748;
  assign n71214 = (n70799 & n71212) | (n70799 & n71213) | (n71212 & n71213);
  assign n34344 = ~n71211 & n71214;
  assign n34345 = x154 & x199;
  assign n34346 = n34344 & n34345;
  assign n34347 = n34344 | n34345;
  assign n34348 = ~n34346 & n34347;
  assign n34349 = n71088 & n34348;
  assign n34350 = n71088 | n34348;
  assign n34351 = ~n34349 & n34350;
  assign n34352 = x153 & x200;
  assign n34353 = n34351 & n34352;
  assign n34354 = n34351 | n34352;
  assign n34355 = ~n34353 & n34354;
  assign n57618 = n33857 | n33859;
  assign n57750 = n34355 & n57618;
  assign n57751 = n33857 & n34355;
  assign n57752 = (n70942 & n57750) | (n70942 & n57751) | (n57750 & n57751);
  assign n57753 = n34355 | n57618;
  assign n57754 = n33857 | n34355;
  assign n57755 = (n70942 & n57753) | (n70942 & n57754) | (n57753 & n57754);
  assign n34358 = ~n57752 & n57755;
  assign n34359 = x152 & x201;
  assign n34360 = n34358 & n34359;
  assign n34361 = n34358 | n34359;
  assign n34362 = ~n34360 & n34361;
  assign n57756 = n33864 & n34362;
  assign n71215 = (n34362 & n57508) | (n34362 & n57756) | (n57508 & n57756);
  assign n71216 = (n34362 & n57507) | (n34362 & n57756) | (n57507 & n57756);
  assign n71217 = (n70794 & n71215) | (n70794 & n71216) | (n71215 & n71216);
  assign n57758 = n33864 | n34362;
  assign n71218 = n57508 | n57758;
  assign n71219 = n57507 | n57758;
  assign n71220 = (n70794 & n71218) | (n70794 & n71219) | (n71218 & n71219);
  assign n34365 = ~n71217 & n71220;
  assign n34366 = x151 & x202;
  assign n34367 = n34365 & n34366;
  assign n34368 = n34365 | n34366;
  assign n34369 = ~n34367 & n34368;
  assign n34370 = n71083 & n34369;
  assign n34371 = n71083 | n34369;
  assign n34372 = ~n34370 & n34371;
  assign n34373 = x150 & x203;
  assign n34374 = n34372 & n34373;
  assign n34375 = n34372 | n34373;
  assign n34376 = ~n34374 & n34375;
  assign n57613 = n33878 | n33880;
  assign n57760 = n34376 & n57613;
  assign n57761 = n33878 & n34376;
  assign n57762 = (n57365 & n57760) | (n57365 & n57761) | (n57760 & n57761);
  assign n57763 = n34376 | n57613;
  assign n57764 = n33878 | n34376;
  assign n57765 = (n57365 & n57763) | (n57365 & n57764) | (n57763 & n57764);
  assign n34379 = ~n57762 & n57765;
  assign n34380 = x149 & x204;
  assign n34381 = n34379 & n34380;
  assign n34382 = n34379 | n34380;
  assign n34383 = ~n34381 & n34382;
  assign n57766 = n33885 & n34383;
  assign n57767 = (n34383 & n71059) | (n34383 & n57766) | (n71059 & n57766);
  assign n57768 = n33885 | n34383;
  assign n57769 = n71059 | n57768;
  assign n34386 = ~n57767 & n57769;
  assign n34387 = x148 & x205;
  assign n34388 = n34386 & n34387;
  assign n34389 = n34386 | n34387;
  assign n34390 = ~n34388 & n34389;
  assign n57770 = n33892 & n34390;
  assign n57771 = (n34390 & n57522) | (n34390 & n57770) | (n57522 & n57770);
  assign n57772 = n33892 | n34390;
  assign n57773 = n57522 | n57772;
  assign n34393 = ~n57771 & n57773;
  assign n34394 = x147 & x206;
  assign n34395 = n34393 & n34394;
  assign n34396 = n34393 | n34394;
  assign n34397 = ~n34395 & n34396;
  assign n57774 = n33899 & n34397;
  assign n57775 = (n34397 & n57526) | (n34397 & n57774) | (n57526 & n57774);
  assign n57776 = n33899 | n34397;
  assign n57777 = n57526 | n57776;
  assign n34400 = ~n57775 & n57777;
  assign n34401 = x146 & x207;
  assign n34402 = n34400 & n34401;
  assign n34403 = n34400 | n34401;
  assign n34404 = ~n34402 & n34403;
  assign n57778 = n33906 & n34404;
  assign n57779 = (n34404 & n57530) | (n34404 & n57778) | (n57530 & n57778);
  assign n57780 = n33906 | n34404;
  assign n57781 = n57530 | n57780;
  assign n34407 = ~n57779 & n57781;
  assign n34408 = x145 & x208;
  assign n34409 = n34407 & n34408;
  assign n34410 = n34407 | n34408;
  assign n34411 = ~n34409 & n34410;
  assign n57782 = n33913 & n34411;
  assign n57783 = (n34411 & n57534) | (n34411 & n57782) | (n57534 & n57782);
  assign n57784 = n33913 | n34411;
  assign n57785 = n57534 | n57784;
  assign n34414 = ~n57783 & n57785;
  assign n34415 = x144 & x209;
  assign n34416 = n34414 & n34415;
  assign n34417 = n34414 | n34415;
  assign n34418 = ~n34416 & n34417;
  assign n57786 = n33920 & n34418;
  assign n57787 = (n34418 & n57538) | (n34418 & n57786) | (n57538 & n57786);
  assign n57788 = n33920 | n34418;
  assign n57789 = n57538 | n57788;
  assign n34421 = ~n57787 & n57789;
  assign n34422 = x143 & x210;
  assign n34423 = n34421 & n34422;
  assign n34424 = n34421 | n34422;
  assign n34425 = ~n34423 & n34424;
  assign n57790 = n33927 & n34425;
  assign n57791 = (n34425 & n57542) | (n34425 & n57790) | (n57542 & n57790);
  assign n57792 = n33927 | n34425;
  assign n57793 = n57542 | n57792;
  assign n34428 = ~n57791 & n57793;
  assign n34429 = x142 & x211;
  assign n34430 = n34428 & n34429;
  assign n34431 = n34428 | n34429;
  assign n34432 = ~n34430 & n34431;
  assign n57794 = n33934 & n34432;
  assign n57795 = (n34432 & n57546) | (n34432 & n57794) | (n57546 & n57794);
  assign n57796 = n33934 | n34432;
  assign n57797 = n57546 | n57796;
  assign n34435 = ~n57795 & n57797;
  assign n34436 = x141 & x212;
  assign n34437 = n34435 & n34436;
  assign n34438 = n34435 | n34436;
  assign n34439 = ~n34437 & n34438;
  assign n57798 = n33941 & n34439;
  assign n57799 = (n34439 & n57550) | (n34439 & n57798) | (n57550 & n57798);
  assign n57800 = n33941 | n34439;
  assign n57801 = n57550 | n57800;
  assign n34442 = ~n57799 & n57801;
  assign n34443 = x140 & x213;
  assign n34444 = n34442 & n34443;
  assign n34445 = n34442 | n34443;
  assign n34446 = ~n34444 & n34445;
  assign n57802 = n33948 & n34446;
  assign n57803 = (n34446 & n57554) | (n34446 & n57802) | (n57554 & n57802);
  assign n57804 = n33948 | n34446;
  assign n57805 = n57554 | n57804;
  assign n34449 = ~n57803 & n57805;
  assign n34450 = x139 & x214;
  assign n34451 = n34449 & n34450;
  assign n34452 = n34449 | n34450;
  assign n34453 = ~n34451 & n34452;
  assign n57806 = n33955 & n34453;
  assign n57807 = (n34453 & n57558) | (n34453 & n57806) | (n57558 & n57806);
  assign n57808 = n33955 | n34453;
  assign n57809 = n57558 | n57808;
  assign n34456 = ~n57807 & n57809;
  assign n34457 = x138 & x215;
  assign n34458 = n34456 & n34457;
  assign n34459 = n34456 | n34457;
  assign n34460 = ~n34458 & n34459;
  assign n57810 = n33962 & n34460;
  assign n57811 = (n34460 & n57562) | (n34460 & n57810) | (n57562 & n57810);
  assign n57812 = n33962 | n34460;
  assign n57813 = n57562 | n57812;
  assign n34463 = ~n57811 & n57813;
  assign n34464 = x137 & x216;
  assign n34465 = n34463 & n34464;
  assign n34466 = n34463 | n34464;
  assign n34467 = ~n34465 & n34466;
  assign n57814 = n33969 & n34467;
  assign n57815 = (n34467 & n57566) | (n34467 & n57814) | (n57566 & n57814);
  assign n57816 = n33969 | n34467;
  assign n57817 = n57566 | n57816;
  assign n34470 = ~n57815 & n57817;
  assign n34471 = x136 & x217;
  assign n34472 = n34470 & n34471;
  assign n34473 = n34470 | n34471;
  assign n34474 = ~n34472 & n34473;
  assign n57818 = n33976 & n34474;
  assign n57819 = (n34474 & n57570) | (n34474 & n57818) | (n57570 & n57818);
  assign n57820 = n33976 | n34474;
  assign n57821 = n57570 | n57820;
  assign n34477 = ~n57819 & n57821;
  assign n34478 = x135 & x218;
  assign n34479 = n34477 & n34478;
  assign n34480 = n34477 | n34478;
  assign n34481 = ~n34479 & n34480;
  assign n57822 = n33983 & n34481;
  assign n57823 = (n34481 & n57574) | (n34481 & n57822) | (n57574 & n57822);
  assign n57824 = n33983 | n34481;
  assign n57825 = n57574 | n57824;
  assign n34484 = ~n57823 & n57825;
  assign n34485 = x134 & x219;
  assign n34486 = n34484 & n34485;
  assign n34487 = n34484 | n34485;
  assign n34488 = ~n34486 & n34487;
  assign n57826 = n33990 & n34488;
  assign n57827 = (n34488 & n57578) | (n34488 & n57826) | (n57578 & n57826);
  assign n57828 = n33990 | n34488;
  assign n57829 = n57578 | n57828;
  assign n34491 = ~n57827 & n57829;
  assign n34492 = x133 & x220;
  assign n34493 = n34491 & n34492;
  assign n34494 = n34491 | n34492;
  assign n34495 = ~n34493 & n34494;
  assign n57830 = n33997 & n34495;
  assign n57831 = (n34495 & n57582) | (n34495 & n57830) | (n57582 & n57830);
  assign n57832 = n33997 | n34495;
  assign n57833 = n57582 | n57832;
  assign n34498 = ~n57831 & n57833;
  assign n34499 = x132 & x221;
  assign n34500 = n34498 & n34499;
  assign n34501 = n34498 | n34499;
  assign n34502 = ~n34500 & n34501;
  assign n57834 = n34004 & n34502;
  assign n57835 = (n34502 & n57586) | (n34502 & n57834) | (n57586 & n57834);
  assign n57836 = n34004 | n34502;
  assign n57837 = n57586 | n57836;
  assign n34505 = ~n57835 & n57837;
  assign n34506 = x131 & x222;
  assign n34507 = n34505 & n34506;
  assign n34508 = n34505 | n34506;
  assign n34509 = ~n34507 & n34508;
  assign n57838 = n34011 & n34509;
  assign n57839 = (n34509 & n57590) | (n34509 & n57838) | (n57590 & n57838);
  assign n57840 = n34011 | n34509;
  assign n57841 = n57590 | n57840;
  assign n34512 = ~n57839 & n57841;
  assign n34513 = x130 & x223;
  assign n34514 = n34512 & n34513;
  assign n34515 = n34512 | n34513;
  assign n34516 = ~n34514 & n34515;
  assign n57842 = n34018 & n34516;
  assign n57843 = (n34516 & n57595) | (n34516 & n57842) | (n57595 & n57842);
  assign n57844 = n34018 | n34516;
  assign n57845 = n57595 | n57844;
  assign n34519 = ~n57843 & n57845;
  assign n34520 = x129 & x224;
  assign n34521 = n34519 & n34520;
  assign n34522 = n34519 | n34520;
  assign n34523 = ~n34521 & n34522;
  assign n57611 = n34025 | n34027;
  assign n57846 = n34523 & n57611;
  assign n57847 = n34025 & n34523;
  assign n57848 = (n57360 & n57846) | (n57360 & n57847) | (n57846 & n57847);
  assign n57849 = n34523 | n57611;
  assign n57850 = n34025 | n34523;
  assign n57851 = (n57360 & n57849) | (n57360 & n57850) | (n57849 & n57850);
  assign n34526 = ~n57848 & n57851;
  assign n34527 = x128 & x225;
  assign n34528 = n34526 & n34527;
  assign n34529 = n34526 | n34527;
  assign n34530 = ~n34528 & n34529;
  assign n57609 = n34032 | n34034;
  assign n71221 = n34530 & n57609;
  assign n71222 = n34032 & n34530;
  assign n71223 = (n57358 & n71221) | (n57358 & n71222) | (n71221 & n71222);
  assign n71224 = n34530 | n57609;
  assign n71225 = n34032 | n34530;
  assign n71226 = (n57358 & n71224) | (n57358 & n71225) | (n71224 & n71225);
  assign n34533 = ~n71223 & n71226;
  assign n34534 = x127 & x226;
  assign n34535 = n34533 & n34534;
  assign n34536 = n34533 | n34534;
  assign n34537 = ~n34535 & n34536;
  assign n57607 = n34039 | n34041;
  assign n71227 = n34537 & n57607;
  assign n71228 = n34039 & n34537;
  assign n71229 = (n57356 & n71227) | (n57356 & n71228) | (n71227 & n71228);
  assign n71230 = n34537 | n57607;
  assign n71231 = n34039 | n34537;
  assign n71232 = (n57356 & n71230) | (n57356 & n71231) | (n71230 & n71231);
  assign n34540 = ~n71229 & n71232;
  assign n34541 = x126 & x227;
  assign n34542 = n34540 & n34541;
  assign n34543 = n34540 | n34541;
  assign n34544 = ~n34542 & n34543;
  assign n34545 = n57606 & n34544;
  assign n34546 = n57606 | n34544;
  assign n34547 = ~n34545 & n34546;
  assign n34548 = x125 & x228;
  assign n34549 = n34547 & n34548;
  assign n34550 = n34547 | n34548;
  assign n34551 = ~n34549 & n34550;
  assign n34552 = n57604 & n34551;
  assign n34553 = n57604 | n34551;
  assign n34554 = ~n34552 & n34553;
  assign n34555 = x124 & x229;
  assign n34556 = n34554 & n34555;
  assign n34557 = n34554 | n34555;
  assign n34558 = ~n34556 & n34557;
  assign n34559 = n34146 & n34558;
  assign n34560 = n34146 | n34558;
  assign n34561 = ~n34559 & n34560;
  assign n34562 = x123 & x230;
  assign n34563 = n34561 & n34562;
  assign n34564 = n34561 | n34562;
  assign n34565 = ~n34563 & n34564;
  assign n34566 = n34145 & n34565;
  assign n34567 = n34145 | n34565;
  assign n34568 = ~n34566 & n34567;
  assign n34569 = x122 & x231;
  assign n34570 = n34568 & n34569;
  assign n34571 = n34568 | n34569;
  assign n34572 = ~n34570 & n34571;
  assign n34573 = n34144 & n34572;
  assign n34574 = n34144 | n34572;
  assign n34575 = ~n34573 & n34574;
  assign n34576 = x121 & x232;
  assign n34577 = n34575 & n34576;
  assign n34578 = n34575 | n34576;
  assign n34579 = ~n34577 & n34578;
  assign n34580 = n34143 & n34579;
  assign n34581 = n34143 | n34579;
  assign n34582 = ~n34580 & n34581;
  assign n34583 = x120 & x233;
  assign n34584 = n34582 & n34583;
  assign n34585 = n34582 | n34583;
  assign n34586 = ~n34584 & n34585;
  assign n34587 = n34142 & n34586;
  assign n34588 = n34142 | n34586;
  assign n34589 = ~n34587 & n34588;
  assign n34590 = x119 & x234;
  assign n34591 = n34589 & n34590;
  assign n34592 = n34589 | n34590;
  assign n34593 = ~n34591 & n34592;
  assign n34594 = n34141 & n34593;
  assign n34595 = n34141 | n34593;
  assign n34596 = ~n34594 & n34595;
  assign n34597 = x118 & x235;
  assign n34598 = n34596 & n34597;
  assign n34599 = n34596 | n34597;
  assign n34600 = ~n34598 & n34599;
  assign n34601 = n34140 & n34600;
  assign n34602 = n34140 | n34600;
  assign n34603 = ~n34601 & n34602;
  assign n34604 = x117 & x236;
  assign n34605 = n34603 & n34604;
  assign n34606 = n34603 | n34604;
  assign n34607 = ~n34605 & n34606;
  assign n34608 = n34139 & n34607;
  assign n34609 = n34139 | n34607;
  assign n34610 = ~n34608 & n34609;
  assign n34611 = x116 & x237;
  assign n34612 = n34610 & n34611;
  assign n34613 = n34610 | n34611;
  assign n34614 = ~n34612 & n34613;
  assign n34615 = n71078 & n34614;
  assign n34616 = n71078 | n34614;
  assign n34617 = ~n34615 & n34616;
  assign n34618 = x115 & x238;
  assign n34619 = n34617 & n34618;
  assign n34620 = n34617 | n34618;
  assign n34621 = ~n34619 & n34620;
  assign n34622 = n57602 & n34621;
  assign n34623 = n57602 | n34621;
  assign n34624 = ~n34622 & n34623;
  assign n34625 = x114 & x239;
  assign n34626 = n34624 & n34625;
  assign n34627 = n34624 | n34625;
  assign n34628 = ~n34626 & n34627;
  assign n34629 = n57600 & n34628;
  assign n34630 = n57600 | n34628;
  assign n34631 = ~n34629 & n34630;
  assign n57852 = n34626 | n57600;
  assign n57853 = (n34626 & n34628) | (n34626 & n57852) | (n34628 & n57852);
  assign n57854 = n34619 | n57602;
  assign n57855 = (n34619 & n34621) | (n34619 & n57854) | (n34621 & n57854);
  assign n71233 = n34612 | n71078;
  assign n71234 = (n34612 & n34614) | (n34612 & n71233) | (n34614 & n71233);
  assign n34635 = n34605 | n34608;
  assign n34636 = n34598 | n34601;
  assign n34637 = n34591 | n34594;
  assign n34638 = n34584 | n34587;
  assign n34639 = n34577 | n34580;
  assign n34640 = n34570 | n34573;
  assign n34641 = n34563 | n34566;
  assign n57856 = n34556 | n34558;
  assign n57857 = (n34146 & n34556) | (n34146 & n57856) | (n34556 & n57856);
  assign n57858 = n34549 | n34551;
  assign n57859 = (n34549 & n57604) | (n34549 & n57858) | (n57604 & n57858);
  assign n57608 = (n34039 & n57356) | (n34039 & n57607) | (n57356 & n57607);
  assign n57610 = (n34032 & n57358) | (n34032 & n57609) | (n57358 & n57609);
  assign n57872 = n34360 | n34362;
  assign n71237 = n33864 | n34360;
  assign n71238 = (n34360 & n34362) | (n34360 & n71237) | (n34362 & n71237);
  assign n71239 = (n57508 & n57872) | (n57508 & n71238) | (n57872 & n71238);
  assign n71240 = (n57507 & n57872) | (n57507 & n71238) | (n57872 & n71238);
  assign n71241 = (n70794 & n71239) | (n70794 & n71240) | (n71239 & n71240);
  assign n57877 = n34339 | n34341;
  assign n71242 = n33843 | n34339;
  assign n71243 = (n34339 & n34341) | (n34339 & n71242) | (n34341 & n71242);
  assign n71244 = (n57498 & n57877) | (n57498 & n71243) | (n57877 & n71243);
  assign n71245 = (n57497 & n57877) | (n57497 & n71243) | (n57877 & n71243);
  assign n71246 = (n70799 & n71244) | (n70799 & n71245) | (n71244 & n71245);
  assign n57627 = (n57245 & n71090) | (n57245 & n57626) | (n71090 & n57626);
  assign n57882 = n34318 | n34320;
  assign n71247 = n33822 | n34318;
  assign n71248 = (n34318 & n34320) | (n34318 & n71247) | (n34320 & n71247);
  assign n71249 = (n57488 & n57882) | (n57488 & n71248) | (n57882 & n71248);
  assign n71250 = (n57487 & n57882) | (n57487 & n71248) | (n57882 & n71248);
  assign n71251 = (n57141 & n71249) | (n57141 & n71250) | (n71249 & n71250);
  assign n57632 = (n57235 & n71092) | (n57235 & n57631) | (n71092 & n57631);
  assign n57887 = n34297 | n34299;
  assign n71252 = n33801 | n34297;
  assign n71253 = (n34297 & n34299) | (n34297 & n71252) | (n34299 & n71252);
  assign n71254 = (n57478 & n57887) | (n57478 & n71253) | (n57887 & n71253);
  assign n71255 = (n57477 & n57887) | (n57477 & n71253) | (n57887 & n71253);
  assign n71256 = (n57146 & n71254) | (n57146 & n71255) | (n71254 & n71255);
  assign n57637 = (n57225 & n71094) | (n57225 & n57636) | (n71094 & n57636);
  assign n57892 = n34276 | n34278;
  assign n71257 = n33780 | n34276;
  assign n71258 = (n34276 & n34278) | (n34276 & n71257) | (n34278 & n71257);
  assign n71259 = (n57467 & n57892) | (n57467 & n71258) | (n57892 & n71258);
  assign n71260 = (n57468 & n57892) | (n57468 & n71258) | (n57892 & n71258);
  assign n71261 = (n57151 & n71259) | (n57151 & n71260) | (n71259 & n71260);
  assign n71264 = n33752 | n34248;
  assign n71265 = (n34248 & n34250) | (n34248 & n71264) | (n34250 & n71264);
  assign n71266 = n34248 | n34250;
  assign n71267 = (n34248 & n57646) | (n34248 & n71266) | (n57646 & n71266);
  assign n71268 = (n57396 & n71265) | (n57396 & n71267) | (n71265 & n71267);
  assign n71269 = (n70966 & n71265) | (n70966 & n71267) | (n71265 & n71267);
  assign n71270 = (n70684 & n71268) | (n70684 & n71269) | (n71268 & n71269);
  assign n34694 = x175 & x179;
  assign n71274 = n34694 & n57665;
  assign n71275 = n34694 & n71109;
  assign n71276 = (n70695 & n71274) | (n70695 & n71275) | (n71274 & n71275);
  assign n71277 = (n34694 & n71120) | (n34694 & n71276) | (n71120 & n71276);
  assign n71278 = (n34694 & n71119) | (n34694 & n71276) | (n71119 & n71276);
  assign n71279 = (n69887 & n71277) | (n69887 & n71278) | (n71277 & n71278);
  assign n71280 = n34694 | n57665;
  assign n71281 = n34694 | n71109;
  assign n71282 = (n70695 & n71280) | (n70695 & n71281) | (n71280 & n71281);
  assign n71283 = n71120 | n71282;
  assign n71284 = n71119 | n71282;
  assign n71285 = (n69887 & n71283) | (n69887 & n71284) | (n71283 & n71284);
  assign n34697 = ~n71279 & n71285;
  assign n71286 = n33710 | n34206;
  assign n71287 = (n34206 & n34208) | (n34206 & n71286) | (n34208 & n71286);
  assign n57922 = n34697 & n71287;
  assign n71288 = n34206 & n34697;
  assign n71289 = (n34208 & n34697) | (n34208 & n71288) | (n34697 & n71288);
  assign n71290 = (n57922 & n70995) | (n57922 & n71289) | (n70995 & n71289);
  assign n71291 = (n57922 & n70994) | (n57922 & n71289) | (n70994 & n71289);
  assign n71292 = (n70013 & n71290) | (n70013 & n71291) | (n71290 & n71291);
  assign n57925 = n34697 | n71287;
  assign n71293 = n34206 | n34697;
  assign n71294 = n34208 | n71293;
  assign n71295 = (n57925 & n70995) | (n57925 & n71294) | (n70995 & n71294);
  assign n71296 = (n57925 & n70994) | (n57925 & n71294) | (n70994 & n71294);
  assign n71297 = (n70013 & n71295) | (n70013 & n71296) | (n71295 & n71296);
  assign n34700 = ~n71292 & n71297;
  assign n34701 = x174 & x180;
  assign n34702 = n34700 & n34701;
  assign n34703 = n34700 | n34701;
  assign n34704 = ~n34702 & n34703;
  assign n71298 = n34213 | n34215;
  assign n71299 = (n34213 & n57659) | (n34213 & n71298) | (n57659 & n71298);
  assign n57928 = n34704 & n71299;
  assign n71300 = n33717 | n34213;
  assign n71301 = (n34213 & n34215) | (n34213 & n71300) | (n34215 & n71300);
  assign n57929 = n34704 & n71301;
  assign n71302 = (n57928 & n57929) | (n57928 & n70971) | (n57929 & n70971);
  assign n71303 = (n57928 & n57929) | (n57928 & n70970) | (n57929 & n70970);
  assign n71304 = (n70133 & n71302) | (n70133 & n71303) | (n71302 & n71303);
  assign n57931 = n34704 | n71299;
  assign n57932 = n34704 | n71301;
  assign n71305 = (n57931 & n57932) | (n57931 & n70971) | (n57932 & n70971);
  assign n71306 = (n57931 & n57932) | (n57931 & n70970) | (n57932 & n70970);
  assign n71307 = (n70133 & n71305) | (n70133 & n71306) | (n71305 & n71306);
  assign n34707 = ~n71304 & n71307;
  assign n34708 = x173 & x181;
  assign n34709 = n34707 & n34708;
  assign n34710 = n34707 | n34708;
  assign n34711 = ~n34709 & n34710;
  assign n71271 = n34220 | n34222;
  assign n71273 = (n34220 & n71142) | (n34220 & n71271) | (n71142 & n71271);
  assign n71308 = n34711 & n71273;
  assign n71272 = (n34220 & n71144) | (n34220 & n71271) | (n71144 & n71271);
  assign n71309 = n34711 & n71272;
  assign n71310 = (n70822 & n71308) | (n70822 & n71309) | (n71308 & n71309);
  assign n71311 = n34711 | n71273;
  assign n71312 = n34711 | n71272;
  assign n71313 = (n70822 & n71311) | (n70822 & n71312) | (n71311 & n71312);
  assign n34714 = ~n71310 & n71313;
  assign n34715 = x172 & x182;
  assign n34716 = n34714 & n34715;
  assign n34717 = n34714 | n34715;
  assign n34718 = ~n34716 & n34717;
  assign n71314 = n34227 | n34229;
  assign n71315 = (n34227 & n57654) | (n34227 & n71314) | (n57654 & n71314);
  assign n57934 = n34718 & n71315;
  assign n71316 = n33731 | n34227;
  assign n71317 = (n34227 & n34229) | (n34227 & n71316) | (n34229 & n71316);
  assign n57935 = n34718 & n71317;
  assign n71318 = (n57403 & n57934) | (n57403 & n57935) | (n57934 & n57935);
  assign n71319 = (n57402 & n57934) | (n57402 & n57935) | (n57934 & n57935);
  assign n71320 = (n70574 & n71318) | (n70574 & n71319) | (n71318 & n71319);
  assign n57937 = n34718 | n71315;
  assign n57938 = n34718 | n71317;
  assign n71321 = (n57403 & n57937) | (n57403 & n57938) | (n57937 & n57938);
  assign n71322 = (n57402 & n57937) | (n57402 & n57938) | (n57937 & n57938);
  assign n71323 = (n70574 & n71321) | (n70574 & n71322) | (n71321 & n71322);
  assign n34721 = ~n71320 & n71323;
  assign n34722 = x171 & x183;
  assign n34723 = n34721 & n34722;
  assign n34724 = n34721 | n34722;
  assign n34725 = ~n34723 & n34724;
  assign n57940 = n34234 & n34725;
  assign n71324 = (n34725 & n57698) | (n34725 & n57940) | (n57698 & n57940);
  assign n71325 = (n34725 & n57699) | (n34725 & n57940) | (n57699 & n57940);
  assign n71326 = (n57167 & n71324) | (n57167 & n71325) | (n71324 & n71325);
  assign n57942 = n34234 | n34725;
  assign n71327 = n57698 | n57942;
  assign n71328 = n57699 | n57942;
  assign n71329 = (n57167 & n71327) | (n57167 & n71328) | (n71327 & n71328);
  assign n34728 = ~n71326 & n71329;
  assign n34729 = x170 & x184;
  assign n34730 = n34728 & n34729;
  assign n34731 = n34728 | n34729;
  assign n34732 = ~n34730 & n34731;
  assign n57904 = n34241 | n34243;
  assign n57944 = n34732 & n57904;
  assign n57945 = n34241 & n34732;
  assign n71330 = (n57944 & n57945) | (n57944 & n71105) | (n57945 & n71105);
  assign n71331 = (n57944 & n57945) | (n57944 & n71107) | (n57945 & n71107);
  assign n71332 = (n70816 & n71330) | (n70816 & n71331) | (n71330 & n71331);
  assign n57947 = n34732 | n57904;
  assign n57948 = n34241 | n34732;
  assign n71333 = (n57947 & n57948) | (n57947 & n71105) | (n57948 & n71105);
  assign n71334 = (n57947 & n57948) | (n57947 & n71107) | (n57948 & n71107);
  assign n71335 = (n70816 & n71333) | (n70816 & n71334) | (n71333 & n71334);
  assign n34735 = ~n71332 & n71335;
  assign n34736 = x169 & x185;
  assign n34737 = n34735 & n34736;
  assign n34738 = n34735 | n34736;
  assign n34739 = ~n34737 & n34738;
  assign n34740 = n71270 & n34739;
  assign n34741 = n71270 | n34739;
  assign n34742 = ~n34740 & n34741;
  assign n34743 = x168 & x186;
  assign n34744 = n34742 & n34743;
  assign n34745 = n34742 | n34743;
  assign n34746 = ~n34744 & n34745;
  assign n57899 = n34255 | n34257;
  assign n57950 = n34746 & n57899;
  assign n57951 = n34255 & n34746;
  assign n57952 = (n71103 & n57950) | (n71103 & n57951) | (n57950 & n57951);
  assign n57953 = n34746 | n57899;
  assign n57954 = n34255 | n34746;
  assign n57955 = (n71103 & n57953) | (n71103 & n57954) | (n57953 & n57954);
  assign n34749 = ~n57952 & n57955;
  assign n34750 = x167 & x187;
  assign n34751 = n34749 & n34750;
  assign n34752 = n34749 | n34750;
  assign n34753 = ~n34751 & n34752;
  assign n57897 = n34262 | n57710;
  assign n71336 = n34753 & n57897;
  assign n71262 = n33766 | n34262;
  assign n71263 = (n34262 & n34264) | (n34262 & n71262) | (n34264 & n71262);
  assign n71337 = n34753 & n71263;
  assign n71338 = (n70964 & n71336) | (n70964 & n71337) | (n71336 & n71337);
  assign n71339 = n34753 | n57897;
  assign n71340 = n34753 | n71263;
  assign n71341 = (n70964 & n71339) | (n70964 & n71340) | (n71339 & n71340);
  assign n34756 = ~n71338 & n71341;
  assign n34757 = x166 & x188;
  assign n34758 = n34756 & n34757;
  assign n34759 = n34756 | n34757;
  assign n34760 = ~n34758 & n34759;
  assign n57894 = n34269 | n34271;
  assign n57956 = n34760 & n57894;
  assign n57957 = n34269 & n34760;
  assign n71342 = (n57639 & n57956) | (n57639 & n57957) | (n57956 & n57957);
  assign n71343 = (n57956 & n57957) | (n57956 & n71096) | (n57957 & n71096);
  assign n71344 = (n57154 & n71342) | (n57154 & n71343) | (n71342 & n71343);
  assign n57959 = n34760 | n57894;
  assign n57960 = n34269 | n34760;
  assign n71345 = (n57639 & n57959) | (n57639 & n57960) | (n57959 & n57960);
  assign n71346 = (n57959 & n57960) | (n57959 & n71096) | (n57960 & n71096);
  assign n71347 = (n57154 & n71345) | (n57154 & n71346) | (n71345 & n71346);
  assign n34763 = ~n71344 & n71347;
  assign n34764 = x165 & x189;
  assign n34765 = n34763 & n34764;
  assign n34766 = n34763 | n34764;
  assign n34767 = ~n34765 & n34766;
  assign n34768 = n71261 & n34767;
  assign n34769 = n71261 | n34767;
  assign n34770 = ~n34768 & n34769;
  assign n34771 = x164 & x190;
  assign n34772 = n34770 & n34771;
  assign n34773 = n34770 | n34771;
  assign n34774 = ~n34772 & n34773;
  assign n57889 = n34283 | n34285;
  assign n57962 = n34774 & n57889;
  assign n57963 = n34283 & n34774;
  assign n57964 = (n57637 & n57962) | (n57637 & n57963) | (n57962 & n57963);
  assign n57965 = n34774 | n57889;
  assign n57966 = n34283 | n34774;
  assign n57967 = (n57637 & n57965) | (n57637 & n57966) | (n57965 & n57966);
  assign n34777 = ~n57964 & n57967;
  assign n34778 = x163 & x191;
  assign n34779 = n34777 & n34778;
  assign n34780 = n34777 | n34778;
  assign n34781 = ~n34779 & n34780;
  assign n57968 = n34290 & n34781;
  assign n57969 = (n34781 & n57722) | (n34781 & n57968) | (n57722 & n57968);
  assign n57970 = n34290 | n34781;
  assign n57971 = n57722 | n57970;
  assign n34784 = ~n57969 & n57971;
  assign n34785 = x162 & x192;
  assign n34786 = n34784 & n34785;
  assign n34787 = n34784 | n34785;
  assign n34788 = ~n34786 & n34787;
  assign n34789 = n71256 & n34788;
  assign n34790 = n71256 | n34788;
  assign n34791 = ~n34789 & n34790;
  assign n34792 = x161 & x193;
  assign n34793 = n34791 & n34792;
  assign n34794 = n34791 | n34792;
  assign n34795 = ~n34793 & n34794;
  assign n57884 = n34304 | n34306;
  assign n57972 = n34795 & n57884;
  assign n57973 = n34304 & n34795;
  assign n57974 = (n57632 & n57972) | (n57632 & n57973) | (n57972 & n57973);
  assign n57975 = n34795 | n57884;
  assign n57976 = n34304 | n34795;
  assign n57977 = (n57632 & n57975) | (n57632 & n57976) | (n57975 & n57976);
  assign n34798 = ~n57974 & n57977;
  assign n34799 = x160 & x194;
  assign n34800 = n34798 & n34799;
  assign n34801 = n34798 | n34799;
  assign n34802 = ~n34800 & n34801;
  assign n57978 = n34311 & n34802;
  assign n57979 = (n34802 & n57732) | (n34802 & n57978) | (n57732 & n57978);
  assign n57980 = n34311 | n34802;
  assign n57981 = n57732 | n57980;
  assign n34805 = ~n57979 & n57981;
  assign n34806 = x159 & x195;
  assign n34807 = n34805 & n34806;
  assign n34808 = n34805 | n34806;
  assign n34809 = ~n34807 & n34808;
  assign n34810 = n71251 & n34809;
  assign n34811 = n71251 | n34809;
  assign n34812 = ~n34810 & n34811;
  assign n34813 = x158 & x196;
  assign n34814 = n34812 & n34813;
  assign n34815 = n34812 | n34813;
  assign n34816 = ~n34814 & n34815;
  assign n57879 = n34325 | n34327;
  assign n57982 = n34816 & n57879;
  assign n57983 = n34325 & n34816;
  assign n57984 = (n57627 & n57982) | (n57627 & n57983) | (n57982 & n57983);
  assign n57985 = n34816 | n57879;
  assign n57986 = n34325 | n34816;
  assign n57987 = (n57627 & n57985) | (n57627 & n57986) | (n57985 & n57986);
  assign n34819 = ~n57984 & n57987;
  assign n34820 = x157 & x197;
  assign n34821 = n34819 & n34820;
  assign n34822 = n34819 | n34820;
  assign n34823 = ~n34821 & n34822;
  assign n57988 = n34332 & n34823;
  assign n57989 = (n34823 & n57742) | (n34823 & n57988) | (n57742 & n57988);
  assign n57990 = n34332 | n34823;
  assign n57991 = n57742 | n57990;
  assign n34826 = ~n57989 & n57991;
  assign n34827 = x156 & x198;
  assign n34828 = n34826 & n34827;
  assign n34829 = n34826 | n34827;
  assign n34830 = ~n34828 & n34829;
  assign n34831 = n71246 & n34830;
  assign n34832 = n71246 | n34830;
  assign n34833 = ~n34831 & n34832;
  assign n34834 = x155 & x199;
  assign n34835 = n34833 & n34834;
  assign n34836 = n34833 | n34834;
  assign n34837 = ~n34835 & n34836;
  assign n57874 = n34346 | n34348;
  assign n57992 = n34837 & n57874;
  assign n57993 = n34346 & n34837;
  assign n57994 = (n71088 & n57992) | (n71088 & n57993) | (n57992 & n57993);
  assign n57995 = n34837 | n57874;
  assign n57996 = n34346 | n34837;
  assign n57997 = (n71088 & n57995) | (n71088 & n57996) | (n57995 & n57996);
  assign n34840 = ~n57994 & n57997;
  assign n34841 = x154 & x200;
  assign n34842 = n34840 & n34841;
  assign n34843 = n34840 | n34841;
  assign n34844 = ~n34842 & n34843;
  assign n57998 = n34353 & n34844;
  assign n71348 = (n34844 & n57751) | (n34844 & n57998) | (n57751 & n57998);
  assign n71349 = (n34844 & n57750) | (n34844 & n57998) | (n57750 & n57998);
  assign n71350 = (n70942 & n71348) | (n70942 & n71349) | (n71348 & n71349);
  assign n58000 = n34353 | n34844;
  assign n71351 = n57751 | n58000;
  assign n71352 = n57750 | n58000;
  assign n71353 = (n70942 & n71351) | (n70942 & n71352) | (n71351 & n71352);
  assign n34847 = ~n71350 & n71353;
  assign n34848 = x153 & x201;
  assign n34849 = n34847 & n34848;
  assign n34850 = n34847 | n34848;
  assign n34851 = ~n34849 & n34850;
  assign n34852 = n71241 & n34851;
  assign n34853 = n71241 | n34851;
  assign n34854 = ~n34852 & n34853;
  assign n34855 = x152 & x202;
  assign n34856 = n34854 & n34855;
  assign n34857 = n34854 | n34855;
  assign n34858 = ~n34856 & n34857;
  assign n57869 = n34367 | n34369;
  assign n58002 = n34858 & n57869;
  assign n58003 = n34367 & n34858;
  assign n58004 = (n71083 & n58002) | (n71083 & n58003) | (n58002 & n58003);
  assign n58005 = n34858 | n57869;
  assign n58006 = n34367 | n34858;
  assign n58007 = (n71083 & n58005) | (n71083 & n58006) | (n58005 & n58006);
  assign n34861 = ~n58004 & n58007;
  assign n34862 = x151 & x203;
  assign n34863 = n34861 & n34862;
  assign n34864 = n34861 | n34862;
  assign n34865 = ~n34863 & n34864;
  assign n58008 = n34374 & n34865;
  assign n71354 = (n34865 & n57761) | (n34865 & n58008) | (n57761 & n58008);
  assign n71355 = (n34865 & n57760) | (n34865 & n58008) | (n57760 & n58008);
  assign n71356 = (n57365 & n71354) | (n57365 & n71355) | (n71354 & n71355);
  assign n58010 = n34374 | n34865;
  assign n71357 = n57761 | n58010;
  assign n71358 = n57760 | n58010;
  assign n71359 = (n57365 & n71357) | (n57365 & n71358) | (n71357 & n71358);
  assign n34868 = ~n71356 & n71359;
  assign n34869 = x150 & x204;
  assign n34870 = n34868 & n34869;
  assign n34871 = n34868 | n34869;
  assign n34872 = ~n34870 & n34871;
  assign n57867 = n34381 | n34383;
  assign n71360 = n34872 & n57867;
  assign n71235 = n33885 | n34381;
  assign n71236 = (n34381 & n34383) | (n34381 & n71235) | (n34383 & n71235);
  assign n71361 = n34872 & n71236;
  assign n71362 = (n71059 & n71360) | (n71059 & n71361) | (n71360 & n71361);
  assign n71363 = n34872 | n57867;
  assign n71364 = n34872 | n71236;
  assign n71365 = (n71059 & n71363) | (n71059 & n71364) | (n71363 & n71364);
  assign n34875 = ~n71362 & n71365;
  assign n34876 = x149 & x205;
  assign n34877 = n34875 & n34876;
  assign n34878 = n34875 | n34876;
  assign n34879 = ~n34877 & n34878;
  assign n58012 = n34388 & n34879;
  assign n71366 = (n34879 & n57770) | (n34879 & n58012) | (n57770 & n58012);
  assign n71367 = (n34390 & n34879) | (n34390 & n58012) | (n34879 & n58012);
  assign n71368 = (n57522 & n71366) | (n57522 & n71367) | (n71366 & n71367);
  assign n58014 = n34388 | n34879;
  assign n71369 = n57770 | n58014;
  assign n71370 = n34390 | n58014;
  assign n71371 = (n57522 & n71369) | (n57522 & n71370) | (n71369 & n71370);
  assign n34882 = ~n71368 & n71371;
  assign n34883 = x148 & x206;
  assign n34884 = n34882 & n34883;
  assign n34885 = n34882 | n34883;
  assign n34886 = ~n34884 & n34885;
  assign n58016 = n34395 & n34886;
  assign n58017 = (n34886 & n57775) | (n34886 & n58016) | (n57775 & n58016);
  assign n58018 = n34395 | n34886;
  assign n58019 = n57775 | n58018;
  assign n34889 = ~n58017 & n58019;
  assign n34890 = x147 & x207;
  assign n34891 = n34889 & n34890;
  assign n34892 = n34889 | n34890;
  assign n34893 = ~n34891 & n34892;
  assign n58020 = n34402 & n34893;
  assign n58021 = (n34893 & n57779) | (n34893 & n58020) | (n57779 & n58020);
  assign n58022 = n34402 | n34893;
  assign n58023 = n57779 | n58022;
  assign n34896 = ~n58021 & n58023;
  assign n34897 = x146 & x208;
  assign n34898 = n34896 & n34897;
  assign n34899 = n34896 | n34897;
  assign n34900 = ~n34898 & n34899;
  assign n58024 = n34409 & n34900;
  assign n58025 = (n34900 & n57783) | (n34900 & n58024) | (n57783 & n58024);
  assign n58026 = n34409 | n34900;
  assign n58027 = n57783 | n58026;
  assign n34903 = ~n58025 & n58027;
  assign n34904 = x145 & x209;
  assign n34905 = n34903 & n34904;
  assign n34906 = n34903 | n34904;
  assign n34907 = ~n34905 & n34906;
  assign n58028 = n34416 & n34907;
  assign n58029 = (n34907 & n57787) | (n34907 & n58028) | (n57787 & n58028);
  assign n58030 = n34416 | n34907;
  assign n58031 = n57787 | n58030;
  assign n34910 = ~n58029 & n58031;
  assign n34911 = x144 & x210;
  assign n34912 = n34910 & n34911;
  assign n34913 = n34910 | n34911;
  assign n34914 = ~n34912 & n34913;
  assign n58032 = n34423 & n34914;
  assign n58033 = (n34914 & n57791) | (n34914 & n58032) | (n57791 & n58032);
  assign n58034 = n34423 | n34914;
  assign n58035 = n57791 | n58034;
  assign n34917 = ~n58033 & n58035;
  assign n34918 = x143 & x211;
  assign n34919 = n34917 & n34918;
  assign n34920 = n34917 | n34918;
  assign n34921 = ~n34919 & n34920;
  assign n58036 = n34430 & n34921;
  assign n58037 = (n34921 & n57795) | (n34921 & n58036) | (n57795 & n58036);
  assign n58038 = n34430 | n34921;
  assign n58039 = n57795 | n58038;
  assign n34924 = ~n58037 & n58039;
  assign n34925 = x142 & x212;
  assign n34926 = n34924 & n34925;
  assign n34927 = n34924 | n34925;
  assign n34928 = ~n34926 & n34927;
  assign n58040 = n34437 & n34928;
  assign n58041 = (n34928 & n57799) | (n34928 & n58040) | (n57799 & n58040);
  assign n58042 = n34437 | n34928;
  assign n58043 = n57799 | n58042;
  assign n34931 = ~n58041 & n58043;
  assign n34932 = x141 & x213;
  assign n34933 = n34931 & n34932;
  assign n34934 = n34931 | n34932;
  assign n34935 = ~n34933 & n34934;
  assign n58044 = n34444 & n34935;
  assign n58045 = (n34935 & n57803) | (n34935 & n58044) | (n57803 & n58044);
  assign n58046 = n34444 | n34935;
  assign n58047 = n57803 | n58046;
  assign n34938 = ~n58045 & n58047;
  assign n34939 = x140 & x214;
  assign n34940 = n34938 & n34939;
  assign n34941 = n34938 | n34939;
  assign n34942 = ~n34940 & n34941;
  assign n58048 = n34451 & n34942;
  assign n58049 = (n34942 & n57807) | (n34942 & n58048) | (n57807 & n58048);
  assign n58050 = n34451 | n34942;
  assign n58051 = n57807 | n58050;
  assign n34945 = ~n58049 & n58051;
  assign n34946 = x139 & x215;
  assign n34947 = n34945 & n34946;
  assign n34948 = n34945 | n34946;
  assign n34949 = ~n34947 & n34948;
  assign n58052 = n34458 & n34949;
  assign n58053 = (n34949 & n57811) | (n34949 & n58052) | (n57811 & n58052);
  assign n58054 = n34458 | n34949;
  assign n58055 = n57811 | n58054;
  assign n34952 = ~n58053 & n58055;
  assign n34953 = x138 & x216;
  assign n34954 = n34952 & n34953;
  assign n34955 = n34952 | n34953;
  assign n34956 = ~n34954 & n34955;
  assign n58056 = n34465 & n34956;
  assign n58057 = (n34956 & n57815) | (n34956 & n58056) | (n57815 & n58056);
  assign n58058 = n34465 | n34956;
  assign n58059 = n57815 | n58058;
  assign n34959 = ~n58057 & n58059;
  assign n34960 = x137 & x217;
  assign n34961 = n34959 & n34960;
  assign n34962 = n34959 | n34960;
  assign n34963 = ~n34961 & n34962;
  assign n58060 = n34472 & n34963;
  assign n58061 = (n34963 & n57819) | (n34963 & n58060) | (n57819 & n58060);
  assign n58062 = n34472 | n34963;
  assign n58063 = n57819 | n58062;
  assign n34966 = ~n58061 & n58063;
  assign n34967 = x136 & x218;
  assign n34968 = n34966 & n34967;
  assign n34969 = n34966 | n34967;
  assign n34970 = ~n34968 & n34969;
  assign n58064 = n34479 & n34970;
  assign n58065 = (n34970 & n57823) | (n34970 & n58064) | (n57823 & n58064);
  assign n58066 = n34479 | n34970;
  assign n58067 = n57823 | n58066;
  assign n34973 = ~n58065 & n58067;
  assign n34974 = x135 & x219;
  assign n34975 = n34973 & n34974;
  assign n34976 = n34973 | n34974;
  assign n34977 = ~n34975 & n34976;
  assign n58068 = n34486 & n34977;
  assign n58069 = (n34977 & n57827) | (n34977 & n58068) | (n57827 & n58068);
  assign n58070 = n34486 | n34977;
  assign n58071 = n57827 | n58070;
  assign n34980 = ~n58069 & n58071;
  assign n34981 = x134 & x220;
  assign n34982 = n34980 & n34981;
  assign n34983 = n34980 | n34981;
  assign n34984 = ~n34982 & n34983;
  assign n58072 = n34493 & n34984;
  assign n58073 = (n34984 & n57831) | (n34984 & n58072) | (n57831 & n58072);
  assign n58074 = n34493 | n34984;
  assign n58075 = n57831 | n58074;
  assign n34987 = ~n58073 & n58075;
  assign n34988 = x133 & x221;
  assign n34989 = n34987 & n34988;
  assign n34990 = n34987 | n34988;
  assign n34991 = ~n34989 & n34990;
  assign n58076 = n34500 & n34991;
  assign n58077 = (n34991 & n57835) | (n34991 & n58076) | (n57835 & n58076);
  assign n58078 = n34500 | n34991;
  assign n58079 = n57835 | n58078;
  assign n34994 = ~n58077 & n58079;
  assign n34995 = x132 & x222;
  assign n34996 = n34994 & n34995;
  assign n34997 = n34994 | n34995;
  assign n34998 = ~n34996 & n34997;
  assign n58080 = n34507 & n34998;
  assign n58081 = (n34998 & n57839) | (n34998 & n58080) | (n57839 & n58080);
  assign n58082 = n34507 | n34998;
  assign n58083 = n57839 | n58082;
  assign n35001 = ~n58081 & n58083;
  assign n35002 = x131 & x223;
  assign n35003 = n35001 & n35002;
  assign n35004 = n35001 | n35002;
  assign n35005 = ~n35003 & n35004;
  assign n58084 = n34514 & n35005;
  assign n58085 = (n35005 & n57843) | (n35005 & n58084) | (n57843 & n58084);
  assign n58086 = n34514 | n35005;
  assign n58087 = n57843 | n58086;
  assign n35008 = ~n58085 & n58087;
  assign n35009 = x130 & x224;
  assign n35010 = n35008 & n35009;
  assign n35011 = n35008 | n35009;
  assign n35012 = ~n35010 & n35011;
  assign n58088 = n34521 & n35012;
  assign n58089 = (n35012 & n57848) | (n35012 & n58088) | (n57848 & n58088);
  assign n58090 = n34521 | n35012;
  assign n58091 = n57848 | n58090;
  assign n35015 = ~n58089 & n58091;
  assign n35016 = x129 & x225;
  assign n35017 = n35015 & n35016;
  assign n35018 = n35015 | n35016;
  assign n35019 = ~n35017 & n35018;
  assign n57864 = n34528 | n34530;
  assign n58092 = n35019 & n57864;
  assign n58093 = n34528 & n35019;
  assign n58094 = (n57610 & n58092) | (n57610 & n58093) | (n58092 & n58093);
  assign n58095 = n35019 | n57864;
  assign n58096 = n34528 | n35019;
  assign n58097 = (n57610 & n58095) | (n57610 & n58096) | (n58095 & n58096);
  assign n35022 = ~n58094 & n58097;
  assign n35023 = x128 & x226;
  assign n35024 = n35022 & n35023;
  assign n35025 = n35022 | n35023;
  assign n35026 = ~n35024 & n35025;
  assign n57862 = n34535 | n34537;
  assign n71372 = n35026 & n57862;
  assign n71373 = n34535 & n35026;
  assign n71374 = (n57608 & n71372) | (n57608 & n71373) | (n71372 & n71373);
  assign n71375 = n35026 | n57862;
  assign n71376 = n34535 | n35026;
  assign n71377 = (n57608 & n71375) | (n57608 & n71376) | (n71375 & n71376);
  assign n35029 = ~n71374 & n71377;
  assign n35030 = x127 & x227;
  assign n35031 = n35029 & n35030;
  assign n35032 = n35029 | n35030;
  assign n35033 = ~n35031 & n35032;
  assign n57860 = n34542 | n34544;
  assign n71378 = n35033 & n57860;
  assign n71379 = n34542 & n35033;
  assign n71380 = (n57606 & n71378) | (n57606 & n71379) | (n71378 & n71379);
  assign n71381 = n35033 | n57860;
  assign n71382 = n34542 | n35033;
  assign n71383 = (n57606 & n71381) | (n57606 & n71382) | (n71381 & n71382);
  assign n35036 = ~n71380 & n71383;
  assign n35037 = x126 & x228;
  assign n35038 = n35036 & n35037;
  assign n35039 = n35036 | n35037;
  assign n35040 = ~n35038 & n35039;
  assign n35041 = n57859 & n35040;
  assign n35042 = n57859 | n35040;
  assign n35043 = ~n35041 & n35042;
  assign n35044 = x125 & x229;
  assign n35045 = n35043 & n35044;
  assign n35046 = n35043 | n35044;
  assign n35047 = ~n35045 & n35046;
  assign n35048 = n57857 & n35047;
  assign n35049 = n57857 | n35047;
  assign n35050 = ~n35048 & n35049;
  assign n35051 = x124 & x230;
  assign n35052 = n35050 & n35051;
  assign n35053 = n35050 | n35051;
  assign n35054 = ~n35052 & n35053;
  assign n35055 = n34641 & n35054;
  assign n35056 = n34641 | n35054;
  assign n35057 = ~n35055 & n35056;
  assign n35058 = x123 & x231;
  assign n35059 = n35057 & n35058;
  assign n35060 = n35057 | n35058;
  assign n35061 = ~n35059 & n35060;
  assign n35062 = n34640 & n35061;
  assign n35063 = n34640 | n35061;
  assign n35064 = ~n35062 & n35063;
  assign n35065 = x122 & x232;
  assign n35066 = n35064 & n35065;
  assign n35067 = n35064 | n35065;
  assign n35068 = ~n35066 & n35067;
  assign n35069 = n34639 & n35068;
  assign n35070 = n34639 | n35068;
  assign n35071 = ~n35069 & n35070;
  assign n35072 = x121 & x233;
  assign n35073 = n35071 & n35072;
  assign n35074 = n35071 | n35072;
  assign n35075 = ~n35073 & n35074;
  assign n35076 = n34638 & n35075;
  assign n35077 = n34638 | n35075;
  assign n35078 = ~n35076 & n35077;
  assign n35079 = x120 & x234;
  assign n35080 = n35078 & n35079;
  assign n35081 = n35078 | n35079;
  assign n35082 = ~n35080 & n35081;
  assign n35083 = n34637 & n35082;
  assign n35084 = n34637 | n35082;
  assign n35085 = ~n35083 & n35084;
  assign n35086 = x119 & x235;
  assign n35087 = n35085 & n35086;
  assign n35088 = n35085 | n35086;
  assign n35089 = ~n35087 & n35088;
  assign n35090 = n34636 & n35089;
  assign n35091 = n34636 | n35089;
  assign n35092 = ~n35090 & n35091;
  assign n35093 = x118 & x236;
  assign n35094 = n35092 & n35093;
  assign n35095 = n35092 | n35093;
  assign n35096 = ~n35094 & n35095;
  assign n35097 = n34635 & n35096;
  assign n35098 = n34635 | n35096;
  assign n35099 = ~n35097 & n35098;
  assign n35100 = x117 & x237;
  assign n35101 = n35099 & n35100;
  assign n35102 = n35099 | n35100;
  assign n35103 = ~n35101 & n35102;
  assign n35104 = n71234 & n35103;
  assign n35105 = n71234 | n35103;
  assign n35106 = ~n35104 & n35105;
  assign n35107 = x116 & x238;
  assign n35108 = n35106 & n35107;
  assign n35109 = n35106 | n35107;
  assign n35110 = ~n35108 & n35109;
  assign n35111 = n57855 & n35110;
  assign n35112 = n57855 | n35110;
  assign n35113 = ~n35111 & n35112;
  assign n35114 = x115 & x239;
  assign n35115 = n35113 & n35114;
  assign n35116 = n35113 | n35114;
  assign n35117 = ~n35115 & n35116;
  assign n35118 = n57853 & n35117;
  assign n35119 = n57853 | n35117;
  assign n35120 = ~n35118 & n35119;
  assign n58098 = n35115 | n57853;
  assign n58099 = (n35115 & n35117) | (n35115 & n58098) | (n35117 & n58098);
  assign n58100 = n35108 | n57855;
  assign n58101 = (n35108 & n35110) | (n35108 & n58100) | (n35110 & n58100);
  assign n71384 = n35101 | n71234;
  assign n71385 = (n35101 & n35103) | (n35101 & n71384) | (n35103 & n71384);
  assign n35124 = n35094 | n35097;
  assign n35125 = n35087 | n35090;
  assign n35126 = n35080 | n35083;
  assign n35127 = n35073 | n35076;
  assign n35128 = n35066 | n35069;
  assign n35129 = n35059 | n35062;
  assign n58102 = n35052 | n35054;
  assign n58103 = (n34641 & n35052) | (n34641 & n58102) | (n35052 & n58102);
  assign n58104 = n35045 | n35047;
  assign n58105 = (n35045 & n57857) | (n35045 & n58104) | (n57857 & n58104);
  assign n57861 = (n34542 & n57606) | (n34542 & n57860) | (n57606 & n57860);
  assign n57863 = (n34535 & n57608) | (n34535 & n57862) | (n57608 & n57862);
  assign n57868 = (n71059 & n71236) | (n71059 & n57867) | (n71236 & n57867);
  assign n58115 = n34863 | n34865;
  assign n71386 = n34374 | n34863;
  assign n71387 = (n34863 & n34865) | (n34863 & n71386) | (n34865 & n71386);
  assign n71388 = (n57761 & n58115) | (n57761 & n71387) | (n58115 & n71387);
  assign n71389 = (n57760 & n58115) | (n57760 & n71387) | (n58115 & n71387);
  assign n71390 = (n57365 & n71388) | (n57365 & n71389) | (n71388 & n71389);
  assign n58120 = n34842 | n34844;
  assign n71391 = n34353 | n34842;
  assign n71392 = (n34842 & n34844) | (n34842 & n71391) | (n34844 & n71391);
  assign n71393 = (n57751 & n58120) | (n57751 & n71392) | (n58120 & n71392);
  assign n71394 = (n57750 & n58120) | (n57750 & n71392) | (n58120 & n71392);
  assign n71395 = (n70942 & n71393) | (n70942 & n71394) | (n71393 & n71394);
  assign n71402 = n34269 | n34758;
  assign n71403 = (n34758 & n34760) | (n34758 & n71402) | (n34760 & n71402);
  assign n71404 = n34758 | n34760;
  assign n71405 = (n34758 & n57894) | (n34758 & n71404) | (n57894 & n71404);
  assign n71406 = (n57639 & n71403) | (n57639 & n71405) | (n71403 & n71405);
  assign n71407 = (n71096 & n71403) | (n71096 & n71405) | (n71403 & n71405);
  assign n71408 = (n57154 & n71406) | (n57154 & n71407) | (n71406 & n71407);
  assign n57650 = (n70816 & n71105) | (n70816 & n71107) | (n71105 & n71107);
  assign n35182 = x175 & x180;
  assign n71411 = n34697 | n71279;
  assign n71413 = n35182 & n71411;
  assign n71414 = n35182 & n71279;
  assign n71415 = (n71287 & n71413) | (n71287 & n71414) | (n71413 & n71414);
  assign n71416 = (n35182 & n71289) | (n35182 & n71414) | (n71289 & n71414);
  assign n71417 = (n70995 & n71415) | (n70995 & n71416) | (n71415 & n71416);
  assign n71418 = (n70994 & n71415) | (n70994 & n71416) | (n71415 & n71416);
  assign n71419 = (n70013 & n71417) | (n70013 & n71418) | (n71417 & n71418);
  assign n71420 = n35182 | n71411;
  assign n71421 = n35182 | n71279;
  assign n71422 = (n71287 & n71420) | (n71287 & n71421) | (n71420 & n71421);
  assign n71423 = n71289 | n71421;
  assign n71424 = (n70995 & n71422) | (n70995 & n71423) | (n71422 & n71423);
  assign n71425 = (n70994 & n71422) | (n70994 & n71423) | (n71422 & n71423);
  assign n71426 = (n70013 & n71424) | (n70013 & n71425) | (n71424 & n71425);
  assign n35185 = ~n71419 & n71426;
  assign n71427 = n34702 | n34704;
  assign n71432 = (n34702 & n71301) | (n34702 & n71427) | (n71301 & n71427);
  assign n58170 = n35185 & n71432;
  assign n71429 = n35185 & n71427;
  assign n71430 = n34702 & n35185;
  assign n71431 = (n71299 & n71429) | (n71299 & n71430) | (n71429 & n71430);
  assign n71433 = (n58170 & n70971) | (n58170 & n71431) | (n70971 & n71431);
  assign n71434 = (n58170 & n70970) | (n58170 & n71431) | (n70970 & n71431);
  assign n71435 = (n70133 & n71433) | (n70133 & n71434) | (n71433 & n71434);
  assign n58173 = n35185 | n71432;
  assign n71436 = n35185 | n71427;
  assign n71437 = n34702 | n35185;
  assign n71438 = (n71299 & n71436) | (n71299 & n71437) | (n71436 & n71437);
  assign n71439 = (n58173 & n70971) | (n58173 & n71438) | (n70971 & n71438);
  assign n71440 = (n58173 & n70970) | (n58173 & n71438) | (n70970 & n71438);
  assign n71441 = (n70133 & n71439) | (n70133 & n71440) | (n71439 & n71440);
  assign n35188 = ~n71435 & n71441;
  assign n35189 = x174 & x181;
  assign n35190 = n35188 & n35189;
  assign n35191 = n35188 | n35189;
  assign n35192 = ~n35190 & n35191;
  assign n58155 = n34709 | n34711;
  assign n58175 = n35192 & n58155;
  assign n58176 = n34709 & n35192;
  assign n71442 = (n58175 & n58176) | (n58175 & n71273) | (n58176 & n71273);
  assign n71443 = (n58175 & n58176) | (n58175 & n71272) | (n58176 & n71272);
  assign n71444 = (n70822 & n71442) | (n70822 & n71443) | (n71442 & n71443);
  assign n58178 = n35192 | n58155;
  assign n58179 = n34709 | n35192;
  assign n71445 = (n58178 & n58179) | (n58178 & n71273) | (n58179 & n71273);
  assign n71446 = (n58178 & n58179) | (n58178 & n71272) | (n58179 & n71272);
  assign n71447 = (n70822 & n71445) | (n70822 & n71446) | (n71445 & n71446);
  assign n35195 = ~n71444 & n71447;
  assign n35196 = x173 & x182;
  assign n35197 = n35195 & n35196;
  assign n35198 = n35195 | n35196;
  assign n35199 = ~n35197 & n35198;
  assign n58181 = n34716 & n35199;
  assign n58182 = (n35199 & n71320) | (n35199 & n58181) | (n71320 & n58181);
  assign n58183 = n34716 | n35199;
  assign n58184 = n71320 | n58183;
  assign n35202 = ~n58182 & n58184;
  assign n35203 = x172 & x183;
  assign n35204 = n35202 & n35203;
  assign n35205 = n35202 | n35203;
  assign n35206 = ~n35204 & n35205;
  assign n71448 = n34234 | n34723;
  assign n71449 = (n34723 & n34725) | (n34723 & n71448) | (n34725 & n71448);
  assign n58185 = n35206 & n71449;
  assign n58153 = n34723 | n34725;
  assign n58186 = n35206 & n58153;
  assign n71450 = (n57698 & n58185) | (n57698 & n58186) | (n58185 & n58186);
  assign n71451 = (n57699 & n58185) | (n57699 & n58186) | (n58185 & n58186);
  assign n71452 = (n57167 & n71450) | (n57167 & n71451) | (n71450 & n71451);
  assign n58188 = n35206 | n71449;
  assign n58189 = n35206 | n58153;
  assign n71453 = (n57698 & n58188) | (n57698 & n58189) | (n58188 & n58189);
  assign n71454 = (n57699 & n58188) | (n57699 & n58189) | (n58188 & n58189);
  assign n71455 = (n57167 & n71453) | (n57167 & n71454) | (n71453 & n71454);
  assign n35209 = ~n71452 & n71455;
  assign n35210 = x171 & x184;
  assign n35211 = n35209 & n35210;
  assign n35212 = n35209 | n35210;
  assign n35213 = ~n35211 & n35212;
  assign n71456 = n34730 | n34732;
  assign n71457 = (n34730 & n57904) | (n34730 & n71456) | (n57904 & n71456);
  assign n58191 = n35213 & n71457;
  assign n71458 = n34241 | n34730;
  assign n71459 = (n34730 & n34732) | (n34730 & n71458) | (n34732 & n71458);
  assign n58192 = n35213 & n71459;
  assign n58193 = (n57650 & n58191) | (n57650 & n58192) | (n58191 & n58192);
  assign n58194 = n35213 | n71457;
  assign n58195 = n35213 | n71459;
  assign n58196 = (n57650 & n58194) | (n57650 & n58195) | (n58194 & n58195);
  assign n35216 = ~n58193 & n58196;
  assign n35217 = x170 & x185;
  assign n35218 = n35216 & n35217;
  assign n35219 = n35216 | n35217;
  assign n35220 = ~n35218 & n35219;
  assign n58147 = n34737 | n34739;
  assign n58197 = n35220 & n58147;
  assign n58198 = n34737 & n35220;
  assign n58199 = (n71270 & n58197) | (n71270 & n58198) | (n58197 & n58198);
  assign n58200 = n35220 | n58147;
  assign n58201 = n34737 | n35220;
  assign n58202 = (n71270 & n58200) | (n71270 & n58201) | (n58200 & n58201);
  assign n35223 = ~n58199 & n58202;
  assign n35224 = x169 & x186;
  assign n35225 = n35223 & n35224;
  assign n35226 = n35223 | n35224;
  assign n35227 = ~n35225 & n35226;
  assign n58145 = n34744 | n57950;
  assign n71460 = n35227 & n58145;
  assign n71409 = n34255 | n34744;
  assign n71410 = (n34744 & n34746) | (n34744 & n71409) | (n34746 & n71409);
  assign n71461 = n35227 & n71410;
  assign n71462 = (n71103 & n71460) | (n71103 & n71461) | (n71460 & n71461);
  assign n71463 = n35227 | n58145;
  assign n71464 = n35227 | n71410;
  assign n71465 = (n71103 & n71463) | (n71103 & n71464) | (n71463 & n71464);
  assign n35230 = ~n71462 & n71465;
  assign n35231 = x168 & x187;
  assign n35232 = n35230 & n35231;
  assign n35233 = n35230 | n35231;
  assign n35234 = ~n35232 & n35233;
  assign n58142 = n34751 | n34753;
  assign n58203 = n35234 & n58142;
  assign n58204 = n34751 & n35234;
  assign n71466 = (n57897 & n58203) | (n57897 & n58204) | (n58203 & n58204);
  assign n71467 = (n58203 & n58204) | (n58203 & n71263) | (n58204 & n71263);
  assign n71468 = (n70964 & n71466) | (n70964 & n71467) | (n71466 & n71467);
  assign n58206 = n35234 | n58142;
  assign n58207 = n34751 | n35234;
  assign n71469 = (n57897 & n58206) | (n57897 & n58207) | (n58206 & n58207);
  assign n71470 = (n58206 & n58207) | (n58206 & n71263) | (n58207 & n71263);
  assign n71471 = (n70964 & n71469) | (n70964 & n71470) | (n71469 & n71470);
  assign n35237 = ~n71468 & n71471;
  assign n35238 = x167 & x188;
  assign n35239 = n35237 & n35238;
  assign n35240 = n35237 | n35238;
  assign n35241 = ~n35239 & n35240;
  assign n35242 = n71408 & n35241;
  assign n35243 = n71408 | n35241;
  assign n35244 = ~n35242 & n35243;
  assign n35245 = x166 & x189;
  assign n35246 = n35244 & n35245;
  assign n35247 = n35244 | n35245;
  assign n35248 = ~n35246 & n35247;
  assign n58137 = n34765 | n34767;
  assign n58209 = n35248 & n58137;
  assign n58210 = n34765 & n35248;
  assign n58211 = (n71261 & n58209) | (n71261 & n58210) | (n58209 & n58210);
  assign n58212 = n35248 | n58137;
  assign n58213 = n34765 | n35248;
  assign n58214 = (n71261 & n58212) | (n71261 & n58213) | (n58212 & n58213);
  assign n35251 = ~n58211 & n58214;
  assign n35252 = x165 & x190;
  assign n35253 = n35251 & n35252;
  assign n35254 = n35251 | n35252;
  assign n35255 = ~n35253 & n35254;
  assign n58215 = n34772 & n35255;
  assign n71472 = (n35255 & n57963) | (n35255 & n58215) | (n57963 & n58215);
  assign n71473 = (n35255 & n57962) | (n35255 & n58215) | (n57962 & n58215);
  assign n71474 = (n57637 & n71472) | (n57637 & n71473) | (n71472 & n71473);
  assign n58217 = n34772 | n35255;
  assign n71475 = n57963 | n58217;
  assign n71476 = n57962 | n58217;
  assign n71477 = (n57637 & n71475) | (n57637 & n71476) | (n71475 & n71476);
  assign n35258 = ~n71474 & n71477;
  assign n35259 = x164 & x191;
  assign n35260 = n35258 & n35259;
  assign n35261 = n35258 | n35259;
  assign n35262 = ~n35260 & n35261;
  assign n58135 = n34779 | n34781;
  assign n71478 = n35262 & n58135;
  assign n71400 = n34290 | n34779;
  assign n71401 = (n34779 & n34781) | (n34779 & n71400) | (n34781 & n71400);
  assign n71479 = n35262 & n71401;
  assign n71480 = (n57722 & n71478) | (n57722 & n71479) | (n71478 & n71479);
  assign n71481 = n35262 | n58135;
  assign n71482 = n35262 | n71401;
  assign n71483 = (n57722 & n71481) | (n57722 & n71482) | (n71481 & n71482);
  assign n35265 = ~n71480 & n71483;
  assign n35266 = x163 & x192;
  assign n35267 = n35265 & n35266;
  assign n35268 = n35265 | n35266;
  assign n35269 = ~n35267 & n35268;
  assign n58132 = n34786 | n34788;
  assign n58219 = n35269 & n58132;
  assign n58220 = n34786 & n35269;
  assign n58221 = (n71256 & n58219) | (n71256 & n58220) | (n58219 & n58220);
  assign n58222 = n35269 | n58132;
  assign n58223 = n34786 | n35269;
  assign n58224 = (n71256 & n58222) | (n71256 & n58223) | (n58222 & n58223);
  assign n35272 = ~n58221 & n58224;
  assign n35273 = x162 & x193;
  assign n35274 = n35272 & n35273;
  assign n35275 = n35272 | n35273;
  assign n35276 = ~n35274 & n35275;
  assign n58225 = n34793 & n35276;
  assign n71484 = (n35276 & n57973) | (n35276 & n58225) | (n57973 & n58225);
  assign n71485 = (n35276 & n57972) | (n35276 & n58225) | (n57972 & n58225);
  assign n71486 = (n57632 & n71484) | (n57632 & n71485) | (n71484 & n71485);
  assign n58227 = n34793 | n35276;
  assign n71487 = n57973 | n58227;
  assign n71488 = n57972 | n58227;
  assign n71489 = (n57632 & n71487) | (n57632 & n71488) | (n71487 & n71488);
  assign n35279 = ~n71486 & n71489;
  assign n35280 = x161 & x194;
  assign n35281 = n35279 & n35280;
  assign n35282 = n35279 | n35280;
  assign n35283 = ~n35281 & n35282;
  assign n58130 = n34800 | n34802;
  assign n71490 = n35283 & n58130;
  assign n71398 = n34311 | n34800;
  assign n71399 = (n34800 & n34802) | (n34800 & n71398) | (n34802 & n71398);
  assign n71491 = n35283 & n71399;
  assign n71492 = (n57732 & n71490) | (n57732 & n71491) | (n71490 & n71491);
  assign n71493 = n35283 | n58130;
  assign n71494 = n35283 | n71399;
  assign n71495 = (n57732 & n71493) | (n57732 & n71494) | (n71493 & n71494);
  assign n35286 = ~n71492 & n71495;
  assign n35287 = x160 & x195;
  assign n35288 = n35286 & n35287;
  assign n35289 = n35286 | n35287;
  assign n35290 = ~n35288 & n35289;
  assign n58127 = n34807 | n34809;
  assign n58229 = n35290 & n58127;
  assign n58230 = n34807 & n35290;
  assign n58231 = (n71251 & n58229) | (n71251 & n58230) | (n58229 & n58230);
  assign n58232 = n35290 | n58127;
  assign n58233 = n34807 | n35290;
  assign n58234 = (n71251 & n58232) | (n71251 & n58233) | (n58232 & n58233);
  assign n35293 = ~n58231 & n58234;
  assign n35294 = x159 & x196;
  assign n35295 = n35293 & n35294;
  assign n35296 = n35293 | n35294;
  assign n35297 = ~n35295 & n35296;
  assign n58235 = n34814 & n35297;
  assign n71496 = (n35297 & n57983) | (n35297 & n58235) | (n57983 & n58235);
  assign n71497 = (n35297 & n57982) | (n35297 & n58235) | (n57982 & n58235);
  assign n71498 = (n57627 & n71496) | (n57627 & n71497) | (n71496 & n71497);
  assign n58237 = n34814 | n35297;
  assign n71499 = n57983 | n58237;
  assign n71500 = n57982 | n58237;
  assign n71501 = (n57627 & n71499) | (n57627 & n71500) | (n71499 & n71500);
  assign n35300 = ~n71498 & n71501;
  assign n35301 = x158 & x197;
  assign n35302 = n35300 & n35301;
  assign n35303 = n35300 | n35301;
  assign n35304 = ~n35302 & n35303;
  assign n58125 = n34821 | n34823;
  assign n71502 = n35304 & n58125;
  assign n71396 = n34332 | n34821;
  assign n71397 = (n34821 & n34823) | (n34821 & n71396) | (n34823 & n71396);
  assign n71503 = n35304 & n71397;
  assign n71504 = (n57742 & n71502) | (n57742 & n71503) | (n71502 & n71503);
  assign n71505 = n35304 | n58125;
  assign n71506 = n35304 | n71397;
  assign n71507 = (n57742 & n71505) | (n57742 & n71506) | (n71505 & n71506);
  assign n35307 = ~n71504 & n71507;
  assign n35308 = x157 & x198;
  assign n35309 = n35307 & n35308;
  assign n35310 = n35307 | n35308;
  assign n35311 = ~n35309 & n35310;
  assign n58122 = n34828 | n34830;
  assign n58239 = n35311 & n58122;
  assign n58240 = n34828 & n35311;
  assign n58241 = (n71246 & n58239) | (n71246 & n58240) | (n58239 & n58240);
  assign n58242 = n35311 | n58122;
  assign n58243 = n34828 | n35311;
  assign n58244 = (n71246 & n58242) | (n71246 & n58243) | (n58242 & n58243);
  assign n35314 = ~n58241 & n58244;
  assign n35315 = x156 & x199;
  assign n35316 = n35314 & n35315;
  assign n35317 = n35314 | n35315;
  assign n35318 = ~n35316 & n35317;
  assign n58245 = n34835 & n35318;
  assign n71508 = (n35318 & n57993) | (n35318 & n58245) | (n57993 & n58245);
  assign n71509 = (n35318 & n57992) | (n35318 & n58245) | (n57992 & n58245);
  assign n71510 = (n71088 & n71508) | (n71088 & n71509) | (n71508 & n71509);
  assign n58247 = n34835 | n35318;
  assign n71511 = n57993 | n58247;
  assign n71512 = n57992 | n58247;
  assign n71513 = (n71088 & n71511) | (n71088 & n71512) | (n71511 & n71512);
  assign n35321 = ~n71510 & n71513;
  assign n35322 = x155 & x200;
  assign n35323 = n35321 & n35322;
  assign n35324 = n35321 | n35322;
  assign n35325 = ~n35323 & n35324;
  assign n35326 = n71395 & n35325;
  assign n35327 = n71395 | n35325;
  assign n35328 = ~n35326 & n35327;
  assign n35329 = x154 & x201;
  assign n35330 = n35328 & n35329;
  assign n35331 = n35328 | n35329;
  assign n35332 = ~n35330 & n35331;
  assign n58117 = n34849 | n34851;
  assign n58249 = n35332 & n58117;
  assign n58250 = n34849 & n35332;
  assign n58251 = (n71241 & n58249) | (n71241 & n58250) | (n58249 & n58250);
  assign n58252 = n35332 | n58117;
  assign n58253 = n34849 | n35332;
  assign n58254 = (n71241 & n58252) | (n71241 & n58253) | (n58252 & n58253);
  assign n35335 = ~n58251 & n58254;
  assign n35336 = x153 & x202;
  assign n35337 = n35335 & n35336;
  assign n35338 = n35335 | n35336;
  assign n35339 = ~n35337 & n35338;
  assign n58255 = n34856 & n35339;
  assign n71514 = (n35339 & n58003) | (n35339 & n58255) | (n58003 & n58255);
  assign n71515 = (n35339 & n58002) | (n35339 & n58255) | (n58002 & n58255);
  assign n71516 = (n71083 & n71514) | (n71083 & n71515) | (n71514 & n71515);
  assign n58257 = n34856 | n35339;
  assign n71517 = n58003 | n58257;
  assign n71518 = n58002 | n58257;
  assign n71519 = (n71083 & n71517) | (n71083 & n71518) | (n71517 & n71518);
  assign n35342 = ~n71516 & n71519;
  assign n35343 = x152 & x203;
  assign n35344 = n35342 & n35343;
  assign n35345 = n35342 | n35343;
  assign n35346 = ~n35344 & n35345;
  assign n35347 = n71390 & n35346;
  assign n35348 = n71390 | n35346;
  assign n35349 = ~n35347 & n35348;
  assign n35350 = x151 & x204;
  assign n35351 = n35349 & n35350;
  assign n35352 = n35349 | n35350;
  assign n35353 = ~n35351 & n35352;
  assign n58112 = n34870 | n34872;
  assign n58259 = n35353 & n58112;
  assign n58260 = n34870 & n35353;
  assign n58261 = (n57868 & n58259) | (n57868 & n58260) | (n58259 & n58260);
  assign n58262 = n35353 | n58112;
  assign n58263 = n34870 | n35353;
  assign n58264 = (n57868 & n58262) | (n57868 & n58263) | (n58262 & n58263);
  assign n35356 = ~n58261 & n58264;
  assign n35357 = x150 & x205;
  assign n35358 = n35356 & n35357;
  assign n35359 = n35356 | n35357;
  assign n35360 = ~n35358 & n35359;
  assign n58265 = n34877 & n35360;
  assign n58266 = (n35360 & n71368) | (n35360 & n58265) | (n71368 & n58265);
  assign n58267 = n34877 | n35360;
  assign n58268 = n71368 | n58267;
  assign n35363 = ~n58266 & n58268;
  assign n35364 = x149 & x206;
  assign n35365 = n35363 & n35364;
  assign n35366 = n35363 | n35364;
  assign n35367 = ~n35365 & n35366;
  assign n58269 = n34884 & n35367;
  assign n58270 = (n35367 & n58017) | (n35367 & n58269) | (n58017 & n58269);
  assign n58271 = n34884 | n35367;
  assign n58272 = n58017 | n58271;
  assign n35370 = ~n58270 & n58272;
  assign n35371 = x148 & x207;
  assign n35372 = n35370 & n35371;
  assign n35373 = n35370 | n35371;
  assign n35374 = ~n35372 & n35373;
  assign n58273 = n34891 & n35374;
  assign n58274 = (n35374 & n58021) | (n35374 & n58273) | (n58021 & n58273);
  assign n58275 = n34891 | n35374;
  assign n58276 = n58021 | n58275;
  assign n35377 = ~n58274 & n58276;
  assign n35378 = x147 & x208;
  assign n35379 = n35377 & n35378;
  assign n35380 = n35377 | n35378;
  assign n35381 = ~n35379 & n35380;
  assign n58277 = n34898 & n35381;
  assign n58278 = (n35381 & n58025) | (n35381 & n58277) | (n58025 & n58277);
  assign n58279 = n34898 | n35381;
  assign n58280 = n58025 | n58279;
  assign n35384 = ~n58278 & n58280;
  assign n35385 = x146 & x209;
  assign n35386 = n35384 & n35385;
  assign n35387 = n35384 | n35385;
  assign n35388 = ~n35386 & n35387;
  assign n58281 = n34905 & n35388;
  assign n58282 = (n35388 & n58029) | (n35388 & n58281) | (n58029 & n58281);
  assign n58283 = n34905 | n35388;
  assign n58284 = n58029 | n58283;
  assign n35391 = ~n58282 & n58284;
  assign n35392 = x145 & x210;
  assign n35393 = n35391 & n35392;
  assign n35394 = n35391 | n35392;
  assign n35395 = ~n35393 & n35394;
  assign n58285 = n34912 & n35395;
  assign n58286 = (n35395 & n58033) | (n35395 & n58285) | (n58033 & n58285);
  assign n58287 = n34912 | n35395;
  assign n58288 = n58033 | n58287;
  assign n35398 = ~n58286 & n58288;
  assign n35399 = x144 & x211;
  assign n35400 = n35398 & n35399;
  assign n35401 = n35398 | n35399;
  assign n35402 = ~n35400 & n35401;
  assign n58289 = n34919 & n35402;
  assign n58290 = (n35402 & n58037) | (n35402 & n58289) | (n58037 & n58289);
  assign n58291 = n34919 | n35402;
  assign n58292 = n58037 | n58291;
  assign n35405 = ~n58290 & n58292;
  assign n35406 = x143 & x212;
  assign n35407 = n35405 & n35406;
  assign n35408 = n35405 | n35406;
  assign n35409 = ~n35407 & n35408;
  assign n58293 = n34926 & n35409;
  assign n58294 = (n35409 & n58041) | (n35409 & n58293) | (n58041 & n58293);
  assign n58295 = n34926 | n35409;
  assign n58296 = n58041 | n58295;
  assign n35412 = ~n58294 & n58296;
  assign n35413 = x142 & x213;
  assign n35414 = n35412 & n35413;
  assign n35415 = n35412 | n35413;
  assign n35416 = ~n35414 & n35415;
  assign n58297 = n34933 & n35416;
  assign n58298 = (n35416 & n58045) | (n35416 & n58297) | (n58045 & n58297);
  assign n58299 = n34933 | n35416;
  assign n58300 = n58045 | n58299;
  assign n35419 = ~n58298 & n58300;
  assign n35420 = x141 & x214;
  assign n35421 = n35419 & n35420;
  assign n35422 = n35419 | n35420;
  assign n35423 = ~n35421 & n35422;
  assign n58301 = n34940 & n35423;
  assign n58302 = (n35423 & n58049) | (n35423 & n58301) | (n58049 & n58301);
  assign n58303 = n34940 | n35423;
  assign n58304 = n58049 | n58303;
  assign n35426 = ~n58302 & n58304;
  assign n35427 = x140 & x215;
  assign n35428 = n35426 & n35427;
  assign n35429 = n35426 | n35427;
  assign n35430 = ~n35428 & n35429;
  assign n58305 = n34947 & n35430;
  assign n58306 = (n35430 & n58053) | (n35430 & n58305) | (n58053 & n58305);
  assign n58307 = n34947 | n35430;
  assign n58308 = n58053 | n58307;
  assign n35433 = ~n58306 & n58308;
  assign n35434 = x139 & x216;
  assign n35435 = n35433 & n35434;
  assign n35436 = n35433 | n35434;
  assign n35437 = ~n35435 & n35436;
  assign n58309 = n34954 & n35437;
  assign n58310 = (n35437 & n58057) | (n35437 & n58309) | (n58057 & n58309);
  assign n58311 = n34954 | n35437;
  assign n58312 = n58057 | n58311;
  assign n35440 = ~n58310 & n58312;
  assign n35441 = x138 & x217;
  assign n35442 = n35440 & n35441;
  assign n35443 = n35440 | n35441;
  assign n35444 = ~n35442 & n35443;
  assign n58313 = n34961 & n35444;
  assign n58314 = (n35444 & n58061) | (n35444 & n58313) | (n58061 & n58313);
  assign n58315 = n34961 | n35444;
  assign n58316 = n58061 | n58315;
  assign n35447 = ~n58314 & n58316;
  assign n35448 = x137 & x218;
  assign n35449 = n35447 & n35448;
  assign n35450 = n35447 | n35448;
  assign n35451 = ~n35449 & n35450;
  assign n58317 = n34968 & n35451;
  assign n58318 = (n35451 & n58065) | (n35451 & n58317) | (n58065 & n58317);
  assign n58319 = n34968 | n35451;
  assign n58320 = n58065 | n58319;
  assign n35454 = ~n58318 & n58320;
  assign n35455 = x136 & x219;
  assign n35456 = n35454 & n35455;
  assign n35457 = n35454 | n35455;
  assign n35458 = ~n35456 & n35457;
  assign n58321 = n34975 & n35458;
  assign n58322 = (n35458 & n58069) | (n35458 & n58321) | (n58069 & n58321);
  assign n58323 = n34975 | n35458;
  assign n58324 = n58069 | n58323;
  assign n35461 = ~n58322 & n58324;
  assign n35462 = x135 & x220;
  assign n35463 = n35461 & n35462;
  assign n35464 = n35461 | n35462;
  assign n35465 = ~n35463 & n35464;
  assign n58325 = n34982 & n35465;
  assign n58326 = (n35465 & n58073) | (n35465 & n58325) | (n58073 & n58325);
  assign n58327 = n34982 | n35465;
  assign n58328 = n58073 | n58327;
  assign n35468 = ~n58326 & n58328;
  assign n35469 = x134 & x221;
  assign n35470 = n35468 & n35469;
  assign n35471 = n35468 | n35469;
  assign n35472 = ~n35470 & n35471;
  assign n58329 = n34989 & n35472;
  assign n58330 = (n35472 & n58077) | (n35472 & n58329) | (n58077 & n58329);
  assign n58331 = n34989 | n35472;
  assign n58332 = n58077 | n58331;
  assign n35475 = ~n58330 & n58332;
  assign n35476 = x133 & x222;
  assign n35477 = n35475 & n35476;
  assign n35478 = n35475 | n35476;
  assign n35479 = ~n35477 & n35478;
  assign n58333 = n34996 & n35479;
  assign n58334 = (n35479 & n58081) | (n35479 & n58333) | (n58081 & n58333);
  assign n58335 = n34996 | n35479;
  assign n58336 = n58081 | n58335;
  assign n35482 = ~n58334 & n58336;
  assign n35483 = x132 & x223;
  assign n35484 = n35482 & n35483;
  assign n35485 = n35482 | n35483;
  assign n35486 = ~n35484 & n35485;
  assign n58337 = n35003 & n35486;
  assign n58338 = (n35486 & n58085) | (n35486 & n58337) | (n58085 & n58337);
  assign n58339 = n35003 | n35486;
  assign n58340 = n58085 | n58339;
  assign n35489 = ~n58338 & n58340;
  assign n35490 = x131 & x224;
  assign n35491 = n35489 & n35490;
  assign n35492 = n35489 | n35490;
  assign n35493 = ~n35491 & n35492;
  assign n58341 = n35010 & n35493;
  assign n58342 = (n35493 & n58089) | (n35493 & n58341) | (n58089 & n58341);
  assign n58343 = n35010 | n35493;
  assign n58344 = n58089 | n58343;
  assign n35496 = ~n58342 & n58344;
  assign n35497 = x130 & x225;
  assign n35498 = n35496 & n35497;
  assign n35499 = n35496 | n35497;
  assign n35500 = ~n35498 & n35499;
  assign n58345 = n35017 & n35500;
  assign n58346 = (n35500 & n58094) | (n35500 & n58345) | (n58094 & n58345);
  assign n58347 = n35017 | n35500;
  assign n58348 = n58094 | n58347;
  assign n35503 = ~n58346 & n58348;
  assign n35504 = x129 & x226;
  assign n35505 = n35503 & n35504;
  assign n35506 = n35503 | n35504;
  assign n35507 = ~n35505 & n35506;
  assign n58110 = n35024 | n35026;
  assign n58349 = n35507 & n58110;
  assign n58350 = n35024 & n35507;
  assign n58351 = (n57863 & n58349) | (n57863 & n58350) | (n58349 & n58350);
  assign n58352 = n35507 | n58110;
  assign n58353 = n35024 | n35507;
  assign n58354 = (n57863 & n58352) | (n57863 & n58353) | (n58352 & n58353);
  assign n35510 = ~n58351 & n58354;
  assign n35511 = x128 & x227;
  assign n35512 = n35510 & n35511;
  assign n35513 = n35510 | n35511;
  assign n35514 = ~n35512 & n35513;
  assign n58108 = n35031 | n35033;
  assign n71520 = n35514 & n58108;
  assign n71521 = n35031 & n35514;
  assign n71522 = (n57861 & n71520) | (n57861 & n71521) | (n71520 & n71521);
  assign n71523 = n35514 | n58108;
  assign n71524 = n35031 | n35514;
  assign n71525 = (n57861 & n71523) | (n57861 & n71524) | (n71523 & n71524);
  assign n35517 = ~n71522 & n71525;
  assign n35518 = x127 & x228;
  assign n35519 = n35517 & n35518;
  assign n35520 = n35517 | n35518;
  assign n35521 = ~n35519 & n35520;
  assign n58106 = n35038 | n35040;
  assign n71526 = n35521 & n58106;
  assign n71527 = n35038 & n35521;
  assign n71528 = (n57859 & n71526) | (n57859 & n71527) | (n71526 & n71527);
  assign n71529 = n35521 | n58106;
  assign n71530 = n35038 | n35521;
  assign n71531 = (n57859 & n71529) | (n57859 & n71530) | (n71529 & n71530);
  assign n35524 = ~n71528 & n71531;
  assign n35525 = x126 & x229;
  assign n35526 = n35524 & n35525;
  assign n35527 = n35524 | n35525;
  assign n35528 = ~n35526 & n35527;
  assign n35529 = n58105 & n35528;
  assign n35530 = n58105 | n35528;
  assign n35531 = ~n35529 & n35530;
  assign n35532 = x125 & x230;
  assign n35533 = n35531 & n35532;
  assign n35534 = n35531 | n35532;
  assign n35535 = ~n35533 & n35534;
  assign n35536 = n58103 & n35535;
  assign n35537 = n58103 | n35535;
  assign n35538 = ~n35536 & n35537;
  assign n35539 = x124 & x231;
  assign n35540 = n35538 & n35539;
  assign n35541 = n35538 | n35539;
  assign n35542 = ~n35540 & n35541;
  assign n35543 = n35129 & n35542;
  assign n35544 = n35129 | n35542;
  assign n35545 = ~n35543 & n35544;
  assign n35546 = x123 & x232;
  assign n35547 = n35545 & n35546;
  assign n35548 = n35545 | n35546;
  assign n35549 = ~n35547 & n35548;
  assign n35550 = n35128 & n35549;
  assign n35551 = n35128 | n35549;
  assign n35552 = ~n35550 & n35551;
  assign n35553 = x122 & x233;
  assign n35554 = n35552 & n35553;
  assign n35555 = n35552 | n35553;
  assign n35556 = ~n35554 & n35555;
  assign n35557 = n35127 & n35556;
  assign n35558 = n35127 | n35556;
  assign n35559 = ~n35557 & n35558;
  assign n35560 = x121 & x234;
  assign n35561 = n35559 & n35560;
  assign n35562 = n35559 | n35560;
  assign n35563 = ~n35561 & n35562;
  assign n35564 = n35126 & n35563;
  assign n35565 = n35126 | n35563;
  assign n35566 = ~n35564 & n35565;
  assign n35567 = x120 & x235;
  assign n35568 = n35566 & n35567;
  assign n35569 = n35566 | n35567;
  assign n35570 = ~n35568 & n35569;
  assign n35571 = n35125 & n35570;
  assign n35572 = n35125 | n35570;
  assign n35573 = ~n35571 & n35572;
  assign n35574 = x119 & x236;
  assign n35575 = n35573 & n35574;
  assign n35576 = n35573 | n35574;
  assign n35577 = ~n35575 & n35576;
  assign n35578 = n35124 & n35577;
  assign n35579 = n35124 | n35577;
  assign n35580 = ~n35578 & n35579;
  assign n35581 = x118 & x237;
  assign n35582 = n35580 & n35581;
  assign n35583 = n35580 | n35581;
  assign n35584 = ~n35582 & n35583;
  assign n35585 = n71385 & n35584;
  assign n35586 = n71385 | n35584;
  assign n35587 = ~n35585 & n35586;
  assign n35588 = x117 & x238;
  assign n35589 = n35587 & n35588;
  assign n35590 = n35587 | n35588;
  assign n35591 = ~n35589 & n35590;
  assign n35592 = n58101 & n35591;
  assign n35593 = n58101 | n35591;
  assign n35594 = ~n35592 & n35593;
  assign n35595 = x116 & x239;
  assign n35596 = n35594 & n35595;
  assign n35597 = n35594 | n35595;
  assign n35598 = ~n35596 & n35597;
  assign n35599 = n58099 & n35598;
  assign n35600 = n58099 | n35598;
  assign n35601 = ~n35599 & n35600;
  assign n58355 = n35596 | n58099;
  assign n58356 = (n35596 & n35598) | (n35596 & n58355) | (n35598 & n58355);
  assign n58357 = n35589 | n58101;
  assign n58358 = (n35589 & n35591) | (n35589 & n58357) | (n35591 & n58357);
  assign n71532 = n35582 | n71385;
  assign n71533 = (n35582 & n35584) | (n35582 & n71532) | (n35584 & n71532);
  assign n35605 = n35575 | n35578;
  assign n35606 = n35568 | n35571;
  assign n35607 = n35561 | n35564;
  assign n35608 = n35554 | n35557;
  assign n35609 = n35547 | n35550;
  assign n58359 = n35540 | n35542;
  assign n58360 = (n35129 & n35540) | (n35129 & n58359) | (n35540 & n58359);
  assign n58361 = n35533 | n35535;
  assign n58362 = (n35533 & n58103) | (n35533 & n58361) | (n58103 & n58361);
  assign n58107 = (n35038 & n57859) | (n35038 & n58106) | (n57859 & n58106);
  assign n58109 = (n35031 & n57861) | (n35031 & n58108) | (n57861 & n58108);
  assign n58375 = n35337 | n35339;
  assign n71536 = n34856 | n35337;
  assign n71537 = (n35337 & n35339) | (n35337 & n71536) | (n35339 & n71536);
  assign n71538 = (n58003 & n58375) | (n58003 & n71537) | (n58375 & n71537);
  assign n71539 = (n58002 & n58375) | (n58002 & n71537) | (n58375 & n71537);
  assign n71540 = (n71083 & n71538) | (n71083 & n71539) | (n71538 & n71539);
  assign n58380 = n35316 | n35318;
  assign n71541 = n34835 | n35316;
  assign n71542 = (n35316 & n35318) | (n35316 & n71541) | (n35318 & n71541);
  assign n71543 = (n57993 & n58380) | (n57993 & n71542) | (n58380 & n71542);
  assign n71544 = (n57992 & n58380) | (n57992 & n71542) | (n58380 & n71542);
  assign n71545 = (n71088 & n71543) | (n71088 & n71544) | (n71543 & n71544);
  assign n58126 = (n57742 & n71397) | (n57742 & n58125) | (n71397 & n58125);
  assign n58385 = n35295 | n35297;
  assign n71546 = n34814 | n35295;
  assign n71547 = (n35295 & n35297) | (n35295 & n71546) | (n35297 & n71546);
  assign n71548 = (n57983 & n58385) | (n57983 & n71547) | (n58385 & n71547);
  assign n71549 = (n57982 & n58385) | (n57982 & n71547) | (n58385 & n71547);
  assign n71550 = (n57627 & n71548) | (n57627 & n71549) | (n71548 & n71549);
  assign n58131 = (n57732 & n71399) | (n57732 & n58130) | (n71399 & n58130);
  assign n58390 = n35274 | n35276;
  assign n71551 = n34793 | n35274;
  assign n71552 = (n35274 & n35276) | (n35274 & n71551) | (n35276 & n71551);
  assign n71553 = (n57973 & n58390) | (n57973 & n71552) | (n58390 & n71552);
  assign n71554 = (n57972 & n58390) | (n57972 & n71552) | (n58390 & n71552);
  assign n71555 = (n57632 & n71553) | (n57632 & n71554) | (n71553 & n71554);
  assign n58136 = (n57722 & n71401) | (n57722 & n58135) | (n71401 & n58135);
  assign n58395 = n35253 | n35255;
  assign n71556 = n34772 | n35253;
  assign n71557 = (n35253 & n35255) | (n35253 & n71556) | (n35255 & n71556);
  assign n71558 = (n57963 & n58395) | (n57963 & n71557) | (n58395 & n71557);
  assign n71559 = (n57962 & n58395) | (n57962 & n71557) | (n58395 & n71557);
  assign n71560 = (n57637 & n71558) | (n57637 & n71559) | (n71558 & n71559);
  assign n71561 = n34765 | n35246;
  assign n71562 = (n35246 & n35248) | (n35246 & n71561) | (n35248 & n71561);
  assign n58398 = n35246 | n58209;
  assign n58399 = (n71261 & n71562) | (n71261 & n58398) | (n71562 & n58398);
  assign n71563 = n34751 | n35232;
  assign n71564 = (n35232 & n35234) | (n35232 & n71563) | (n35234 & n71563);
  assign n71565 = n35232 | n35234;
  assign n71566 = (n35232 & n58142) | (n35232 & n71565) | (n58142 & n71565);
  assign n71567 = (n57897 & n71564) | (n57897 & n71566) | (n71564 & n71566);
  assign n71568 = (n71263 & n71564) | (n71263 & n71566) | (n71564 & n71566);
  assign n71569 = (n70964 & n71567) | (n70964 & n71568) | (n71567 & n71568);
  assign n58410 = n35204 | n58185;
  assign n58411 = n35204 | n58186;
  assign n71572 = (n57698 & n58410) | (n57698 & n58411) | (n58410 & n58411);
  assign n71573 = (n57699 & n58410) | (n57699 & n58411) | (n58410 & n58411);
  assign n71574 = (n57167 & n71572) | (n57167 & n71573) | (n71572 & n71573);
  assign n35662 = x175 & x181;
  assign n58419 = n35662 & n71419;
  assign n58420 = (n35662 & n71435) | (n35662 & n58419) | (n71435 & n58419);
  assign n58421 = n35662 | n71419;
  assign n58422 = n71435 | n58421;
  assign n35665 = ~n58420 & n58422;
  assign n71575 = n35190 | n35192;
  assign n71576 = (n35190 & n58155) | (n35190 & n71575) | (n58155 & n71575);
  assign n58423 = n35665 & n71576;
  assign n71577 = n34709 | n35190;
  assign n71578 = (n35190 & n35192) | (n35190 & n71577) | (n35192 & n71577);
  assign n58424 = n35665 & n71578;
  assign n71579 = (n58423 & n58424) | (n58423 & n71273) | (n58424 & n71273);
  assign n71580 = (n58423 & n58424) | (n58423 & n71272) | (n58424 & n71272);
  assign n71581 = (n70822 & n71579) | (n70822 & n71580) | (n71579 & n71580);
  assign n58426 = n35665 | n71576;
  assign n58427 = n35665 | n71578;
  assign n71582 = (n58426 & n58427) | (n58426 & n71273) | (n58427 & n71273);
  assign n71583 = (n58426 & n58427) | (n58426 & n71272) | (n58427 & n71272);
  assign n71584 = (n70822 & n71582) | (n70822 & n71583) | (n71582 & n71583);
  assign n35668 = ~n71581 & n71584;
  assign n35669 = x174 & x182;
  assign n35670 = n35668 & n35669;
  assign n35671 = n35668 | n35669;
  assign n35672 = ~n35670 & n35671;
  assign n71585 = n34716 | n35197;
  assign n71586 = (n35197 & n35199) | (n35197 & n71585) | (n35199 & n71585);
  assign n58429 = n35672 & n71586;
  assign n58414 = n35197 | n35199;
  assign n58430 = n35672 & n58414;
  assign n58431 = (n71320 & n58429) | (n71320 & n58430) | (n58429 & n58430);
  assign n58432 = n35672 | n71586;
  assign n58433 = n35672 | n58414;
  assign n58434 = (n71320 & n58432) | (n71320 & n58433) | (n58432 & n58433);
  assign n35675 = ~n58431 & n58434;
  assign n35676 = x173 & x183;
  assign n35677 = n35675 & n35676;
  assign n35678 = n35675 | n35676;
  assign n35679 = ~n35677 & n35678;
  assign n35680 = n71574 & n35679;
  assign n35681 = n71574 | n35679;
  assign n35682 = ~n35680 & n35681;
  assign n35683 = x172 & x184;
  assign n35684 = n35682 & n35683;
  assign n35685 = n35682 | n35683;
  assign n35686 = ~n35684 & n35685;
  assign n58435 = n35211 & n35686;
  assign n71587 = (n35686 & n58191) | (n35686 & n58435) | (n58191 & n58435);
  assign n71588 = (n35686 & n58192) | (n35686 & n58435) | (n58192 & n58435);
  assign n71589 = (n57650 & n71587) | (n57650 & n71588) | (n71587 & n71588);
  assign n58437 = n35211 | n35686;
  assign n71590 = n58191 | n58437;
  assign n71591 = n58192 | n58437;
  assign n71592 = (n57650 & n71590) | (n57650 & n71591) | (n71590 & n71591);
  assign n35689 = ~n71589 & n71592;
  assign n35690 = x171 & x185;
  assign n35691 = n35689 & n35690;
  assign n35692 = n35689 | n35690;
  assign n35693 = ~n35691 & n35692;
  assign n58407 = n35218 | n58197;
  assign n71593 = n35693 & n58407;
  assign n71570 = n34737 | n35218;
  assign n71571 = (n35218 & n35220) | (n35218 & n71570) | (n35220 & n71570);
  assign n71594 = n35693 & n71571;
  assign n71595 = (n71270 & n71593) | (n71270 & n71594) | (n71593 & n71594);
  assign n71596 = n35693 | n58407;
  assign n71597 = n35693 | n71571;
  assign n71598 = (n71270 & n71596) | (n71270 & n71597) | (n71596 & n71597);
  assign n35696 = ~n71595 & n71598;
  assign n35697 = x170 & x186;
  assign n35698 = n35696 & n35697;
  assign n35699 = n35696 | n35697;
  assign n35700 = ~n35698 & n35699;
  assign n58405 = n35225 | n35227;
  assign n58439 = n35700 & n58405;
  assign n58440 = n35225 & n35700;
  assign n71599 = (n58145 & n58439) | (n58145 & n58440) | (n58439 & n58440);
  assign n71600 = (n58439 & n58440) | (n58439 & n71410) | (n58440 & n71410);
  assign n71601 = (n71103 & n71599) | (n71103 & n71600) | (n71599 & n71600);
  assign n58442 = n35700 | n58405;
  assign n58443 = n35225 | n35700;
  assign n71602 = (n58145 & n58442) | (n58145 & n58443) | (n58442 & n58443);
  assign n71603 = (n58442 & n58443) | (n58442 & n71410) | (n58443 & n71410);
  assign n71604 = (n71103 & n71602) | (n71103 & n71603) | (n71602 & n71603);
  assign n35703 = ~n71601 & n71604;
  assign n35704 = x169 & x187;
  assign n35705 = n35703 & n35704;
  assign n35706 = n35703 | n35704;
  assign n35707 = ~n35705 & n35706;
  assign n35708 = n71569 & n35707;
  assign n35709 = n71569 | n35707;
  assign n35710 = ~n35708 & n35709;
  assign n35711 = x168 & x188;
  assign n35712 = n35710 & n35711;
  assign n35713 = n35710 | n35711;
  assign n35714 = ~n35712 & n35713;
  assign n58400 = n35239 | n35241;
  assign n58445 = n35714 & n58400;
  assign n58446 = n35239 & n35714;
  assign n58447 = (n71408 & n58445) | (n71408 & n58446) | (n58445 & n58446);
  assign n58448 = n35714 | n58400;
  assign n58449 = n35239 | n35714;
  assign n58450 = (n71408 & n58448) | (n71408 & n58449) | (n58448 & n58449);
  assign n35717 = ~n58447 & n58450;
  assign n35718 = x167 & x189;
  assign n35719 = n35717 & n35718;
  assign n35720 = n35717 | n35718;
  assign n35721 = ~n35719 & n35720;
  assign n35722 = n58399 & n35721;
  assign n35723 = n58399 | n35721;
  assign n35724 = ~n35722 & n35723;
  assign n35725 = x166 & x190;
  assign n35726 = n35724 & n35725;
  assign n35727 = n35724 | n35725;
  assign n35728 = ~n35726 & n35727;
  assign n35729 = n71560 & n35728;
  assign n35730 = n71560 | n35728;
  assign n35731 = ~n35729 & n35730;
  assign n35732 = x165 & x191;
  assign n35733 = n35731 & n35732;
  assign n35734 = n35731 | n35732;
  assign n35735 = ~n35733 & n35734;
  assign n58392 = n35260 | n35262;
  assign n58451 = n35735 & n58392;
  assign n58452 = n35260 & n35735;
  assign n58453 = (n58136 & n58451) | (n58136 & n58452) | (n58451 & n58452);
  assign n58454 = n35735 | n58392;
  assign n58455 = n35260 | n35735;
  assign n58456 = (n58136 & n58454) | (n58136 & n58455) | (n58454 & n58455);
  assign n35738 = ~n58453 & n58456;
  assign n35739 = x164 & x192;
  assign n35740 = n35738 & n35739;
  assign n35741 = n35738 | n35739;
  assign n35742 = ~n35740 & n35741;
  assign n58457 = n35267 & n35742;
  assign n58458 = (n35742 & n58221) | (n35742 & n58457) | (n58221 & n58457);
  assign n58459 = n35267 | n35742;
  assign n58460 = n58221 | n58459;
  assign n35745 = ~n58458 & n58460;
  assign n35746 = x163 & x193;
  assign n35747 = n35745 & n35746;
  assign n35748 = n35745 | n35746;
  assign n35749 = ~n35747 & n35748;
  assign n35750 = n71555 & n35749;
  assign n35751 = n71555 | n35749;
  assign n35752 = ~n35750 & n35751;
  assign n35753 = x162 & x194;
  assign n35754 = n35752 & n35753;
  assign n35755 = n35752 | n35753;
  assign n35756 = ~n35754 & n35755;
  assign n58387 = n35281 | n35283;
  assign n58461 = n35756 & n58387;
  assign n58462 = n35281 & n35756;
  assign n58463 = (n58131 & n58461) | (n58131 & n58462) | (n58461 & n58462);
  assign n58464 = n35756 | n58387;
  assign n58465 = n35281 | n35756;
  assign n58466 = (n58131 & n58464) | (n58131 & n58465) | (n58464 & n58465);
  assign n35759 = ~n58463 & n58466;
  assign n35760 = x161 & x195;
  assign n35761 = n35759 & n35760;
  assign n35762 = n35759 | n35760;
  assign n35763 = ~n35761 & n35762;
  assign n58467 = n35288 & n35763;
  assign n58468 = (n35763 & n58231) | (n35763 & n58467) | (n58231 & n58467);
  assign n58469 = n35288 | n35763;
  assign n58470 = n58231 | n58469;
  assign n35766 = ~n58468 & n58470;
  assign n35767 = x160 & x196;
  assign n35768 = n35766 & n35767;
  assign n35769 = n35766 | n35767;
  assign n35770 = ~n35768 & n35769;
  assign n35771 = n71550 & n35770;
  assign n35772 = n71550 | n35770;
  assign n35773 = ~n35771 & n35772;
  assign n35774 = x159 & x197;
  assign n35775 = n35773 & n35774;
  assign n35776 = n35773 | n35774;
  assign n35777 = ~n35775 & n35776;
  assign n58382 = n35302 | n35304;
  assign n58471 = n35777 & n58382;
  assign n58472 = n35302 & n35777;
  assign n58473 = (n58126 & n58471) | (n58126 & n58472) | (n58471 & n58472);
  assign n58474 = n35777 | n58382;
  assign n58475 = n35302 | n35777;
  assign n58476 = (n58126 & n58474) | (n58126 & n58475) | (n58474 & n58475);
  assign n35780 = ~n58473 & n58476;
  assign n35781 = x158 & x198;
  assign n35782 = n35780 & n35781;
  assign n35783 = n35780 | n35781;
  assign n35784 = ~n35782 & n35783;
  assign n58477 = n35309 & n35784;
  assign n58478 = (n35784 & n58241) | (n35784 & n58477) | (n58241 & n58477);
  assign n58479 = n35309 | n35784;
  assign n58480 = n58241 | n58479;
  assign n35787 = ~n58478 & n58480;
  assign n35788 = x157 & x199;
  assign n35789 = n35787 & n35788;
  assign n35790 = n35787 | n35788;
  assign n35791 = ~n35789 & n35790;
  assign n35792 = n71545 & n35791;
  assign n35793 = n71545 | n35791;
  assign n35794 = ~n35792 & n35793;
  assign n35795 = x156 & x200;
  assign n35796 = n35794 & n35795;
  assign n35797 = n35794 | n35795;
  assign n35798 = ~n35796 & n35797;
  assign n58377 = n35323 | n35325;
  assign n58481 = n35798 & n58377;
  assign n58482 = n35323 & n35798;
  assign n58483 = (n71395 & n58481) | (n71395 & n58482) | (n58481 & n58482);
  assign n58484 = n35798 | n58377;
  assign n58485 = n35323 | n35798;
  assign n58486 = (n71395 & n58484) | (n71395 & n58485) | (n58484 & n58485);
  assign n35801 = ~n58483 & n58486;
  assign n35802 = x155 & x201;
  assign n35803 = n35801 & n35802;
  assign n35804 = n35801 | n35802;
  assign n35805 = ~n35803 & n35804;
  assign n58487 = n35330 & n35805;
  assign n71605 = (n35805 & n58250) | (n35805 & n58487) | (n58250 & n58487);
  assign n71606 = (n35805 & n58249) | (n35805 & n58487) | (n58249 & n58487);
  assign n71607 = (n71241 & n71605) | (n71241 & n71606) | (n71605 & n71606);
  assign n58489 = n35330 | n35805;
  assign n71608 = n58250 | n58489;
  assign n71609 = n58249 | n58489;
  assign n71610 = (n71241 & n71608) | (n71241 & n71609) | (n71608 & n71609);
  assign n35808 = ~n71607 & n71610;
  assign n35809 = x154 & x202;
  assign n35810 = n35808 & n35809;
  assign n35811 = n35808 | n35809;
  assign n35812 = ~n35810 & n35811;
  assign n35813 = n71540 & n35812;
  assign n35814 = n71540 | n35812;
  assign n35815 = ~n35813 & n35814;
  assign n35816 = x153 & x203;
  assign n35817 = n35815 & n35816;
  assign n35818 = n35815 | n35816;
  assign n35819 = ~n35817 & n35818;
  assign n58372 = n35344 | n35346;
  assign n58491 = n35819 & n58372;
  assign n58492 = n35344 & n35819;
  assign n58493 = (n71390 & n58491) | (n71390 & n58492) | (n58491 & n58492);
  assign n58494 = n35819 | n58372;
  assign n58495 = n35344 | n35819;
  assign n58496 = (n71390 & n58494) | (n71390 & n58495) | (n58494 & n58495);
  assign n35822 = ~n58493 & n58496;
  assign n35823 = x152 & x204;
  assign n35824 = n35822 & n35823;
  assign n35825 = n35822 | n35823;
  assign n35826 = ~n35824 & n35825;
  assign n58497 = n35351 & n35826;
  assign n71611 = (n35826 & n58260) | (n35826 & n58497) | (n58260 & n58497);
  assign n71612 = (n35826 & n58259) | (n35826 & n58497) | (n58259 & n58497);
  assign n71613 = (n57868 & n71611) | (n57868 & n71612) | (n71611 & n71612);
  assign n58499 = n35351 | n35826;
  assign n71614 = n58260 | n58499;
  assign n71615 = n58259 | n58499;
  assign n71616 = (n57868 & n71614) | (n57868 & n71615) | (n71614 & n71615);
  assign n35829 = ~n71613 & n71616;
  assign n35830 = x151 & x205;
  assign n35831 = n35829 & n35830;
  assign n35832 = n35829 | n35830;
  assign n35833 = ~n35831 & n35832;
  assign n58370 = n35358 | n35360;
  assign n71617 = n35833 & n58370;
  assign n71534 = n34877 | n35358;
  assign n71535 = (n35358 & n35360) | (n35358 & n71534) | (n35360 & n71534);
  assign n71618 = n35833 & n71535;
  assign n71619 = (n71368 & n71617) | (n71368 & n71618) | (n71617 & n71618);
  assign n71620 = n35833 | n58370;
  assign n71621 = n35833 | n71535;
  assign n71622 = (n71368 & n71620) | (n71368 & n71621) | (n71620 & n71621);
  assign n35836 = ~n71619 & n71622;
  assign n35837 = x150 & x206;
  assign n35838 = n35836 & n35837;
  assign n35839 = n35836 | n35837;
  assign n35840 = ~n35838 & n35839;
  assign n58501 = n35365 & n35840;
  assign n71623 = (n35840 & n58269) | (n35840 & n58501) | (n58269 & n58501);
  assign n71624 = (n35367 & n35840) | (n35367 & n58501) | (n35840 & n58501);
  assign n71625 = (n58017 & n71623) | (n58017 & n71624) | (n71623 & n71624);
  assign n58503 = n35365 | n35840;
  assign n71626 = n58269 | n58503;
  assign n71627 = n35367 | n58503;
  assign n71628 = (n58017 & n71626) | (n58017 & n71627) | (n71626 & n71627);
  assign n35843 = ~n71625 & n71628;
  assign n35844 = x149 & x207;
  assign n35845 = n35843 & n35844;
  assign n35846 = n35843 | n35844;
  assign n35847 = ~n35845 & n35846;
  assign n58505 = n35372 & n35847;
  assign n58506 = (n35847 & n58274) | (n35847 & n58505) | (n58274 & n58505);
  assign n58507 = n35372 | n35847;
  assign n58508 = n58274 | n58507;
  assign n35850 = ~n58506 & n58508;
  assign n35851 = x148 & x208;
  assign n35852 = n35850 & n35851;
  assign n35853 = n35850 | n35851;
  assign n35854 = ~n35852 & n35853;
  assign n58509 = n35379 & n35854;
  assign n58510 = (n35854 & n58278) | (n35854 & n58509) | (n58278 & n58509);
  assign n58511 = n35379 | n35854;
  assign n58512 = n58278 | n58511;
  assign n35857 = ~n58510 & n58512;
  assign n35858 = x147 & x209;
  assign n35859 = n35857 & n35858;
  assign n35860 = n35857 | n35858;
  assign n35861 = ~n35859 & n35860;
  assign n58513 = n35386 & n35861;
  assign n58514 = (n35861 & n58282) | (n35861 & n58513) | (n58282 & n58513);
  assign n58515 = n35386 | n35861;
  assign n58516 = n58282 | n58515;
  assign n35864 = ~n58514 & n58516;
  assign n35865 = x146 & x210;
  assign n35866 = n35864 & n35865;
  assign n35867 = n35864 | n35865;
  assign n35868 = ~n35866 & n35867;
  assign n58517 = n35393 & n35868;
  assign n58518 = (n35868 & n58286) | (n35868 & n58517) | (n58286 & n58517);
  assign n58519 = n35393 | n35868;
  assign n58520 = n58286 | n58519;
  assign n35871 = ~n58518 & n58520;
  assign n35872 = x145 & x211;
  assign n35873 = n35871 & n35872;
  assign n35874 = n35871 | n35872;
  assign n35875 = ~n35873 & n35874;
  assign n58521 = n35400 & n35875;
  assign n58522 = (n35875 & n58290) | (n35875 & n58521) | (n58290 & n58521);
  assign n58523 = n35400 | n35875;
  assign n58524 = n58290 | n58523;
  assign n35878 = ~n58522 & n58524;
  assign n35879 = x144 & x212;
  assign n35880 = n35878 & n35879;
  assign n35881 = n35878 | n35879;
  assign n35882 = ~n35880 & n35881;
  assign n58525 = n35407 & n35882;
  assign n58526 = (n35882 & n58294) | (n35882 & n58525) | (n58294 & n58525);
  assign n58527 = n35407 | n35882;
  assign n58528 = n58294 | n58527;
  assign n35885 = ~n58526 & n58528;
  assign n35886 = x143 & x213;
  assign n35887 = n35885 & n35886;
  assign n35888 = n35885 | n35886;
  assign n35889 = ~n35887 & n35888;
  assign n58529 = n35414 & n35889;
  assign n58530 = (n35889 & n58298) | (n35889 & n58529) | (n58298 & n58529);
  assign n58531 = n35414 | n35889;
  assign n58532 = n58298 | n58531;
  assign n35892 = ~n58530 & n58532;
  assign n35893 = x142 & x214;
  assign n35894 = n35892 & n35893;
  assign n35895 = n35892 | n35893;
  assign n35896 = ~n35894 & n35895;
  assign n58533 = n35421 & n35896;
  assign n58534 = (n35896 & n58302) | (n35896 & n58533) | (n58302 & n58533);
  assign n58535 = n35421 | n35896;
  assign n58536 = n58302 | n58535;
  assign n35899 = ~n58534 & n58536;
  assign n35900 = x141 & x215;
  assign n35901 = n35899 & n35900;
  assign n35902 = n35899 | n35900;
  assign n35903 = ~n35901 & n35902;
  assign n58537 = n35428 & n35903;
  assign n58538 = (n35903 & n58306) | (n35903 & n58537) | (n58306 & n58537);
  assign n58539 = n35428 | n35903;
  assign n58540 = n58306 | n58539;
  assign n35906 = ~n58538 & n58540;
  assign n35907 = x140 & x216;
  assign n35908 = n35906 & n35907;
  assign n35909 = n35906 | n35907;
  assign n35910 = ~n35908 & n35909;
  assign n58541 = n35435 & n35910;
  assign n58542 = (n35910 & n58310) | (n35910 & n58541) | (n58310 & n58541);
  assign n58543 = n35435 | n35910;
  assign n58544 = n58310 | n58543;
  assign n35913 = ~n58542 & n58544;
  assign n35914 = x139 & x217;
  assign n35915 = n35913 & n35914;
  assign n35916 = n35913 | n35914;
  assign n35917 = ~n35915 & n35916;
  assign n58545 = n35442 & n35917;
  assign n58546 = (n35917 & n58314) | (n35917 & n58545) | (n58314 & n58545);
  assign n58547 = n35442 | n35917;
  assign n58548 = n58314 | n58547;
  assign n35920 = ~n58546 & n58548;
  assign n35921 = x138 & x218;
  assign n35922 = n35920 & n35921;
  assign n35923 = n35920 | n35921;
  assign n35924 = ~n35922 & n35923;
  assign n58549 = n35449 & n35924;
  assign n58550 = (n35924 & n58318) | (n35924 & n58549) | (n58318 & n58549);
  assign n58551 = n35449 | n35924;
  assign n58552 = n58318 | n58551;
  assign n35927 = ~n58550 & n58552;
  assign n35928 = x137 & x219;
  assign n35929 = n35927 & n35928;
  assign n35930 = n35927 | n35928;
  assign n35931 = ~n35929 & n35930;
  assign n58553 = n35456 & n35931;
  assign n58554 = (n35931 & n58322) | (n35931 & n58553) | (n58322 & n58553);
  assign n58555 = n35456 | n35931;
  assign n58556 = n58322 | n58555;
  assign n35934 = ~n58554 & n58556;
  assign n35935 = x136 & x220;
  assign n35936 = n35934 & n35935;
  assign n35937 = n35934 | n35935;
  assign n35938 = ~n35936 & n35937;
  assign n58557 = n35463 & n35938;
  assign n58558 = (n35938 & n58326) | (n35938 & n58557) | (n58326 & n58557);
  assign n58559 = n35463 | n35938;
  assign n58560 = n58326 | n58559;
  assign n35941 = ~n58558 & n58560;
  assign n35942 = x135 & x221;
  assign n35943 = n35941 & n35942;
  assign n35944 = n35941 | n35942;
  assign n35945 = ~n35943 & n35944;
  assign n58561 = n35470 & n35945;
  assign n58562 = (n35945 & n58330) | (n35945 & n58561) | (n58330 & n58561);
  assign n58563 = n35470 | n35945;
  assign n58564 = n58330 | n58563;
  assign n35948 = ~n58562 & n58564;
  assign n35949 = x134 & x222;
  assign n35950 = n35948 & n35949;
  assign n35951 = n35948 | n35949;
  assign n35952 = ~n35950 & n35951;
  assign n58565 = n35477 & n35952;
  assign n58566 = (n35952 & n58334) | (n35952 & n58565) | (n58334 & n58565);
  assign n58567 = n35477 | n35952;
  assign n58568 = n58334 | n58567;
  assign n35955 = ~n58566 & n58568;
  assign n35956 = x133 & x223;
  assign n35957 = n35955 & n35956;
  assign n35958 = n35955 | n35956;
  assign n35959 = ~n35957 & n35958;
  assign n58569 = n35484 & n35959;
  assign n58570 = (n35959 & n58338) | (n35959 & n58569) | (n58338 & n58569);
  assign n58571 = n35484 | n35959;
  assign n58572 = n58338 | n58571;
  assign n35962 = ~n58570 & n58572;
  assign n35963 = x132 & x224;
  assign n35964 = n35962 & n35963;
  assign n35965 = n35962 | n35963;
  assign n35966 = ~n35964 & n35965;
  assign n58573 = n35491 & n35966;
  assign n58574 = (n35966 & n58342) | (n35966 & n58573) | (n58342 & n58573);
  assign n58575 = n35491 | n35966;
  assign n58576 = n58342 | n58575;
  assign n35969 = ~n58574 & n58576;
  assign n35970 = x131 & x225;
  assign n35971 = n35969 & n35970;
  assign n35972 = n35969 | n35970;
  assign n35973 = ~n35971 & n35972;
  assign n58577 = n35498 & n35973;
  assign n58578 = (n35973 & n58346) | (n35973 & n58577) | (n58346 & n58577);
  assign n58579 = n35498 | n35973;
  assign n58580 = n58346 | n58579;
  assign n35976 = ~n58578 & n58580;
  assign n35977 = x130 & x226;
  assign n35978 = n35976 & n35977;
  assign n35979 = n35976 | n35977;
  assign n35980 = ~n35978 & n35979;
  assign n58581 = n35505 & n35980;
  assign n58582 = (n35980 & n58351) | (n35980 & n58581) | (n58351 & n58581);
  assign n58583 = n35505 | n35980;
  assign n58584 = n58351 | n58583;
  assign n35983 = ~n58582 & n58584;
  assign n35984 = x129 & x227;
  assign n35985 = n35983 & n35984;
  assign n35986 = n35983 | n35984;
  assign n35987 = ~n35985 & n35986;
  assign n58367 = n35512 | n35514;
  assign n58585 = n35987 & n58367;
  assign n58586 = n35512 & n35987;
  assign n58587 = (n58109 & n58585) | (n58109 & n58586) | (n58585 & n58586);
  assign n58588 = n35987 | n58367;
  assign n58589 = n35512 | n35987;
  assign n58590 = (n58109 & n58588) | (n58109 & n58589) | (n58588 & n58589);
  assign n35990 = ~n58587 & n58590;
  assign n35991 = x128 & x228;
  assign n35992 = n35990 & n35991;
  assign n35993 = n35990 | n35991;
  assign n35994 = ~n35992 & n35993;
  assign n58365 = n35519 | n35521;
  assign n71629 = n35994 & n58365;
  assign n71630 = n35519 & n35994;
  assign n71631 = (n58107 & n71629) | (n58107 & n71630) | (n71629 & n71630);
  assign n71632 = n35994 | n58365;
  assign n71633 = n35519 | n35994;
  assign n71634 = (n58107 & n71632) | (n58107 & n71633) | (n71632 & n71633);
  assign n35997 = ~n71631 & n71634;
  assign n35998 = x127 & x229;
  assign n35999 = n35997 & n35998;
  assign n36000 = n35997 | n35998;
  assign n36001 = ~n35999 & n36000;
  assign n58363 = n35526 | n35528;
  assign n71635 = n36001 & n58363;
  assign n71636 = n35526 & n36001;
  assign n71637 = (n58105 & n71635) | (n58105 & n71636) | (n71635 & n71636);
  assign n71638 = n36001 | n58363;
  assign n71639 = n35526 | n36001;
  assign n71640 = (n58105 & n71638) | (n58105 & n71639) | (n71638 & n71639);
  assign n36004 = ~n71637 & n71640;
  assign n36005 = x126 & x230;
  assign n36006 = n36004 & n36005;
  assign n36007 = n36004 | n36005;
  assign n36008 = ~n36006 & n36007;
  assign n36009 = n58362 & n36008;
  assign n36010 = n58362 | n36008;
  assign n36011 = ~n36009 & n36010;
  assign n36012 = x125 & x231;
  assign n36013 = n36011 & n36012;
  assign n36014 = n36011 | n36012;
  assign n36015 = ~n36013 & n36014;
  assign n36016 = n58360 & n36015;
  assign n36017 = n58360 | n36015;
  assign n36018 = ~n36016 & n36017;
  assign n36019 = x124 & x232;
  assign n36020 = n36018 & n36019;
  assign n36021 = n36018 | n36019;
  assign n36022 = ~n36020 & n36021;
  assign n36023 = n35609 & n36022;
  assign n36024 = n35609 | n36022;
  assign n36025 = ~n36023 & n36024;
  assign n36026 = x123 & x233;
  assign n36027 = n36025 & n36026;
  assign n36028 = n36025 | n36026;
  assign n36029 = ~n36027 & n36028;
  assign n36030 = n35608 & n36029;
  assign n36031 = n35608 | n36029;
  assign n36032 = ~n36030 & n36031;
  assign n36033 = x122 & x234;
  assign n36034 = n36032 & n36033;
  assign n36035 = n36032 | n36033;
  assign n36036 = ~n36034 & n36035;
  assign n36037 = n35607 & n36036;
  assign n36038 = n35607 | n36036;
  assign n36039 = ~n36037 & n36038;
  assign n36040 = x121 & x235;
  assign n36041 = n36039 & n36040;
  assign n36042 = n36039 | n36040;
  assign n36043 = ~n36041 & n36042;
  assign n36044 = n35606 & n36043;
  assign n36045 = n35606 | n36043;
  assign n36046 = ~n36044 & n36045;
  assign n36047 = x120 & x236;
  assign n36048 = n36046 & n36047;
  assign n36049 = n36046 | n36047;
  assign n36050 = ~n36048 & n36049;
  assign n36051 = n35605 & n36050;
  assign n36052 = n35605 | n36050;
  assign n36053 = ~n36051 & n36052;
  assign n36054 = x119 & x237;
  assign n36055 = n36053 & n36054;
  assign n36056 = n36053 | n36054;
  assign n36057 = ~n36055 & n36056;
  assign n36058 = n71533 & n36057;
  assign n36059 = n71533 | n36057;
  assign n36060 = ~n36058 & n36059;
  assign n36061 = x118 & x238;
  assign n36062 = n36060 & n36061;
  assign n36063 = n36060 | n36061;
  assign n36064 = ~n36062 & n36063;
  assign n36065 = n58358 & n36064;
  assign n36066 = n58358 | n36064;
  assign n36067 = ~n36065 & n36066;
  assign n36068 = x117 & x239;
  assign n36069 = n36067 & n36068;
  assign n36070 = n36067 | n36068;
  assign n36071 = ~n36069 & n36070;
  assign n36072 = n58356 & n36071;
  assign n36073 = n58356 | n36071;
  assign n36074 = ~n36072 & n36073;
  assign n58591 = n36069 | n58356;
  assign n58592 = (n36069 & n36071) | (n36069 & n58591) | (n36071 & n58591);
  assign n58593 = n36062 | n58358;
  assign n58594 = (n36062 & n36064) | (n36062 & n58593) | (n36064 & n58593);
  assign n71641 = n36055 | n71533;
  assign n71642 = (n36055 & n36057) | (n36055 & n71641) | (n36057 & n71641);
  assign n36078 = n36048 | n36051;
  assign n36079 = n36041 | n36044;
  assign n36080 = n36034 | n36037;
  assign n36081 = n36027 | n36030;
  assign n58595 = n36020 | n36022;
  assign n58596 = (n35609 & n36020) | (n35609 & n58595) | (n36020 & n58595);
  assign n58597 = n36013 | n36015;
  assign n58598 = (n36013 & n58360) | (n36013 & n58597) | (n58360 & n58597);
  assign n58364 = (n35526 & n58105) | (n35526 & n58363) | (n58105 & n58363);
  assign n58366 = (n35519 & n58107) | (n35519 & n58365) | (n58107 & n58365);
  assign n58371 = (n71368 & n71535) | (n71368 & n58370) | (n71535 & n58370);
  assign n58608 = n35824 | n35826;
  assign n71643 = n35351 | n35824;
  assign n71644 = (n35824 & n35826) | (n35824 & n71643) | (n35826 & n71643);
  assign n71645 = (n58260 & n58608) | (n58260 & n71644) | (n58608 & n71644);
  assign n71646 = (n58259 & n58608) | (n58259 & n71644) | (n58608 & n71644);
  assign n71647 = (n57868 & n71645) | (n57868 & n71646) | (n71645 & n71646);
  assign n58613 = n35803 | n35805;
  assign n71648 = n35330 | n35803;
  assign n71649 = (n35803 & n35805) | (n35803 & n71648) | (n35805 & n71648);
  assign n71650 = (n58250 & n58613) | (n58250 & n71649) | (n58613 & n71649);
  assign n71651 = (n58249 & n58613) | (n58249 & n71649) | (n58613 & n71649);
  assign n71652 = (n71241 & n71650) | (n71241 & n71651) | (n71650 & n71651);
  assign n71661 = n35225 | n35698;
  assign n71662 = (n35698 & n35700) | (n35698 & n71661) | (n35700 & n71661);
  assign n71663 = n35698 | n35700;
  assign n71664 = (n35698 & n58405) | (n35698 & n71663) | (n58405 & n71663);
  assign n71665 = (n58145 & n71662) | (n58145 & n71664) | (n71662 & n71664);
  assign n71666 = (n71410 & n71662) | (n71410 & n71664) | (n71662 & n71664);
  assign n71667 = (n71103 & n71665) | (n71103 & n71666) | (n71665 & n71666);
  assign n36134 = x175 & x182;
  assign n71671 = n35665 | n58420;
  assign n71672 = (n58420 & n71576) | (n58420 & n71671) | (n71576 & n71671);
  assign n71673 = (n58420 & n71578) | (n58420 & n71671) | (n71578 & n71671);
  assign n71675 = (n71272 & n71672) | (n71272 & n71673) | (n71672 & n71673);
  assign n71677 = n36134 & n71675;
  assign n71674 = (n71273 & n71672) | (n71273 & n71673) | (n71672 & n71673);
  assign n71678 = n36134 & n71674;
  assign n71679 = (n70822 & n71677) | (n70822 & n71678) | (n71677 & n71678);
  assign n71680 = n36134 | n71675;
  assign n71681 = n36134 | n71674;
  assign n71682 = (n70822 & n71680) | (n70822 & n71681) | (n71680 & n71681);
  assign n36137 = ~n71679 & n71682;
  assign n71668 = n35670 | n35672;
  assign n71670 = (n35670 & n58414) | (n35670 & n71668) | (n58414 & n71668);
  assign n71683 = n36137 & n71670;
  assign n71669 = (n35670 & n71586) | (n35670 & n71668) | (n71586 & n71668);
  assign n71684 = n36137 & n71669;
  assign n71685 = (n71320 & n71683) | (n71320 & n71684) | (n71683 & n71684);
  assign n71686 = n36137 | n71670;
  assign n71687 = n36137 | n71669;
  assign n71688 = (n71320 & n71686) | (n71320 & n71687) | (n71686 & n71687);
  assign n36140 = ~n71685 & n71688;
  assign n36141 = x174 & x183;
  assign n36142 = n36140 & n36141;
  assign n36143 = n36140 | n36141;
  assign n36144 = ~n36142 & n36143;
  assign n58647 = n35677 | n35679;
  assign n58655 = n36144 & n58647;
  assign n58656 = n35677 & n36144;
  assign n58657 = (n71574 & n58655) | (n71574 & n58656) | (n58655 & n58656);
  assign n58658 = n36144 | n58647;
  assign n58659 = n35677 | n36144;
  assign n58660 = (n71574 & n58658) | (n71574 & n58659) | (n58658 & n58659);
  assign n36147 = ~n58657 & n58660;
  assign n36148 = x173 & x184;
  assign n36149 = n36147 & n36148;
  assign n36150 = n36147 | n36148;
  assign n36151 = ~n36149 & n36150;
  assign n71689 = n35211 | n35684;
  assign n71690 = (n35684 & n35686) | (n35684 & n71689) | (n35686 & n71689);
  assign n58661 = n36151 & n71690;
  assign n58645 = n35684 | n35686;
  assign n58662 = n36151 & n58645;
  assign n71691 = (n58191 & n58661) | (n58191 & n58662) | (n58661 & n58662);
  assign n71692 = (n58192 & n58661) | (n58192 & n58662) | (n58661 & n58662);
  assign n71693 = (n57650 & n71691) | (n57650 & n71692) | (n71691 & n71692);
  assign n58664 = n36151 | n71690;
  assign n58665 = n36151 | n58645;
  assign n71694 = (n58191 & n58664) | (n58191 & n58665) | (n58664 & n58665);
  assign n71695 = (n58192 & n58664) | (n58192 & n58665) | (n58664 & n58665);
  assign n71696 = (n57650 & n71694) | (n57650 & n71695) | (n71694 & n71695);
  assign n36154 = ~n71693 & n71696;
  assign n36155 = x172 & x185;
  assign n36156 = n36154 & n36155;
  assign n36157 = n36154 | n36155;
  assign n36158 = ~n36156 & n36157;
  assign n58642 = n35691 | n35693;
  assign n58667 = n36158 & n58642;
  assign n58668 = n35691 & n36158;
  assign n71697 = (n58407 & n58667) | (n58407 & n58668) | (n58667 & n58668);
  assign n71698 = (n58667 & n58668) | (n58667 & n71571) | (n58668 & n71571);
  assign n71699 = (n71270 & n71697) | (n71270 & n71698) | (n71697 & n71698);
  assign n58670 = n36158 | n58642;
  assign n58671 = n35691 | n36158;
  assign n71700 = (n58407 & n58670) | (n58407 & n58671) | (n58670 & n58671);
  assign n71701 = (n58670 & n58671) | (n58670 & n71571) | (n58671 & n71571);
  assign n71702 = (n71270 & n71700) | (n71270 & n71701) | (n71700 & n71701);
  assign n36161 = ~n71699 & n71702;
  assign n36162 = x171 & x186;
  assign n36163 = n36161 & n36162;
  assign n36164 = n36161 | n36162;
  assign n36165 = ~n36163 & n36164;
  assign n36166 = n71667 & n36165;
  assign n36167 = n71667 | n36165;
  assign n36168 = ~n36166 & n36167;
  assign n36169 = x170 & x187;
  assign n36170 = n36168 & n36169;
  assign n36171 = n36168 | n36169;
  assign n36172 = ~n36170 & n36171;
  assign n58637 = n35705 | n35707;
  assign n58673 = n36172 & n58637;
  assign n58674 = n35705 & n36172;
  assign n58675 = (n71569 & n58673) | (n71569 & n58674) | (n58673 & n58674);
  assign n58676 = n36172 | n58637;
  assign n58677 = n35705 | n36172;
  assign n58678 = (n71569 & n58676) | (n71569 & n58677) | (n58676 & n58677);
  assign n36175 = ~n58675 & n58678;
  assign n36176 = x169 & x188;
  assign n36177 = n36175 & n36176;
  assign n36178 = n36175 | n36176;
  assign n36179 = ~n36177 & n36178;
  assign n58635 = n35712 | n58445;
  assign n71703 = n36179 & n58635;
  assign n71659 = n35239 | n35712;
  assign n71660 = (n35712 & n35714) | (n35712 & n71659) | (n35714 & n71659);
  assign n71704 = n36179 & n71660;
  assign n71705 = (n71408 & n71703) | (n71408 & n71704) | (n71703 & n71704);
  assign n71706 = n36179 | n58635;
  assign n71707 = n36179 | n71660;
  assign n71708 = (n71408 & n71706) | (n71408 & n71707) | (n71706 & n71707);
  assign n36182 = ~n71705 & n71708;
  assign n36183 = x168 & x189;
  assign n36184 = n36182 & n36183;
  assign n36185 = n36182 | n36183;
  assign n36186 = ~n36184 & n36185;
  assign n58632 = n35719 | n35721;
  assign n58679 = n36186 & n58632;
  assign n58680 = n35719 & n36186;
  assign n58681 = (n58399 & n58679) | (n58399 & n58680) | (n58679 & n58680);
  assign n58682 = n36186 | n58632;
  assign n58683 = n35719 | n36186;
  assign n58684 = (n58399 & n58682) | (n58399 & n58683) | (n58682 & n58683);
  assign n36189 = ~n58681 & n58684;
  assign n36190 = x167 & x190;
  assign n36191 = n36189 & n36190;
  assign n36192 = n36189 | n36190;
  assign n36193 = ~n36191 & n36192;
  assign n58630 = n35726 | n35728;
  assign n58685 = n36193 & n58630;
  assign n58686 = n35726 & n36193;
  assign n58687 = (n71560 & n58685) | (n71560 & n58686) | (n58685 & n58686);
  assign n58688 = n36193 | n58630;
  assign n58689 = n35726 | n36193;
  assign n58690 = (n71560 & n58688) | (n71560 & n58689) | (n58688 & n58689);
  assign n36196 = ~n58687 & n58690;
  assign n36197 = x166 & x191;
  assign n36198 = n36196 & n36197;
  assign n36199 = n36196 | n36197;
  assign n36200 = ~n36198 & n36199;
  assign n58691 = n35733 & n36200;
  assign n71709 = (n36200 & n58452) | (n36200 & n58691) | (n58452 & n58691);
  assign n71710 = (n36200 & n58451) | (n36200 & n58691) | (n58451 & n58691);
  assign n71711 = (n58136 & n71709) | (n58136 & n71710) | (n71709 & n71710);
  assign n58693 = n35733 | n36200;
  assign n71712 = n58452 | n58693;
  assign n71713 = n58451 | n58693;
  assign n71714 = (n58136 & n71712) | (n58136 & n71713) | (n71712 & n71713);
  assign n36203 = ~n71711 & n71714;
  assign n36204 = x165 & x192;
  assign n36205 = n36203 & n36204;
  assign n36206 = n36203 | n36204;
  assign n36207 = ~n36205 & n36206;
  assign n58628 = n35740 | n35742;
  assign n71715 = n36207 & n58628;
  assign n71657 = n35267 | n35740;
  assign n71658 = (n35740 & n35742) | (n35740 & n71657) | (n35742 & n71657);
  assign n71716 = n36207 & n71658;
  assign n71717 = (n58221 & n71715) | (n58221 & n71716) | (n71715 & n71716);
  assign n71718 = n36207 | n58628;
  assign n71719 = n36207 | n71658;
  assign n71720 = (n58221 & n71718) | (n58221 & n71719) | (n71718 & n71719);
  assign n36210 = ~n71717 & n71720;
  assign n36211 = x164 & x193;
  assign n36212 = n36210 & n36211;
  assign n36213 = n36210 | n36211;
  assign n36214 = ~n36212 & n36213;
  assign n58625 = n35747 | n35749;
  assign n58695 = n36214 & n58625;
  assign n58696 = n35747 & n36214;
  assign n58697 = (n71555 & n58695) | (n71555 & n58696) | (n58695 & n58696);
  assign n58698 = n36214 | n58625;
  assign n58699 = n35747 | n36214;
  assign n58700 = (n71555 & n58698) | (n71555 & n58699) | (n58698 & n58699);
  assign n36217 = ~n58697 & n58700;
  assign n36218 = x163 & x194;
  assign n36219 = n36217 & n36218;
  assign n36220 = n36217 | n36218;
  assign n36221 = ~n36219 & n36220;
  assign n58701 = n35754 & n36221;
  assign n71721 = (n36221 & n58462) | (n36221 & n58701) | (n58462 & n58701);
  assign n71722 = (n36221 & n58461) | (n36221 & n58701) | (n58461 & n58701);
  assign n71723 = (n58131 & n71721) | (n58131 & n71722) | (n71721 & n71722);
  assign n58703 = n35754 | n36221;
  assign n71724 = n58462 | n58703;
  assign n71725 = n58461 | n58703;
  assign n71726 = (n58131 & n71724) | (n58131 & n71725) | (n71724 & n71725);
  assign n36224 = ~n71723 & n71726;
  assign n36225 = x162 & x195;
  assign n36226 = n36224 & n36225;
  assign n36227 = n36224 | n36225;
  assign n36228 = ~n36226 & n36227;
  assign n58623 = n35761 | n35763;
  assign n71727 = n36228 & n58623;
  assign n71655 = n35288 | n35761;
  assign n71656 = (n35761 & n35763) | (n35761 & n71655) | (n35763 & n71655);
  assign n71728 = n36228 & n71656;
  assign n71729 = (n58231 & n71727) | (n58231 & n71728) | (n71727 & n71728);
  assign n71730 = n36228 | n58623;
  assign n71731 = n36228 | n71656;
  assign n71732 = (n58231 & n71730) | (n58231 & n71731) | (n71730 & n71731);
  assign n36231 = ~n71729 & n71732;
  assign n36232 = x161 & x196;
  assign n36233 = n36231 & n36232;
  assign n36234 = n36231 | n36232;
  assign n36235 = ~n36233 & n36234;
  assign n58620 = n35768 | n35770;
  assign n58705 = n36235 & n58620;
  assign n58706 = n35768 & n36235;
  assign n58707 = (n71550 & n58705) | (n71550 & n58706) | (n58705 & n58706);
  assign n58708 = n36235 | n58620;
  assign n58709 = n35768 | n36235;
  assign n58710 = (n71550 & n58708) | (n71550 & n58709) | (n58708 & n58709);
  assign n36238 = ~n58707 & n58710;
  assign n36239 = x160 & x197;
  assign n36240 = n36238 & n36239;
  assign n36241 = n36238 | n36239;
  assign n36242 = ~n36240 & n36241;
  assign n58711 = n35775 & n36242;
  assign n71733 = (n36242 & n58472) | (n36242 & n58711) | (n58472 & n58711);
  assign n71734 = (n36242 & n58471) | (n36242 & n58711) | (n58471 & n58711);
  assign n71735 = (n58126 & n71733) | (n58126 & n71734) | (n71733 & n71734);
  assign n58713 = n35775 | n36242;
  assign n71736 = n58472 | n58713;
  assign n71737 = n58471 | n58713;
  assign n71738 = (n58126 & n71736) | (n58126 & n71737) | (n71736 & n71737);
  assign n36245 = ~n71735 & n71738;
  assign n36246 = x159 & x198;
  assign n36247 = n36245 & n36246;
  assign n36248 = n36245 | n36246;
  assign n36249 = ~n36247 & n36248;
  assign n58618 = n35782 | n35784;
  assign n71739 = n36249 & n58618;
  assign n71653 = n35309 | n35782;
  assign n71654 = (n35782 & n35784) | (n35782 & n71653) | (n35784 & n71653);
  assign n71740 = n36249 & n71654;
  assign n71741 = (n58241 & n71739) | (n58241 & n71740) | (n71739 & n71740);
  assign n71742 = n36249 | n58618;
  assign n71743 = n36249 | n71654;
  assign n71744 = (n58241 & n71742) | (n58241 & n71743) | (n71742 & n71743);
  assign n36252 = ~n71741 & n71744;
  assign n36253 = x158 & x199;
  assign n36254 = n36252 & n36253;
  assign n36255 = n36252 | n36253;
  assign n36256 = ~n36254 & n36255;
  assign n58615 = n35789 | n35791;
  assign n58715 = n36256 & n58615;
  assign n58716 = n35789 & n36256;
  assign n58717 = (n71545 & n58715) | (n71545 & n58716) | (n58715 & n58716);
  assign n58718 = n36256 | n58615;
  assign n58719 = n35789 | n36256;
  assign n58720 = (n71545 & n58718) | (n71545 & n58719) | (n58718 & n58719);
  assign n36259 = ~n58717 & n58720;
  assign n36260 = x157 & x200;
  assign n36261 = n36259 & n36260;
  assign n36262 = n36259 | n36260;
  assign n36263 = ~n36261 & n36262;
  assign n58721 = n35796 & n36263;
  assign n71745 = (n36263 & n58482) | (n36263 & n58721) | (n58482 & n58721);
  assign n71746 = (n36263 & n58481) | (n36263 & n58721) | (n58481 & n58721);
  assign n71747 = (n71395 & n71745) | (n71395 & n71746) | (n71745 & n71746);
  assign n58723 = n35796 | n36263;
  assign n71748 = n58482 | n58723;
  assign n71749 = n58481 | n58723;
  assign n71750 = (n71395 & n71748) | (n71395 & n71749) | (n71748 & n71749);
  assign n36266 = ~n71747 & n71750;
  assign n36267 = x156 & x201;
  assign n36268 = n36266 & n36267;
  assign n36269 = n36266 | n36267;
  assign n36270 = ~n36268 & n36269;
  assign n36271 = n71652 & n36270;
  assign n36272 = n71652 | n36270;
  assign n36273 = ~n36271 & n36272;
  assign n36274 = x155 & x202;
  assign n36275 = n36273 & n36274;
  assign n36276 = n36273 | n36274;
  assign n36277 = ~n36275 & n36276;
  assign n58610 = n35810 | n35812;
  assign n58725 = n36277 & n58610;
  assign n58726 = n35810 & n36277;
  assign n58727 = (n71540 & n58725) | (n71540 & n58726) | (n58725 & n58726);
  assign n58728 = n36277 | n58610;
  assign n58729 = n35810 | n36277;
  assign n58730 = (n71540 & n58728) | (n71540 & n58729) | (n58728 & n58729);
  assign n36280 = ~n58727 & n58730;
  assign n36281 = x154 & x203;
  assign n36282 = n36280 & n36281;
  assign n36283 = n36280 | n36281;
  assign n36284 = ~n36282 & n36283;
  assign n58731 = n35817 & n36284;
  assign n71751 = (n36284 & n58492) | (n36284 & n58731) | (n58492 & n58731);
  assign n71752 = (n36284 & n58491) | (n36284 & n58731) | (n58491 & n58731);
  assign n71753 = (n71390 & n71751) | (n71390 & n71752) | (n71751 & n71752);
  assign n58733 = n35817 | n36284;
  assign n71754 = n58492 | n58733;
  assign n71755 = n58491 | n58733;
  assign n71756 = (n71390 & n71754) | (n71390 & n71755) | (n71754 & n71755);
  assign n36287 = ~n71753 & n71756;
  assign n36288 = x153 & x204;
  assign n36289 = n36287 & n36288;
  assign n36290 = n36287 | n36288;
  assign n36291 = ~n36289 & n36290;
  assign n36292 = n71647 & n36291;
  assign n36293 = n71647 | n36291;
  assign n36294 = ~n36292 & n36293;
  assign n36295 = x152 & x205;
  assign n36296 = n36294 & n36295;
  assign n36297 = n36294 | n36295;
  assign n36298 = ~n36296 & n36297;
  assign n58605 = n35831 | n35833;
  assign n58735 = n36298 & n58605;
  assign n58736 = n35831 & n36298;
  assign n58737 = (n58371 & n58735) | (n58371 & n58736) | (n58735 & n58736);
  assign n58738 = n36298 | n58605;
  assign n58739 = n35831 | n36298;
  assign n58740 = (n58371 & n58738) | (n58371 & n58739) | (n58738 & n58739);
  assign n36301 = ~n58737 & n58740;
  assign n36302 = x151 & x206;
  assign n36303 = n36301 & n36302;
  assign n36304 = n36301 | n36302;
  assign n36305 = ~n36303 & n36304;
  assign n58741 = n35838 & n36305;
  assign n58742 = (n36305 & n71625) | (n36305 & n58741) | (n71625 & n58741);
  assign n58743 = n35838 | n36305;
  assign n58744 = n71625 | n58743;
  assign n36308 = ~n58742 & n58744;
  assign n36309 = x150 & x207;
  assign n36310 = n36308 & n36309;
  assign n36311 = n36308 | n36309;
  assign n36312 = ~n36310 & n36311;
  assign n58745 = n35845 & n36312;
  assign n58746 = (n36312 & n58506) | (n36312 & n58745) | (n58506 & n58745);
  assign n58747 = n35845 | n36312;
  assign n58748 = n58506 | n58747;
  assign n36315 = ~n58746 & n58748;
  assign n36316 = x149 & x208;
  assign n36317 = n36315 & n36316;
  assign n36318 = n36315 | n36316;
  assign n36319 = ~n36317 & n36318;
  assign n58749 = n35852 & n36319;
  assign n58750 = (n36319 & n58510) | (n36319 & n58749) | (n58510 & n58749);
  assign n58751 = n35852 | n36319;
  assign n58752 = n58510 | n58751;
  assign n36322 = ~n58750 & n58752;
  assign n36323 = x148 & x209;
  assign n36324 = n36322 & n36323;
  assign n36325 = n36322 | n36323;
  assign n36326 = ~n36324 & n36325;
  assign n58753 = n35859 & n36326;
  assign n58754 = (n36326 & n58514) | (n36326 & n58753) | (n58514 & n58753);
  assign n58755 = n35859 | n36326;
  assign n58756 = n58514 | n58755;
  assign n36329 = ~n58754 & n58756;
  assign n36330 = x147 & x210;
  assign n36331 = n36329 & n36330;
  assign n36332 = n36329 | n36330;
  assign n36333 = ~n36331 & n36332;
  assign n58757 = n35866 & n36333;
  assign n58758 = (n36333 & n58518) | (n36333 & n58757) | (n58518 & n58757);
  assign n58759 = n35866 | n36333;
  assign n58760 = n58518 | n58759;
  assign n36336 = ~n58758 & n58760;
  assign n36337 = x146 & x211;
  assign n36338 = n36336 & n36337;
  assign n36339 = n36336 | n36337;
  assign n36340 = ~n36338 & n36339;
  assign n58761 = n35873 & n36340;
  assign n58762 = (n36340 & n58522) | (n36340 & n58761) | (n58522 & n58761);
  assign n58763 = n35873 | n36340;
  assign n58764 = n58522 | n58763;
  assign n36343 = ~n58762 & n58764;
  assign n36344 = x145 & x212;
  assign n36345 = n36343 & n36344;
  assign n36346 = n36343 | n36344;
  assign n36347 = ~n36345 & n36346;
  assign n58765 = n35880 & n36347;
  assign n58766 = (n36347 & n58526) | (n36347 & n58765) | (n58526 & n58765);
  assign n58767 = n35880 | n36347;
  assign n58768 = n58526 | n58767;
  assign n36350 = ~n58766 & n58768;
  assign n36351 = x144 & x213;
  assign n36352 = n36350 & n36351;
  assign n36353 = n36350 | n36351;
  assign n36354 = ~n36352 & n36353;
  assign n58769 = n35887 & n36354;
  assign n58770 = (n36354 & n58530) | (n36354 & n58769) | (n58530 & n58769);
  assign n58771 = n35887 | n36354;
  assign n58772 = n58530 | n58771;
  assign n36357 = ~n58770 & n58772;
  assign n36358 = x143 & x214;
  assign n36359 = n36357 & n36358;
  assign n36360 = n36357 | n36358;
  assign n36361 = ~n36359 & n36360;
  assign n58773 = n35894 & n36361;
  assign n58774 = (n36361 & n58534) | (n36361 & n58773) | (n58534 & n58773);
  assign n58775 = n35894 | n36361;
  assign n58776 = n58534 | n58775;
  assign n36364 = ~n58774 & n58776;
  assign n36365 = x142 & x215;
  assign n36366 = n36364 & n36365;
  assign n36367 = n36364 | n36365;
  assign n36368 = ~n36366 & n36367;
  assign n58777 = n35901 & n36368;
  assign n58778 = (n36368 & n58538) | (n36368 & n58777) | (n58538 & n58777);
  assign n58779 = n35901 | n36368;
  assign n58780 = n58538 | n58779;
  assign n36371 = ~n58778 & n58780;
  assign n36372 = x141 & x216;
  assign n36373 = n36371 & n36372;
  assign n36374 = n36371 | n36372;
  assign n36375 = ~n36373 & n36374;
  assign n58781 = n35908 & n36375;
  assign n58782 = (n36375 & n58542) | (n36375 & n58781) | (n58542 & n58781);
  assign n58783 = n35908 | n36375;
  assign n58784 = n58542 | n58783;
  assign n36378 = ~n58782 & n58784;
  assign n36379 = x140 & x217;
  assign n36380 = n36378 & n36379;
  assign n36381 = n36378 | n36379;
  assign n36382 = ~n36380 & n36381;
  assign n58785 = n35915 & n36382;
  assign n58786 = (n36382 & n58546) | (n36382 & n58785) | (n58546 & n58785);
  assign n58787 = n35915 | n36382;
  assign n58788 = n58546 | n58787;
  assign n36385 = ~n58786 & n58788;
  assign n36386 = x139 & x218;
  assign n36387 = n36385 & n36386;
  assign n36388 = n36385 | n36386;
  assign n36389 = ~n36387 & n36388;
  assign n58789 = n35922 & n36389;
  assign n58790 = (n36389 & n58550) | (n36389 & n58789) | (n58550 & n58789);
  assign n58791 = n35922 | n36389;
  assign n58792 = n58550 | n58791;
  assign n36392 = ~n58790 & n58792;
  assign n36393 = x138 & x219;
  assign n36394 = n36392 & n36393;
  assign n36395 = n36392 | n36393;
  assign n36396 = ~n36394 & n36395;
  assign n58793 = n35929 & n36396;
  assign n58794 = (n36396 & n58554) | (n36396 & n58793) | (n58554 & n58793);
  assign n58795 = n35929 | n36396;
  assign n58796 = n58554 | n58795;
  assign n36399 = ~n58794 & n58796;
  assign n36400 = x137 & x220;
  assign n36401 = n36399 & n36400;
  assign n36402 = n36399 | n36400;
  assign n36403 = ~n36401 & n36402;
  assign n58797 = n35936 & n36403;
  assign n58798 = (n36403 & n58558) | (n36403 & n58797) | (n58558 & n58797);
  assign n58799 = n35936 | n36403;
  assign n58800 = n58558 | n58799;
  assign n36406 = ~n58798 & n58800;
  assign n36407 = x136 & x221;
  assign n36408 = n36406 & n36407;
  assign n36409 = n36406 | n36407;
  assign n36410 = ~n36408 & n36409;
  assign n58801 = n35943 & n36410;
  assign n58802 = (n36410 & n58562) | (n36410 & n58801) | (n58562 & n58801);
  assign n58803 = n35943 | n36410;
  assign n58804 = n58562 | n58803;
  assign n36413 = ~n58802 & n58804;
  assign n36414 = x135 & x222;
  assign n36415 = n36413 & n36414;
  assign n36416 = n36413 | n36414;
  assign n36417 = ~n36415 & n36416;
  assign n58805 = n35950 & n36417;
  assign n58806 = (n36417 & n58566) | (n36417 & n58805) | (n58566 & n58805);
  assign n58807 = n35950 | n36417;
  assign n58808 = n58566 | n58807;
  assign n36420 = ~n58806 & n58808;
  assign n36421 = x134 & x223;
  assign n36422 = n36420 & n36421;
  assign n36423 = n36420 | n36421;
  assign n36424 = ~n36422 & n36423;
  assign n58809 = n35957 & n36424;
  assign n58810 = (n36424 & n58570) | (n36424 & n58809) | (n58570 & n58809);
  assign n58811 = n35957 | n36424;
  assign n58812 = n58570 | n58811;
  assign n36427 = ~n58810 & n58812;
  assign n36428 = x133 & x224;
  assign n36429 = n36427 & n36428;
  assign n36430 = n36427 | n36428;
  assign n36431 = ~n36429 & n36430;
  assign n58813 = n35964 & n36431;
  assign n58814 = (n36431 & n58574) | (n36431 & n58813) | (n58574 & n58813);
  assign n58815 = n35964 | n36431;
  assign n58816 = n58574 | n58815;
  assign n36434 = ~n58814 & n58816;
  assign n36435 = x132 & x225;
  assign n36436 = n36434 & n36435;
  assign n36437 = n36434 | n36435;
  assign n36438 = ~n36436 & n36437;
  assign n58817 = n35971 & n36438;
  assign n58818 = (n36438 & n58578) | (n36438 & n58817) | (n58578 & n58817);
  assign n58819 = n35971 | n36438;
  assign n58820 = n58578 | n58819;
  assign n36441 = ~n58818 & n58820;
  assign n36442 = x131 & x226;
  assign n36443 = n36441 & n36442;
  assign n36444 = n36441 | n36442;
  assign n36445 = ~n36443 & n36444;
  assign n58821 = n35978 & n36445;
  assign n58822 = (n36445 & n58582) | (n36445 & n58821) | (n58582 & n58821);
  assign n58823 = n35978 | n36445;
  assign n58824 = n58582 | n58823;
  assign n36448 = ~n58822 & n58824;
  assign n36449 = x130 & x227;
  assign n36450 = n36448 & n36449;
  assign n36451 = n36448 | n36449;
  assign n36452 = ~n36450 & n36451;
  assign n58825 = n35985 & n36452;
  assign n58826 = (n36452 & n58587) | (n36452 & n58825) | (n58587 & n58825);
  assign n58827 = n35985 | n36452;
  assign n58828 = n58587 | n58827;
  assign n36455 = ~n58826 & n58828;
  assign n36456 = x129 & x228;
  assign n36457 = n36455 & n36456;
  assign n36458 = n36455 | n36456;
  assign n36459 = ~n36457 & n36458;
  assign n58603 = n35992 | n35994;
  assign n58829 = n36459 & n58603;
  assign n58830 = n35992 & n36459;
  assign n58831 = (n58366 & n58829) | (n58366 & n58830) | (n58829 & n58830);
  assign n58832 = n36459 | n58603;
  assign n58833 = n35992 | n36459;
  assign n58834 = (n58366 & n58832) | (n58366 & n58833) | (n58832 & n58833);
  assign n36462 = ~n58831 & n58834;
  assign n36463 = x128 & x229;
  assign n36464 = n36462 & n36463;
  assign n36465 = n36462 | n36463;
  assign n36466 = ~n36464 & n36465;
  assign n58601 = n35999 | n36001;
  assign n71757 = n36466 & n58601;
  assign n71758 = n35999 & n36466;
  assign n71759 = (n58364 & n71757) | (n58364 & n71758) | (n71757 & n71758);
  assign n71760 = n36466 | n58601;
  assign n71761 = n35999 | n36466;
  assign n71762 = (n58364 & n71760) | (n58364 & n71761) | (n71760 & n71761);
  assign n36469 = ~n71759 & n71762;
  assign n36470 = x127 & x230;
  assign n36471 = n36469 & n36470;
  assign n36472 = n36469 | n36470;
  assign n36473 = ~n36471 & n36472;
  assign n58599 = n36006 | n36008;
  assign n71763 = n36473 & n58599;
  assign n71764 = n36006 & n36473;
  assign n71765 = (n58362 & n71763) | (n58362 & n71764) | (n71763 & n71764);
  assign n71766 = n36473 | n58599;
  assign n71767 = n36006 | n36473;
  assign n71768 = (n58362 & n71766) | (n58362 & n71767) | (n71766 & n71767);
  assign n36476 = ~n71765 & n71768;
  assign n36477 = x126 & x231;
  assign n36478 = n36476 & n36477;
  assign n36479 = n36476 | n36477;
  assign n36480 = ~n36478 & n36479;
  assign n36481 = n58598 & n36480;
  assign n36482 = n58598 | n36480;
  assign n36483 = ~n36481 & n36482;
  assign n36484 = x125 & x232;
  assign n36485 = n36483 & n36484;
  assign n36486 = n36483 | n36484;
  assign n36487 = ~n36485 & n36486;
  assign n36488 = n58596 & n36487;
  assign n36489 = n58596 | n36487;
  assign n36490 = ~n36488 & n36489;
  assign n36491 = x124 & x233;
  assign n36492 = n36490 & n36491;
  assign n36493 = n36490 | n36491;
  assign n36494 = ~n36492 & n36493;
  assign n36495 = n36081 & n36494;
  assign n36496 = n36081 | n36494;
  assign n36497 = ~n36495 & n36496;
  assign n36498 = x123 & x234;
  assign n36499 = n36497 & n36498;
  assign n36500 = n36497 | n36498;
  assign n36501 = ~n36499 & n36500;
  assign n36502 = n36080 & n36501;
  assign n36503 = n36080 | n36501;
  assign n36504 = ~n36502 & n36503;
  assign n36505 = x122 & x235;
  assign n36506 = n36504 & n36505;
  assign n36507 = n36504 | n36505;
  assign n36508 = ~n36506 & n36507;
  assign n36509 = n36079 & n36508;
  assign n36510 = n36079 | n36508;
  assign n36511 = ~n36509 & n36510;
  assign n36512 = x121 & x236;
  assign n36513 = n36511 & n36512;
  assign n36514 = n36511 | n36512;
  assign n36515 = ~n36513 & n36514;
  assign n36516 = n36078 & n36515;
  assign n36517 = n36078 | n36515;
  assign n36518 = ~n36516 & n36517;
  assign n36519 = x120 & x237;
  assign n36520 = n36518 & n36519;
  assign n36521 = n36518 | n36519;
  assign n36522 = ~n36520 & n36521;
  assign n36523 = n71642 & n36522;
  assign n36524 = n71642 | n36522;
  assign n36525 = ~n36523 & n36524;
  assign n36526 = x119 & x238;
  assign n36527 = n36525 & n36526;
  assign n36528 = n36525 | n36526;
  assign n36529 = ~n36527 & n36528;
  assign n36530 = n58594 & n36529;
  assign n36531 = n58594 | n36529;
  assign n36532 = ~n36530 & n36531;
  assign n36533 = x118 & x239;
  assign n36534 = n36532 & n36533;
  assign n36535 = n36532 | n36533;
  assign n36536 = ~n36534 & n36535;
  assign n36537 = n58592 & n36536;
  assign n36538 = n58592 | n36536;
  assign n36539 = ~n36537 & n36538;
  assign n58835 = n36534 | n58592;
  assign n58836 = (n36534 & n36536) | (n36534 & n58835) | (n36536 & n58835);
  assign n58837 = n36527 | n58594;
  assign n58838 = (n36527 & n36529) | (n36527 & n58837) | (n36529 & n58837);
  assign n71769 = n36520 | n71642;
  assign n71770 = (n36520 & n36522) | (n36520 & n71769) | (n36522 & n71769);
  assign n36543 = n36513 | n36516;
  assign n36544 = n36506 | n36509;
  assign n36545 = n36499 | n36502;
  assign n58839 = n36492 | n36494;
  assign n58840 = (n36081 & n36492) | (n36081 & n58839) | (n36492 & n58839);
  assign n58841 = n36485 | n36487;
  assign n58842 = (n36485 & n58596) | (n36485 & n58841) | (n58596 & n58841);
  assign n58600 = (n36006 & n58362) | (n36006 & n58599) | (n58362 & n58599);
  assign n58602 = (n35999 & n58364) | (n35999 & n58601) | (n58364 & n58601);
  assign n58855 = n36282 | n36284;
  assign n71773 = n35817 | n36282;
  assign n71774 = (n36282 & n36284) | (n36282 & n71773) | (n36284 & n71773);
  assign n71775 = (n58492 & n58855) | (n58492 & n71774) | (n58855 & n71774);
  assign n71776 = (n58491 & n58855) | (n58491 & n71774) | (n58855 & n71774);
  assign n71777 = (n71390 & n71775) | (n71390 & n71776) | (n71775 & n71776);
  assign n58860 = n36261 | n36263;
  assign n71778 = n35796 | n36261;
  assign n71779 = (n36261 & n36263) | (n36261 & n71778) | (n36263 & n71778);
  assign n71780 = (n58482 & n58860) | (n58482 & n71779) | (n58860 & n71779);
  assign n71781 = (n58481 & n58860) | (n58481 & n71779) | (n58860 & n71779);
  assign n71782 = (n71395 & n71780) | (n71395 & n71781) | (n71780 & n71781);
  assign n58619 = (n58241 & n71654) | (n58241 & n58618) | (n71654 & n58618);
  assign n58865 = n36240 | n36242;
  assign n71783 = n35775 | n36240;
  assign n71784 = (n36240 & n36242) | (n36240 & n71783) | (n36242 & n71783);
  assign n71785 = (n58472 & n58865) | (n58472 & n71784) | (n58865 & n71784);
  assign n71786 = (n58471 & n58865) | (n58471 & n71784) | (n58865 & n71784);
  assign n71787 = (n58126 & n71785) | (n58126 & n71786) | (n71785 & n71786);
  assign n58624 = (n58231 & n71656) | (n58231 & n58623) | (n71656 & n58623);
  assign n58870 = n36219 | n36221;
  assign n71788 = n35754 | n36219;
  assign n71789 = (n36219 & n36221) | (n36219 & n71788) | (n36221 & n71788);
  assign n71790 = (n58462 & n58870) | (n58462 & n71789) | (n58870 & n71789);
  assign n71791 = (n58461 & n58870) | (n58461 & n71789) | (n58870 & n71789);
  assign n71792 = (n58131 & n71790) | (n58131 & n71791) | (n71790 & n71791);
  assign n58629 = (n58221 & n71658) | (n58221 & n58628) | (n71658 & n58628);
  assign n58875 = n36198 | n36200;
  assign n71793 = n35733 | n36198;
  assign n71794 = (n36198 & n36200) | (n36198 & n71793) | (n36200 & n71793);
  assign n71795 = (n58452 & n58875) | (n58452 & n71794) | (n58875 & n71794);
  assign n71796 = (n58451 & n58875) | (n58451 & n71794) | (n58875 & n71794);
  assign n71797 = (n58136 & n71795) | (n58136 & n71796) | (n71795 & n71796);
  assign n71804 = n36156 | n36158;
  assign n71805 = (n36156 & n58642) | (n36156 & n71804) | (n58642 & n71804);
  assign n71806 = n35691 | n36156;
  assign n71807 = (n36156 & n36158) | (n36156 & n71806) | (n36158 & n71806);
  assign n71808 = (n58407 & n71805) | (n58407 & n71807) | (n71805 & n71807);
  assign n71809 = (n71571 & n71805) | (n71571 & n71807) | (n71805 & n71807);
  assign n71810 = (n71270 & n71808) | (n71270 & n71809) | (n71808 & n71809);
  assign n36598 = x175 & x183;
  assign n58896 = n71679 & n36598;
  assign n71811 = n36598 & n71679;
  assign n71812 = (n36137 & n36598) | (n36137 & n71811) | (n36598 & n71811);
  assign n71813 = (n58896 & n71670) | (n58896 & n71812) | (n71670 & n71812);
  assign n71814 = (n58896 & n71669) | (n58896 & n71812) | (n71669 & n71812);
  assign n71815 = (n71320 & n71813) | (n71320 & n71814) | (n71813 & n71814);
  assign n58899 = n71679 | n36598;
  assign n71816 = n36598 | n71679;
  assign n71817 = n36137 | n71816;
  assign n71818 = (n58899 & n71670) | (n58899 & n71817) | (n71670 & n71817);
  assign n71819 = (n58899 & n71669) | (n58899 & n71817) | (n71669 & n71817);
  assign n71820 = (n71320 & n71818) | (n71320 & n71819) | (n71818 & n71819);
  assign n36601 = ~n71815 & n71820;
  assign n71821 = n36142 | n36144;
  assign n71822 = (n36142 & n58647) | (n36142 & n71821) | (n58647 & n71821);
  assign n58901 = n36601 & n71822;
  assign n71823 = n35677 | n36142;
  assign n71824 = (n36142 & n36144) | (n36142 & n71823) | (n36144 & n71823);
  assign n58902 = n36601 & n71824;
  assign n58903 = (n71574 & n58901) | (n71574 & n58902) | (n58901 & n58902);
  assign n58904 = n36601 | n71822;
  assign n58905 = n36601 | n71824;
  assign n58906 = (n71574 & n58904) | (n71574 & n58905) | (n58904 & n58905);
  assign n36604 = ~n58903 & n58906;
  assign n36605 = x174 & x184;
  assign n36606 = n36604 & n36605;
  assign n36607 = n36604 | n36605;
  assign n36608 = ~n36606 & n36607;
  assign n58907 = n36149 & n36608;
  assign n58908 = (n36608 & n71693) | (n36608 & n58907) | (n71693 & n58907);
  assign n58909 = n36149 | n36608;
  assign n58910 = n71693 | n58909;
  assign n36611 = ~n58908 & n58910;
  assign n36612 = x173 & x185;
  assign n36613 = n36611 & n36612;
  assign n36614 = n36611 | n36612;
  assign n36615 = ~n36613 & n36614;
  assign n36616 = n71810 & n36615;
  assign n36617 = n71810 | n36615;
  assign n36618 = ~n36616 & n36617;
  assign n36619 = x172 & x186;
  assign n36620 = n36618 & n36619;
  assign n36621 = n36618 | n36619;
  assign n36622 = ~n36620 & n36621;
  assign n58885 = n36163 | n36165;
  assign n58911 = n36622 & n58885;
  assign n58912 = n36163 & n36622;
  assign n58913 = (n71667 & n58911) | (n71667 & n58912) | (n58911 & n58912);
  assign n58914 = n36622 | n58885;
  assign n58915 = n36163 | n36622;
  assign n58916 = (n71667 & n58914) | (n71667 & n58915) | (n58914 & n58915);
  assign n36625 = ~n58913 & n58916;
  assign n36626 = x171 & x187;
  assign n36627 = n36625 & n36626;
  assign n36628 = n36625 | n36626;
  assign n36629 = ~n36627 & n36628;
  assign n58883 = n36170 | n58673;
  assign n71825 = n36629 & n58883;
  assign n71802 = n35705 | n36170;
  assign n71803 = (n36170 & n36172) | (n36170 & n71802) | (n36172 & n71802);
  assign n71826 = n36629 & n71803;
  assign n71827 = (n71569 & n71825) | (n71569 & n71826) | (n71825 & n71826);
  assign n71828 = n36629 | n58883;
  assign n71829 = n36629 | n71803;
  assign n71830 = (n71569 & n71828) | (n71569 & n71829) | (n71828 & n71829);
  assign n36632 = ~n71827 & n71830;
  assign n36633 = x170 & x188;
  assign n36634 = n36632 & n36633;
  assign n36635 = n36632 | n36633;
  assign n36636 = ~n36634 & n36635;
  assign n58880 = n36177 | n36179;
  assign n58917 = n36636 & n58880;
  assign n58918 = n36177 & n36636;
  assign n71831 = (n58635 & n58917) | (n58635 & n58918) | (n58917 & n58918);
  assign n71832 = (n58917 & n58918) | (n58917 & n71660) | (n58918 & n71660);
  assign n71833 = (n71408 & n71831) | (n71408 & n71832) | (n71831 & n71832);
  assign n58920 = n36636 | n58880;
  assign n58921 = n36177 | n36636;
  assign n71834 = (n58635 & n58920) | (n58635 & n58921) | (n58920 & n58921);
  assign n71835 = (n58920 & n58921) | (n58920 & n71660) | (n58921 & n71660);
  assign n71836 = (n71408 & n71834) | (n71408 & n71835) | (n71834 & n71835);
  assign n36639 = ~n71833 & n71836;
  assign n36640 = x169 & x189;
  assign n36641 = n36639 & n36640;
  assign n36642 = n36639 | n36640;
  assign n36643 = ~n36641 & n36642;
  assign n71800 = n36184 | n36186;
  assign n71801 = (n36184 & n58632) | (n36184 & n71800) | (n58632 & n71800);
  assign n71837 = n36643 & n71801;
  assign n71798 = n35719 | n36184;
  assign n71799 = (n36184 & n36186) | (n36184 & n71798) | (n36186 & n71798);
  assign n71838 = n36643 & n71799;
  assign n71839 = (n58399 & n71837) | (n58399 & n71838) | (n71837 & n71838);
  assign n71840 = n36643 | n71801;
  assign n71841 = n36643 | n71799;
  assign n71842 = (n58399 & n71840) | (n58399 & n71841) | (n71840 & n71841);
  assign n36646 = ~n71839 & n71842;
  assign n36647 = x168 & x190;
  assign n36648 = n36646 & n36647;
  assign n36649 = n36646 | n36647;
  assign n36650 = ~n36648 & n36649;
  assign n58923 = n36191 & n36650;
  assign n58924 = (n36650 & n58687) | (n36650 & n58923) | (n58687 & n58923);
  assign n58925 = n36191 | n36650;
  assign n58926 = n58687 | n58925;
  assign n36653 = ~n58924 & n58926;
  assign n36654 = x167 & x191;
  assign n36655 = n36653 & n36654;
  assign n36656 = n36653 | n36654;
  assign n36657 = ~n36655 & n36656;
  assign n36658 = n71797 & n36657;
  assign n36659 = n71797 | n36657;
  assign n36660 = ~n36658 & n36659;
  assign n36661 = x166 & x192;
  assign n36662 = n36660 & n36661;
  assign n36663 = n36660 | n36661;
  assign n36664 = ~n36662 & n36663;
  assign n58872 = n36205 | n36207;
  assign n58927 = n36664 & n58872;
  assign n58928 = n36205 & n36664;
  assign n58929 = (n58629 & n58927) | (n58629 & n58928) | (n58927 & n58928);
  assign n58930 = n36664 | n58872;
  assign n58931 = n36205 | n36664;
  assign n58932 = (n58629 & n58930) | (n58629 & n58931) | (n58930 & n58931);
  assign n36667 = ~n58929 & n58932;
  assign n36668 = x165 & x193;
  assign n36669 = n36667 & n36668;
  assign n36670 = n36667 | n36668;
  assign n36671 = ~n36669 & n36670;
  assign n58933 = n36212 & n36671;
  assign n58934 = (n36671 & n58697) | (n36671 & n58933) | (n58697 & n58933);
  assign n58935 = n36212 | n36671;
  assign n58936 = n58697 | n58935;
  assign n36674 = ~n58934 & n58936;
  assign n36675 = x164 & x194;
  assign n36676 = n36674 & n36675;
  assign n36677 = n36674 | n36675;
  assign n36678 = ~n36676 & n36677;
  assign n36679 = n71792 & n36678;
  assign n36680 = n71792 | n36678;
  assign n36681 = ~n36679 & n36680;
  assign n36682 = x163 & x195;
  assign n36683 = n36681 & n36682;
  assign n36684 = n36681 | n36682;
  assign n36685 = ~n36683 & n36684;
  assign n58867 = n36226 | n36228;
  assign n58937 = n36685 & n58867;
  assign n58938 = n36226 & n36685;
  assign n58939 = (n58624 & n58937) | (n58624 & n58938) | (n58937 & n58938);
  assign n58940 = n36685 | n58867;
  assign n58941 = n36226 | n36685;
  assign n58942 = (n58624 & n58940) | (n58624 & n58941) | (n58940 & n58941);
  assign n36688 = ~n58939 & n58942;
  assign n36689 = x162 & x196;
  assign n36690 = n36688 & n36689;
  assign n36691 = n36688 | n36689;
  assign n36692 = ~n36690 & n36691;
  assign n58943 = n36233 & n36692;
  assign n58944 = (n36692 & n58707) | (n36692 & n58943) | (n58707 & n58943);
  assign n58945 = n36233 | n36692;
  assign n58946 = n58707 | n58945;
  assign n36695 = ~n58944 & n58946;
  assign n36696 = x161 & x197;
  assign n36697 = n36695 & n36696;
  assign n36698 = n36695 | n36696;
  assign n36699 = ~n36697 & n36698;
  assign n36700 = n71787 & n36699;
  assign n36701 = n71787 | n36699;
  assign n36702 = ~n36700 & n36701;
  assign n36703 = x160 & x198;
  assign n36704 = n36702 & n36703;
  assign n36705 = n36702 | n36703;
  assign n36706 = ~n36704 & n36705;
  assign n58862 = n36247 | n36249;
  assign n58947 = n36706 & n58862;
  assign n58948 = n36247 & n36706;
  assign n58949 = (n58619 & n58947) | (n58619 & n58948) | (n58947 & n58948);
  assign n58950 = n36706 | n58862;
  assign n58951 = n36247 | n36706;
  assign n58952 = (n58619 & n58950) | (n58619 & n58951) | (n58950 & n58951);
  assign n36709 = ~n58949 & n58952;
  assign n36710 = x159 & x199;
  assign n36711 = n36709 & n36710;
  assign n36712 = n36709 | n36710;
  assign n36713 = ~n36711 & n36712;
  assign n58953 = n36254 & n36713;
  assign n58954 = (n36713 & n58717) | (n36713 & n58953) | (n58717 & n58953);
  assign n58955 = n36254 | n36713;
  assign n58956 = n58717 | n58955;
  assign n36716 = ~n58954 & n58956;
  assign n36717 = x158 & x200;
  assign n36718 = n36716 & n36717;
  assign n36719 = n36716 | n36717;
  assign n36720 = ~n36718 & n36719;
  assign n36721 = n71782 & n36720;
  assign n36722 = n71782 | n36720;
  assign n36723 = ~n36721 & n36722;
  assign n36724 = x157 & x201;
  assign n36725 = n36723 & n36724;
  assign n36726 = n36723 | n36724;
  assign n36727 = ~n36725 & n36726;
  assign n58857 = n36268 | n36270;
  assign n58957 = n36727 & n58857;
  assign n58958 = n36268 & n36727;
  assign n58959 = (n71652 & n58957) | (n71652 & n58958) | (n58957 & n58958);
  assign n58960 = n36727 | n58857;
  assign n58961 = n36268 | n36727;
  assign n58962 = (n71652 & n58960) | (n71652 & n58961) | (n58960 & n58961);
  assign n36730 = ~n58959 & n58962;
  assign n36731 = x156 & x202;
  assign n36732 = n36730 & n36731;
  assign n36733 = n36730 | n36731;
  assign n36734 = ~n36732 & n36733;
  assign n58963 = n36275 & n36734;
  assign n71843 = (n36734 & n58726) | (n36734 & n58963) | (n58726 & n58963);
  assign n71844 = (n36734 & n58725) | (n36734 & n58963) | (n58725 & n58963);
  assign n71845 = (n71540 & n71843) | (n71540 & n71844) | (n71843 & n71844);
  assign n58965 = n36275 | n36734;
  assign n71846 = n58726 | n58965;
  assign n71847 = n58725 | n58965;
  assign n71848 = (n71540 & n71846) | (n71540 & n71847) | (n71846 & n71847);
  assign n36737 = ~n71845 & n71848;
  assign n36738 = x155 & x203;
  assign n36739 = n36737 & n36738;
  assign n36740 = n36737 | n36738;
  assign n36741 = ~n36739 & n36740;
  assign n36742 = n71777 & n36741;
  assign n36743 = n71777 | n36741;
  assign n36744 = ~n36742 & n36743;
  assign n36745 = x154 & x204;
  assign n36746 = n36744 & n36745;
  assign n36747 = n36744 | n36745;
  assign n36748 = ~n36746 & n36747;
  assign n58852 = n36289 | n36291;
  assign n58967 = n36748 & n58852;
  assign n58968 = n36289 & n36748;
  assign n58969 = (n71647 & n58967) | (n71647 & n58968) | (n58967 & n58968);
  assign n58970 = n36748 | n58852;
  assign n58971 = n36289 | n36748;
  assign n58972 = (n71647 & n58970) | (n71647 & n58971) | (n58970 & n58971);
  assign n36751 = ~n58969 & n58972;
  assign n36752 = x153 & x205;
  assign n36753 = n36751 & n36752;
  assign n36754 = n36751 | n36752;
  assign n36755 = ~n36753 & n36754;
  assign n58973 = n36296 & n36755;
  assign n71849 = (n36755 & n58736) | (n36755 & n58973) | (n58736 & n58973);
  assign n71850 = (n36755 & n58735) | (n36755 & n58973) | (n58735 & n58973);
  assign n71851 = (n58371 & n71849) | (n58371 & n71850) | (n71849 & n71850);
  assign n58975 = n36296 | n36755;
  assign n71852 = n58736 | n58975;
  assign n71853 = n58735 | n58975;
  assign n71854 = (n58371 & n71852) | (n58371 & n71853) | (n71852 & n71853);
  assign n36758 = ~n71851 & n71854;
  assign n36759 = x152 & x206;
  assign n36760 = n36758 & n36759;
  assign n36761 = n36758 | n36759;
  assign n36762 = ~n36760 & n36761;
  assign n58850 = n36303 | n36305;
  assign n71855 = n36762 & n58850;
  assign n71771 = n35838 | n36303;
  assign n71772 = (n36303 & n36305) | (n36303 & n71771) | (n36305 & n71771);
  assign n71856 = n36762 & n71772;
  assign n71857 = (n71625 & n71855) | (n71625 & n71856) | (n71855 & n71856);
  assign n71858 = n36762 | n58850;
  assign n71859 = n36762 | n71772;
  assign n71860 = (n71625 & n71858) | (n71625 & n71859) | (n71858 & n71859);
  assign n36765 = ~n71857 & n71860;
  assign n36766 = x151 & x207;
  assign n36767 = n36765 & n36766;
  assign n36768 = n36765 | n36766;
  assign n36769 = ~n36767 & n36768;
  assign n58977 = n36310 & n36769;
  assign n71861 = (n36769 & n58745) | (n36769 & n58977) | (n58745 & n58977);
  assign n71862 = (n36312 & n36769) | (n36312 & n58977) | (n36769 & n58977);
  assign n71863 = (n58506 & n71861) | (n58506 & n71862) | (n71861 & n71862);
  assign n58979 = n36310 | n36769;
  assign n71864 = n58745 | n58979;
  assign n71865 = n36312 | n58979;
  assign n71866 = (n58506 & n71864) | (n58506 & n71865) | (n71864 & n71865);
  assign n36772 = ~n71863 & n71866;
  assign n36773 = x150 & x208;
  assign n36774 = n36772 & n36773;
  assign n36775 = n36772 | n36773;
  assign n36776 = ~n36774 & n36775;
  assign n58981 = n36317 & n36776;
  assign n58982 = (n36776 & n58750) | (n36776 & n58981) | (n58750 & n58981);
  assign n58983 = n36317 | n36776;
  assign n58984 = n58750 | n58983;
  assign n36779 = ~n58982 & n58984;
  assign n36780 = x149 & x209;
  assign n36781 = n36779 & n36780;
  assign n36782 = n36779 | n36780;
  assign n36783 = ~n36781 & n36782;
  assign n58985 = n36324 & n36783;
  assign n58986 = (n36783 & n58754) | (n36783 & n58985) | (n58754 & n58985);
  assign n58987 = n36324 | n36783;
  assign n58988 = n58754 | n58987;
  assign n36786 = ~n58986 & n58988;
  assign n36787 = x148 & x210;
  assign n36788 = n36786 & n36787;
  assign n36789 = n36786 | n36787;
  assign n36790 = ~n36788 & n36789;
  assign n58989 = n36331 & n36790;
  assign n58990 = (n36790 & n58758) | (n36790 & n58989) | (n58758 & n58989);
  assign n58991 = n36331 | n36790;
  assign n58992 = n58758 | n58991;
  assign n36793 = ~n58990 & n58992;
  assign n36794 = x147 & x211;
  assign n36795 = n36793 & n36794;
  assign n36796 = n36793 | n36794;
  assign n36797 = ~n36795 & n36796;
  assign n58993 = n36338 & n36797;
  assign n58994 = (n36797 & n58762) | (n36797 & n58993) | (n58762 & n58993);
  assign n58995 = n36338 | n36797;
  assign n58996 = n58762 | n58995;
  assign n36800 = ~n58994 & n58996;
  assign n36801 = x146 & x212;
  assign n36802 = n36800 & n36801;
  assign n36803 = n36800 | n36801;
  assign n36804 = ~n36802 & n36803;
  assign n58997 = n36345 & n36804;
  assign n58998 = (n36804 & n58766) | (n36804 & n58997) | (n58766 & n58997);
  assign n58999 = n36345 | n36804;
  assign n59000 = n58766 | n58999;
  assign n36807 = ~n58998 & n59000;
  assign n36808 = x145 & x213;
  assign n36809 = n36807 & n36808;
  assign n36810 = n36807 | n36808;
  assign n36811 = ~n36809 & n36810;
  assign n59001 = n36352 & n36811;
  assign n59002 = (n36811 & n58770) | (n36811 & n59001) | (n58770 & n59001);
  assign n59003 = n36352 | n36811;
  assign n59004 = n58770 | n59003;
  assign n36814 = ~n59002 & n59004;
  assign n36815 = x144 & x214;
  assign n36816 = n36814 & n36815;
  assign n36817 = n36814 | n36815;
  assign n36818 = ~n36816 & n36817;
  assign n59005 = n36359 & n36818;
  assign n59006 = (n36818 & n58774) | (n36818 & n59005) | (n58774 & n59005);
  assign n59007 = n36359 | n36818;
  assign n59008 = n58774 | n59007;
  assign n36821 = ~n59006 & n59008;
  assign n36822 = x143 & x215;
  assign n36823 = n36821 & n36822;
  assign n36824 = n36821 | n36822;
  assign n36825 = ~n36823 & n36824;
  assign n59009 = n36366 & n36825;
  assign n59010 = (n36825 & n58778) | (n36825 & n59009) | (n58778 & n59009);
  assign n59011 = n36366 | n36825;
  assign n59012 = n58778 | n59011;
  assign n36828 = ~n59010 & n59012;
  assign n36829 = x142 & x216;
  assign n36830 = n36828 & n36829;
  assign n36831 = n36828 | n36829;
  assign n36832 = ~n36830 & n36831;
  assign n59013 = n36373 & n36832;
  assign n59014 = (n36832 & n58782) | (n36832 & n59013) | (n58782 & n59013);
  assign n59015 = n36373 | n36832;
  assign n59016 = n58782 | n59015;
  assign n36835 = ~n59014 & n59016;
  assign n36836 = x141 & x217;
  assign n36837 = n36835 & n36836;
  assign n36838 = n36835 | n36836;
  assign n36839 = ~n36837 & n36838;
  assign n59017 = n36380 & n36839;
  assign n59018 = (n36839 & n58786) | (n36839 & n59017) | (n58786 & n59017);
  assign n59019 = n36380 | n36839;
  assign n59020 = n58786 | n59019;
  assign n36842 = ~n59018 & n59020;
  assign n36843 = x140 & x218;
  assign n36844 = n36842 & n36843;
  assign n36845 = n36842 | n36843;
  assign n36846 = ~n36844 & n36845;
  assign n59021 = n36387 & n36846;
  assign n59022 = (n36846 & n58790) | (n36846 & n59021) | (n58790 & n59021);
  assign n59023 = n36387 | n36846;
  assign n59024 = n58790 | n59023;
  assign n36849 = ~n59022 & n59024;
  assign n36850 = x139 & x219;
  assign n36851 = n36849 & n36850;
  assign n36852 = n36849 | n36850;
  assign n36853 = ~n36851 & n36852;
  assign n59025 = n36394 & n36853;
  assign n59026 = (n36853 & n58794) | (n36853 & n59025) | (n58794 & n59025);
  assign n59027 = n36394 | n36853;
  assign n59028 = n58794 | n59027;
  assign n36856 = ~n59026 & n59028;
  assign n36857 = x138 & x220;
  assign n36858 = n36856 & n36857;
  assign n36859 = n36856 | n36857;
  assign n36860 = ~n36858 & n36859;
  assign n59029 = n36401 & n36860;
  assign n59030 = (n36860 & n58798) | (n36860 & n59029) | (n58798 & n59029);
  assign n59031 = n36401 | n36860;
  assign n59032 = n58798 | n59031;
  assign n36863 = ~n59030 & n59032;
  assign n36864 = x137 & x221;
  assign n36865 = n36863 & n36864;
  assign n36866 = n36863 | n36864;
  assign n36867 = ~n36865 & n36866;
  assign n59033 = n36408 & n36867;
  assign n59034 = (n36867 & n58802) | (n36867 & n59033) | (n58802 & n59033);
  assign n59035 = n36408 | n36867;
  assign n59036 = n58802 | n59035;
  assign n36870 = ~n59034 & n59036;
  assign n36871 = x136 & x222;
  assign n36872 = n36870 & n36871;
  assign n36873 = n36870 | n36871;
  assign n36874 = ~n36872 & n36873;
  assign n59037 = n36415 & n36874;
  assign n59038 = (n36874 & n58806) | (n36874 & n59037) | (n58806 & n59037);
  assign n59039 = n36415 | n36874;
  assign n59040 = n58806 | n59039;
  assign n36877 = ~n59038 & n59040;
  assign n36878 = x135 & x223;
  assign n36879 = n36877 & n36878;
  assign n36880 = n36877 | n36878;
  assign n36881 = ~n36879 & n36880;
  assign n59041 = n36422 & n36881;
  assign n59042 = (n36881 & n58810) | (n36881 & n59041) | (n58810 & n59041);
  assign n59043 = n36422 | n36881;
  assign n59044 = n58810 | n59043;
  assign n36884 = ~n59042 & n59044;
  assign n36885 = x134 & x224;
  assign n36886 = n36884 & n36885;
  assign n36887 = n36884 | n36885;
  assign n36888 = ~n36886 & n36887;
  assign n59045 = n36429 & n36888;
  assign n59046 = (n36888 & n58814) | (n36888 & n59045) | (n58814 & n59045);
  assign n59047 = n36429 | n36888;
  assign n59048 = n58814 | n59047;
  assign n36891 = ~n59046 & n59048;
  assign n36892 = x133 & x225;
  assign n36893 = n36891 & n36892;
  assign n36894 = n36891 | n36892;
  assign n36895 = ~n36893 & n36894;
  assign n59049 = n36436 & n36895;
  assign n59050 = (n36895 & n58818) | (n36895 & n59049) | (n58818 & n59049);
  assign n59051 = n36436 | n36895;
  assign n59052 = n58818 | n59051;
  assign n36898 = ~n59050 & n59052;
  assign n36899 = x132 & x226;
  assign n36900 = n36898 & n36899;
  assign n36901 = n36898 | n36899;
  assign n36902 = ~n36900 & n36901;
  assign n59053 = n36443 & n36902;
  assign n59054 = (n36902 & n58822) | (n36902 & n59053) | (n58822 & n59053);
  assign n59055 = n36443 | n36902;
  assign n59056 = n58822 | n59055;
  assign n36905 = ~n59054 & n59056;
  assign n36906 = x131 & x227;
  assign n36907 = n36905 & n36906;
  assign n36908 = n36905 | n36906;
  assign n36909 = ~n36907 & n36908;
  assign n59057 = n36450 & n36909;
  assign n59058 = (n36909 & n58826) | (n36909 & n59057) | (n58826 & n59057);
  assign n59059 = n36450 | n36909;
  assign n59060 = n58826 | n59059;
  assign n36912 = ~n59058 & n59060;
  assign n36913 = x130 & x228;
  assign n36914 = n36912 & n36913;
  assign n36915 = n36912 | n36913;
  assign n36916 = ~n36914 & n36915;
  assign n59061 = n36457 & n36916;
  assign n59062 = (n36916 & n58831) | (n36916 & n59061) | (n58831 & n59061);
  assign n59063 = n36457 | n36916;
  assign n59064 = n58831 | n59063;
  assign n36919 = ~n59062 & n59064;
  assign n36920 = x129 & x229;
  assign n36921 = n36919 & n36920;
  assign n36922 = n36919 | n36920;
  assign n36923 = ~n36921 & n36922;
  assign n58847 = n36464 | n36466;
  assign n59065 = n36923 & n58847;
  assign n59066 = n36464 & n36923;
  assign n59067 = (n58602 & n59065) | (n58602 & n59066) | (n59065 & n59066);
  assign n59068 = n36923 | n58847;
  assign n59069 = n36464 | n36923;
  assign n59070 = (n58602 & n59068) | (n58602 & n59069) | (n59068 & n59069);
  assign n36926 = ~n59067 & n59070;
  assign n36927 = x128 & x230;
  assign n36928 = n36926 & n36927;
  assign n36929 = n36926 | n36927;
  assign n36930 = ~n36928 & n36929;
  assign n58845 = n36471 | n36473;
  assign n71867 = n36930 & n58845;
  assign n71868 = n36471 & n36930;
  assign n71869 = (n58600 & n71867) | (n58600 & n71868) | (n71867 & n71868);
  assign n71870 = n36930 | n58845;
  assign n71871 = n36471 | n36930;
  assign n71872 = (n58600 & n71870) | (n58600 & n71871) | (n71870 & n71871);
  assign n36933 = ~n71869 & n71872;
  assign n36934 = x127 & x231;
  assign n36935 = n36933 & n36934;
  assign n36936 = n36933 | n36934;
  assign n36937 = ~n36935 & n36936;
  assign n58843 = n36478 | n36480;
  assign n71873 = n36937 & n58843;
  assign n71874 = n36478 & n36937;
  assign n71875 = (n58598 & n71873) | (n58598 & n71874) | (n71873 & n71874);
  assign n71876 = n36937 | n58843;
  assign n71877 = n36478 | n36937;
  assign n71878 = (n58598 & n71876) | (n58598 & n71877) | (n71876 & n71877);
  assign n36940 = ~n71875 & n71878;
  assign n36941 = x126 & x232;
  assign n36942 = n36940 & n36941;
  assign n36943 = n36940 | n36941;
  assign n36944 = ~n36942 & n36943;
  assign n36945 = n58842 & n36944;
  assign n36946 = n58842 | n36944;
  assign n36947 = ~n36945 & n36946;
  assign n36948 = x125 & x233;
  assign n36949 = n36947 & n36948;
  assign n36950 = n36947 | n36948;
  assign n36951 = ~n36949 & n36950;
  assign n36952 = n58840 & n36951;
  assign n36953 = n58840 | n36951;
  assign n36954 = ~n36952 & n36953;
  assign n36955 = x124 & x234;
  assign n36956 = n36954 & n36955;
  assign n36957 = n36954 | n36955;
  assign n36958 = ~n36956 & n36957;
  assign n36959 = n36545 & n36958;
  assign n36960 = n36545 | n36958;
  assign n36961 = ~n36959 & n36960;
  assign n36962 = x123 & x235;
  assign n36963 = n36961 & n36962;
  assign n36964 = n36961 | n36962;
  assign n36965 = ~n36963 & n36964;
  assign n36966 = n36544 & n36965;
  assign n36967 = n36544 | n36965;
  assign n36968 = ~n36966 & n36967;
  assign n36969 = x122 & x236;
  assign n36970 = n36968 & n36969;
  assign n36971 = n36968 | n36969;
  assign n36972 = ~n36970 & n36971;
  assign n36973 = n36543 & n36972;
  assign n36974 = n36543 | n36972;
  assign n36975 = ~n36973 & n36974;
  assign n36976 = x121 & x237;
  assign n36977 = n36975 & n36976;
  assign n36978 = n36975 | n36976;
  assign n36979 = ~n36977 & n36978;
  assign n36980 = n71770 & n36979;
  assign n36981 = n71770 | n36979;
  assign n36982 = ~n36980 & n36981;
  assign n36983 = x120 & x238;
  assign n36984 = n36982 & n36983;
  assign n36985 = n36982 | n36983;
  assign n36986 = ~n36984 & n36985;
  assign n36987 = n58838 & n36986;
  assign n36988 = n58838 | n36986;
  assign n36989 = ~n36987 & n36988;
  assign n36990 = x119 & x239;
  assign n36991 = n36989 & n36990;
  assign n36992 = n36989 | n36990;
  assign n36993 = ~n36991 & n36992;
  assign n36994 = n58836 & n36993;
  assign n36995 = n58836 | n36993;
  assign n36996 = ~n36994 & n36995;
  assign n59071 = n36991 | n58836;
  assign n59072 = (n36991 & n36993) | (n36991 & n59071) | (n36993 & n59071);
  assign n59073 = n36984 | n58838;
  assign n59074 = (n36984 & n36986) | (n36984 & n59073) | (n36986 & n59073);
  assign n71879 = n36977 | n71770;
  assign n71880 = (n36977 & n36979) | (n36977 & n71879) | (n36979 & n71879);
  assign n37000 = n36970 | n36973;
  assign n37001 = n36963 | n36966;
  assign n59075 = n36956 | n36958;
  assign n59076 = (n36545 & n36956) | (n36545 & n59075) | (n36956 & n59075);
  assign n59077 = n36949 | n36951;
  assign n59078 = (n36949 & n58840) | (n36949 & n59077) | (n58840 & n59077);
  assign n58844 = (n36478 & n58598) | (n36478 & n58843) | (n58598 & n58843);
  assign n58846 = (n36471 & n58600) | (n36471 & n58845) | (n58600 & n58845);
  assign n58851 = (n71625 & n71772) | (n71625 & n58850) | (n71772 & n58850);
  assign n59088 = n36753 | n36755;
  assign n71881 = n36296 | n36753;
  assign n71882 = (n36753 & n36755) | (n36753 & n71881) | (n36755 & n71881);
  assign n71883 = (n58736 & n59088) | (n58736 & n71882) | (n59088 & n71882);
  assign n71884 = (n58735 & n59088) | (n58735 & n71882) | (n59088 & n71882);
  assign n71885 = (n58371 & n71883) | (n58371 & n71884) | (n71883 & n71884);
  assign n59093 = n36732 | n36734;
  assign n71886 = n36275 | n36732;
  assign n71887 = (n36732 & n36734) | (n36732 & n71886) | (n36734 & n71886);
  assign n71888 = (n58726 & n59093) | (n58726 & n71887) | (n59093 & n71887);
  assign n71889 = (n58725 & n59093) | (n58725 & n71887) | (n59093 & n71887);
  assign n71890 = (n71540 & n71888) | (n71540 & n71889) | (n71888 & n71889);
  assign n71899 = n36177 | n36634;
  assign n71900 = (n36634 & n36636) | (n36634 & n71899) | (n36636 & n71899);
  assign n71901 = n36634 | n36636;
  assign n71902 = (n36634 & n58880) | (n36634 & n71901) | (n58880 & n71901);
  assign n71903 = (n58635 & n71900) | (n58635 & n71902) | (n71900 & n71902);
  assign n71904 = (n71660 & n71900) | (n71660 & n71902) | (n71900 & n71902);
  assign n71905 = (n71408 & n71903) | (n71408 & n71904) | (n71903 & n71904);
  assign n37054 = x175 & x184;
  assign n71908 = n37054 & n71814;
  assign n71909 = n37054 & n71813;
  assign n71910 = (n71320 & n71908) | (n71320 & n71909) | (n71908 & n71909);
  assign n71911 = (n37054 & n58901) | (n37054 & n71910) | (n58901 & n71910);
  assign n71912 = (n37054 & n58902) | (n37054 & n71910) | (n58902 & n71910);
  assign n71913 = (n71574 & n71911) | (n71574 & n71912) | (n71911 & n71912);
  assign n71914 = n37054 | n71814;
  assign n71915 = n37054 | n71813;
  assign n71916 = (n71320 & n71914) | (n71320 & n71915) | (n71914 & n71915);
  assign n71917 = n58901 | n71916;
  assign n71918 = n58902 | n71916;
  assign n71919 = (n71574 & n71917) | (n71574 & n71918) | (n71917 & n71918);
  assign n37057 = ~n71913 & n71919;
  assign n71920 = n36149 | n36606;
  assign n71921 = (n36606 & n36608) | (n36606 & n71920) | (n36608 & n71920);
  assign n59134 = n37057 & n71921;
  assign n71922 = n36606 & n37057;
  assign n71923 = (n36608 & n37057) | (n36608 & n71922) | (n37057 & n71922);
  assign n59136 = (n71693 & n59134) | (n71693 & n71923) | (n59134 & n71923);
  assign n59137 = n37057 | n71921;
  assign n71924 = n36606 | n37057;
  assign n71925 = n36608 | n71924;
  assign n59139 = (n71693 & n59137) | (n71693 & n71925) | (n59137 & n71925);
  assign n37060 = ~n59136 & n59139;
  assign n37061 = x174 & x185;
  assign n37062 = n37060 & n37061;
  assign n37063 = n37060 | n37061;
  assign n37064 = ~n37062 & n37063;
  assign n59125 = n36613 | n36615;
  assign n59140 = n37064 & n59125;
  assign n59141 = n36613 & n37064;
  assign n59142 = (n71810 & n59140) | (n71810 & n59141) | (n59140 & n59141);
  assign n59143 = n37064 | n59125;
  assign n59144 = n36613 | n37064;
  assign n59145 = (n71810 & n59143) | (n71810 & n59144) | (n59143 & n59144);
  assign n37067 = ~n59142 & n59145;
  assign n37068 = x173 & x186;
  assign n37069 = n37067 & n37068;
  assign n37070 = n37067 | n37068;
  assign n37071 = ~n37069 & n37070;
  assign n59123 = n36620 | n58911;
  assign n71926 = n37071 & n59123;
  assign n71906 = n36163 | n36620;
  assign n71907 = (n36620 & n36622) | (n36620 & n71906) | (n36622 & n71906);
  assign n71927 = n37071 & n71907;
  assign n71928 = (n71667 & n71926) | (n71667 & n71927) | (n71926 & n71927);
  assign n71929 = n37071 | n59123;
  assign n71930 = n37071 | n71907;
  assign n71931 = (n71667 & n71929) | (n71667 & n71930) | (n71929 & n71930);
  assign n37074 = ~n71928 & n71931;
  assign n37075 = x172 & x187;
  assign n37076 = n37074 & n37075;
  assign n37077 = n37074 | n37075;
  assign n37078 = ~n37076 & n37077;
  assign n59120 = n36627 | n36629;
  assign n59146 = n37078 & n59120;
  assign n59147 = n36627 & n37078;
  assign n71932 = (n58883 & n59146) | (n58883 & n59147) | (n59146 & n59147);
  assign n71933 = (n59146 & n59147) | (n59146 & n71803) | (n59147 & n71803);
  assign n71934 = (n71569 & n71932) | (n71569 & n71933) | (n71932 & n71933);
  assign n59149 = n37078 | n59120;
  assign n59150 = n36627 | n37078;
  assign n71935 = (n58883 & n59149) | (n58883 & n59150) | (n59149 & n59150);
  assign n71936 = (n59149 & n59150) | (n59149 & n71803) | (n59150 & n71803);
  assign n71937 = (n71569 & n71935) | (n71569 & n71936) | (n71935 & n71936);
  assign n37081 = ~n71934 & n71937;
  assign n37082 = x171 & x188;
  assign n37083 = n37081 & n37082;
  assign n37084 = n37081 | n37082;
  assign n37085 = ~n37083 & n37084;
  assign n37086 = n71905 & n37085;
  assign n37087 = n71905 | n37085;
  assign n37088 = ~n37086 & n37087;
  assign n37089 = x170 & x189;
  assign n37090 = n37088 & n37089;
  assign n37091 = n37088 | n37089;
  assign n37092 = ~n37090 & n37091;
  assign n59115 = n36641 | n36643;
  assign n59152 = n37092 & n59115;
  assign n59153 = n36641 & n37092;
  assign n71938 = (n59152 & n59153) | (n59152 & n71801) | (n59153 & n71801);
  assign n71939 = (n59152 & n59153) | (n59152 & n71799) | (n59153 & n71799);
  assign n71940 = (n58399 & n71938) | (n58399 & n71939) | (n71938 & n71939);
  assign n59155 = n37092 | n59115;
  assign n59156 = n36641 | n37092;
  assign n71941 = (n59155 & n59156) | (n59155 & n71801) | (n59156 & n71801);
  assign n71942 = (n59155 & n59156) | (n59155 & n71799) | (n59156 & n71799);
  assign n71943 = (n58399 & n71941) | (n58399 & n71942) | (n71941 & n71942);
  assign n37095 = ~n71940 & n71943;
  assign n37096 = x169 & x190;
  assign n37097 = n37095 & n37096;
  assign n37098 = n37095 | n37096;
  assign n37099 = ~n37097 & n37098;
  assign n59113 = n36648 | n36650;
  assign n71944 = n37099 & n59113;
  assign n71897 = n36191 | n36648;
  assign n71898 = (n36648 & n36650) | (n36648 & n71897) | (n36650 & n71897);
  assign n71945 = n37099 & n71898;
  assign n71946 = (n58687 & n71944) | (n58687 & n71945) | (n71944 & n71945);
  assign n71947 = n37099 | n59113;
  assign n71948 = n37099 | n71898;
  assign n71949 = (n58687 & n71947) | (n58687 & n71948) | (n71947 & n71948);
  assign n37102 = ~n71946 & n71949;
  assign n37103 = x168 & x191;
  assign n37104 = n37102 & n37103;
  assign n37105 = n37102 | n37103;
  assign n37106 = ~n37104 & n37105;
  assign n59110 = n36655 | n36657;
  assign n59158 = n37106 & n59110;
  assign n59159 = n36655 & n37106;
  assign n59160 = (n71797 & n59158) | (n71797 & n59159) | (n59158 & n59159);
  assign n59161 = n37106 | n59110;
  assign n59162 = n36655 | n37106;
  assign n59163 = (n71797 & n59161) | (n71797 & n59162) | (n59161 & n59162);
  assign n37109 = ~n59160 & n59163;
  assign n37110 = x167 & x192;
  assign n37111 = n37109 & n37110;
  assign n37112 = n37109 | n37110;
  assign n37113 = ~n37111 & n37112;
  assign n59164 = n36662 & n37113;
  assign n71950 = (n37113 & n58928) | (n37113 & n59164) | (n58928 & n59164);
  assign n71951 = (n37113 & n58927) | (n37113 & n59164) | (n58927 & n59164);
  assign n71952 = (n58629 & n71950) | (n58629 & n71951) | (n71950 & n71951);
  assign n59166 = n36662 | n37113;
  assign n71953 = n58928 | n59166;
  assign n71954 = n58927 | n59166;
  assign n71955 = (n58629 & n71953) | (n58629 & n71954) | (n71953 & n71954);
  assign n37116 = ~n71952 & n71955;
  assign n37117 = x166 & x193;
  assign n37118 = n37116 & n37117;
  assign n37119 = n37116 | n37117;
  assign n37120 = ~n37118 & n37119;
  assign n59108 = n36669 | n36671;
  assign n71956 = n37120 & n59108;
  assign n71895 = n36212 | n36669;
  assign n71896 = (n36669 & n36671) | (n36669 & n71895) | (n36671 & n71895);
  assign n71957 = n37120 & n71896;
  assign n71958 = (n58697 & n71956) | (n58697 & n71957) | (n71956 & n71957);
  assign n71959 = n37120 | n59108;
  assign n71960 = n37120 | n71896;
  assign n71961 = (n58697 & n71959) | (n58697 & n71960) | (n71959 & n71960);
  assign n37123 = ~n71958 & n71961;
  assign n37124 = x165 & x194;
  assign n37125 = n37123 & n37124;
  assign n37126 = n37123 | n37124;
  assign n37127 = ~n37125 & n37126;
  assign n59105 = n36676 | n36678;
  assign n59168 = n37127 & n59105;
  assign n59169 = n36676 & n37127;
  assign n59170 = (n71792 & n59168) | (n71792 & n59169) | (n59168 & n59169);
  assign n59171 = n37127 | n59105;
  assign n59172 = n36676 | n37127;
  assign n59173 = (n71792 & n59171) | (n71792 & n59172) | (n59171 & n59172);
  assign n37130 = ~n59170 & n59173;
  assign n37131 = x164 & x195;
  assign n37132 = n37130 & n37131;
  assign n37133 = n37130 | n37131;
  assign n37134 = ~n37132 & n37133;
  assign n59174 = n36683 & n37134;
  assign n71962 = (n37134 & n58938) | (n37134 & n59174) | (n58938 & n59174);
  assign n71963 = (n37134 & n58937) | (n37134 & n59174) | (n58937 & n59174);
  assign n71964 = (n58624 & n71962) | (n58624 & n71963) | (n71962 & n71963);
  assign n59176 = n36683 | n37134;
  assign n71965 = n58938 | n59176;
  assign n71966 = n58937 | n59176;
  assign n71967 = (n58624 & n71965) | (n58624 & n71966) | (n71965 & n71966);
  assign n37137 = ~n71964 & n71967;
  assign n37138 = x163 & x196;
  assign n37139 = n37137 & n37138;
  assign n37140 = n37137 | n37138;
  assign n37141 = ~n37139 & n37140;
  assign n59103 = n36690 | n36692;
  assign n71968 = n37141 & n59103;
  assign n71893 = n36233 | n36690;
  assign n71894 = (n36690 & n36692) | (n36690 & n71893) | (n36692 & n71893);
  assign n71969 = n37141 & n71894;
  assign n71970 = (n58707 & n71968) | (n58707 & n71969) | (n71968 & n71969);
  assign n71971 = n37141 | n59103;
  assign n71972 = n37141 | n71894;
  assign n71973 = (n58707 & n71971) | (n58707 & n71972) | (n71971 & n71972);
  assign n37144 = ~n71970 & n71973;
  assign n37145 = x162 & x197;
  assign n37146 = n37144 & n37145;
  assign n37147 = n37144 | n37145;
  assign n37148 = ~n37146 & n37147;
  assign n59100 = n36697 | n36699;
  assign n59178 = n37148 & n59100;
  assign n59179 = n36697 & n37148;
  assign n59180 = (n71787 & n59178) | (n71787 & n59179) | (n59178 & n59179);
  assign n59181 = n37148 | n59100;
  assign n59182 = n36697 | n37148;
  assign n59183 = (n71787 & n59181) | (n71787 & n59182) | (n59181 & n59182);
  assign n37151 = ~n59180 & n59183;
  assign n37152 = x161 & x198;
  assign n37153 = n37151 & n37152;
  assign n37154 = n37151 | n37152;
  assign n37155 = ~n37153 & n37154;
  assign n59184 = n36704 & n37155;
  assign n71974 = (n37155 & n58948) | (n37155 & n59184) | (n58948 & n59184);
  assign n71975 = (n37155 & n58947) | (n37155 & n59184) | (n58947 & n59184);
  assign n71976 = (n58619 & n71974) | (n58619 & n71975) | (n71974 & n71975);
  assign n59186 = n36704 | n37155;
  assign n71977 = n58948 | n59186;
  assign n71978 = n58947 | n59186;
  assign n71979 = (n58619 & n71977) | (n58619 & n71978) | (n71977 & n71978);
  assign n37158 = ~n71976 & n71979;
  assign n37159 = x160 & x199;
  assign n37160 = n37158 & n37159;
  assign n37161 = n37158 | n37159;
  assign n37162 = ~n37160 & n37161;
  assign n59098 = n36711 | n36713;
  assign n71980 = n37162 & n59098;
  assign n71891 = n36254 | n36711;
  assign n71892 = (n36711 & n36713) | (n36711 & n71891) | (n36713 & n71891);
  assign n71981 = n37162 & n71892;
  assign n71982 = (n58717 & n71980) | (n58717 & n71981) | (n71980 & n71981);
  assign n71983 = n37162 | n59098;
  assign n71984 = n37162 | n71892;
  assign n71985 = (n58717 & n71983) | (n58717 & n71984) | (n71983 & n71984);
  assign n37165 = ~n71982 & n71985;
  assign n37166 = x159 & x200;
  assign n37167 = n37165 & n37166;
  assign n37168 = n37165 | n37166;
  assign n37169 = ~n37167 & n37168;
  assign n59095 = n36718 | n36720;
  assign n59188 = n37169 & n59095;
  assign n59189 = n36718 & n37169;
  assign n59190 = (n71782 & n59188) | (n71782 & n59189) | (n59188 & n59189);
  assign n59191 = n37169 | n59095;
  assign n59192 = n36718 | n37169;
  assign n59193 = (n71782 & n59191) | (n71782 & n59192) | (n59191 & n59192);
  assign n37172 = ~n59190 & n59193;
  assign n37173 = x158 & x201;
  assign n37174 = n37172 & n37173;
  assign n37175 = n37172 | n37173;
  assign n37176 = ~n37174 & n37175;
  assign n59194 = n36725 & n37176;
  assign n71986 = (n37176 & n58958) | (n37176 & n59194) | (n58958 & n59194);
  assign n71987 = (n37176 & n58957) | (n37176 & n59194) | (n58957 & n59194);
  assign n71988 = (n71652 & n71986) | (n71652 & n71987) | (n71986 & n71987);
  assign n59196 = n36725 | n37176;
  assign n71989 = n58958 | n59196;
  assign n71990 = n58957 | n59196;
  assign n71991 = (n71652 & n71989) | (n71652 & n71990) | (n71989 & n71990);
  assign n37179 = ~n71988 & n71991;
  assign n37180 = x157 & x202;
  assign n37181 = n37179 & n37180;
  assign n37182 = n37179 | n37180;
  assign n37183 = ~n37181 & n37182;
  assign n37184 = n71890 & n37183;
  assign n37185 = n71890 | n37183;
  assign n37186 = ~n37184 & n37185;
  assign n37187 = x156 & x203;
  assign n37188 = n37186 & n37187;
  assign n37189 = n37186 | n37187;
  assign n37190 = ~n37188 & n37189;
  assign n59090 = n36739 | n36741;
  assign n59198 = n37190 & n59090;
  assign n59199 = n36739 & n37190;
  assign n59200 = (n71777 & n59198) | (n71777 & n59199) | (n59198 & n59199);
  assign n59201 = n37190 | n59090;
  assign n59202 = n36739 | n37190;
  assign n59203 = (n71777 & n59201) | (n71777 & n59202) | (n59201 & n59202);
  assign n37193 = ~n59200 & n59203;
  assign n37194 = x155 & x204;
  assign n37195 = n37193 & n37194;
  assign n37196 = n37193 | n37194;
  assign n37197 = ~n37195 & n37196;
  assign n59204 = n36746 & n37197;
  assign n71992 = (n37197 & n58968) | (n37197 & n59204) | (n58968 & n59204);
  assign n71993 = (n37197 & n58967) | (n37197 & n59204) | (n58967 & n59204);
  assign n71994 = (n71647 & n71992) | (n71647 & n71993) | (n71992 & n71993);
  assign n59206 = n36746 | n37197;
  assign n71995 = n58968 | n59206;
  assign n71996 = n58967 | n59206;
  assign n71997 = (n71647 & n71995) | (n71647 & n71996) | (n71995 & n71996);
  assign n37200 = ~n71994 & n71997;
  assign n37201 = x154 & x205;
  assign n37202 = n37200 & n37201;
  assign n37203 = n37200 | n37201;
  assign n37204 = ~n37202 & n37203;
  assign n37205 = n71885 & n37204;
  assign n37206 = n71885 | n37204;
  assign n37207 = ~n37205 & n37206;
  assign n37208 = x153 & x206;
  assign n37209 = n37207 & n37208;
  assign n37210 = n37207 | n37208;
  assign n37211 = ~n37209 & n37210;
  assign n59085 = n36760 | n36762;
  assign n59208 = n37211 & n59085;
  assign n59209 = n36760 & n37211;
  assign n59210 = (n58851 & n59208) | (n58851 & n59209) | (n59208 & n59209);
  assign n59211 = n37211 | n59085;
  assign n59212 = n36760 | n37211;
  assign n59213 = (n58851 & n59211) | (n58851 & n59212) | (n59211 & n59212);
  assign n37214 = ~n59210 & n59213;
  assign n37215 = x152 & x207;
  assign n37216 = n37214 & n37215;
  assign n37217 = n37214 | n37215;
  assign n37218 = ~n37216 & n37217;
  assign n59214 = n36767 & n37218;
  assign n59215 = (n37218 & n71863) | (n37218 & n59214) | (n71863 & n59214);
  assign n59216 = n36767 | n37218;
  assign n59217 = n71863 | n59216;
  assign n37221 = ~n59215 & n59217;
  assign n37222 = x151 & x208;
  assign n37223 = n37221 & n37222;
  assign n37224 = n37221 | n37222;
  assign n37225 = ~n37223 & n37224;
  assign n59218 = n36774 & n37225;
  assign n59219 = (n37225 & n58982) | (n37225 & n59218) | (n58982 & n59218);
  assign n59220 = n36774 | n37225;
  assign n59221 = n58982 | n59220;
  assign n37228 = ~n59219 & n59221;
  assign n37229 = x150 & x209;
  assign n37230 = n37228 & n37229;
  assign n37231 = n37228 | n37229;
  assign n37232 = ~n37230 & n37231;
  assign n59222 = n36781 & n37232;
  assign n59223 = (n37232 & n58986) | (n37232 & n59222) | (n58986 & n59222);
  assign n59224 = n36781 | n37232;
  assign n59225 = n58986 | n59224;
  assign n37235 = ~n59223 & n59225;
  assign n37236 = x149 & x210;
  assign n37237 = n37235 & n37236;
  assign n37238 = n37235 | n37236;
  assign n37239 = ~n37237 & n37238;
  assign n59226 = n36788 & n37239;
  assign n59227 = (n37239 & n58990) | (n37239 & n59226) | (n58990 & n59226);
  assign n59228 = n36788 | n37239;
  assign n59229 = n58990 | n59228;
  assign n37242 = ~n59227 & n59229;
  assign n37243 = x148 & x211;
  assign n37244 = n37242 & n37243;
  assign n37245 = n37242 | n37243;
  assign n37246 = ~n37244 & n37245;
  assign n59230 = n36795 & n37246;
  assign n59231 = (n37246 & n58994) | (n37246 & n59230) | (n58994 & n59230);
  assign n59232 = n36795 | n37246;
  assign n59233 = n58994 | n59232;
  assign n37249 = ~n59231 & n59233;
  assign n37250 = x147 & x212;
  assign n37251 = n37249 & n37250;
  assign n37252 = n37249 | n37250;
  assign n37253 = ~n37251 & n37252;
  assign n59234 = n36802 & n37253;
  assign n59235 = (n37253 & n58998) | (n37253 & n59234) | (n58998 & n59234);
  assign n59236 = n36802 | n37253;
  assign n59237 = n58998 | n59236;
  assign n37256 = ~n59235 & n59237;
  assign n37257 = x146 & x213;
  assign n37258 = n37256 & n37257;
  assign n37259 = n37256 | n37257;
  assign n37260 = ~n37258 & n37259;
  assign n59238 = n36809 & n37260;
  assign n59239 = (n37260 & n59002) | (n37260 & n59238) | (n59002 & n59238);
  assign n59240 = n36809 | n37260;
  assign n59241 = n59002 | n59240;
  assign n37263 = ~n59239 & n59241;
  assign n37264 = x145 & x214;
  assign n37265 = n37263 & n37264;
  assign n37266 = n37263 | n37264;
  assign n37267 = ~n37265 & n37266;
  assign n59242 = n36816 & n37267;
  assign n59243 = (n37267 & n59006) | (n37267 & n59242) | (n59006 & n59242);
  assign n59244 = n36816 | n37267;
  assign n59245 = n59006 | n59244;
  assign n37270 = ~n59243 & n59245;
  assign n37271 = x144 & x215;
  assign n37272 = n37270 & n37271;
  assign n37273 = n37270 | n37271;
  assign n37274 = ~n37272 & n37273;
  assign n59246 = n36823 & n37274;
  assign n59247 = (n37274 & n59010) | (n37274 & n59246) | (n59010 & n59246);
  assign n59248 = n36823 | n37274;
  assign n59249 = n59010 | n59248;
  assign n37277 = ~n59247 & n59249;
  assign n37278 = x143 & x216;
  assign n37279 = n37277 & n37278;
  assign n37280 = n37277 | n37278;
  assign n37281 = ~n37279 & n37280;
  assign n59250 = n36830 & n37281;
  assign n59251 = (n37281 & n59014) | (n37281 & n59250) | (n59014 & n59250);
  assign n59252 = n36830 | n37281;
  assign n59253 = n59014 | n59252;
  assign n37284 = ~n59251 & n59253;
  assign n37285 = x142 & x217;
  assign n37286 = n37284 & n37285;
  assign n37287 = n37284 | n37285;
  assign n37288 = ~n37286 & n37287;
  assign n59254 = n36837 & n37288;
  assign n59255 = (n37288 & n59018) | (n37288 & n59254) | (n59018 & n59254);
  assign n59256 = n36837 | n37288;
  assign n59257 = n59018 | n59256;
  assign n37291 = ~n59255 & n59257;
  assign n37292 = x141 & x218;
  assign n37293 = n37291 & n37292;
  assign n37294 = n37291 | n37292;
  assign n37295 = ~n37293 & n37294;
  assign n59258 = n36844 & n37295;
  assign n59259 = (n37295 & n59022) | (n37295 & n59258) | (n59022 & n59258);
  assign n59260 = n36844 | n37295;
  assign n59261 = n59022 | n59260;
  assign n37298 = ~n59259 & n59261;
  assign n37299 = x140 & x219;
  assign n37300 = n37298 & n37299;
  assign n37301 = n37298 | n37299;
  assign n37302 = ~n37300 & n37301;
  assign n59262 = n36851 & n37302;
  assign n59263 = (n37302 & n59026) | (n37302 & n59262) | (n59026 & n59262);
  assign n59264 = n36851 | n37302;
  assign n59265 = n59026 | n59264;
  assign n37305 = ~n59263 & n59265;
  assign n37306 = x139 & x220;
  assign n37307 = n37305 & n37306;
  assign n37308 = n37305 | n37306;
  assign n37309 = ~n37307 & n37308;
  assign n59266 = n36858 & n37309;
  assign n59267 = (n37309 & n59030) | (n37309 & n59266) | (n59030 & n59266);
  assign n59268 = n36858 | n37309;
  assign n59269 = n59030 | n59268;
  assign n37312 = ~n59267 & n59269;
  assign n37313 = x138 & x221;
  assign n37314 = n37312 & n37313;
  assign n37315 = n37312 | n37313;
  assign n37316 = ~n37314 & n37315;
  assign n59270 = n36865 & n37316;
  assign n59271 = (n37316 & n59034) | (n37316 & n59270) | (n59034 & n59270);
  assign n59272 = n36865 | n37316;
  assign n59273 = n59034 | n59272;
  assign n37319 = ~n59271 & n59273;
  assign n37320 = x137 & x222;
  assign n37321 = n37319 & n37320;
  assign n37322 = n37319 | n37320;
  assign n37323 = ~n37321 & n37322;
  assign n59274 = n36872 & n37323;
  assign n59275 = (n37323 & n59038) | (n37323 & n59274) | (n59038 & n59274);
  assign n59276 = n36872 | n37323;
  assign n59277 = n59038 | n59276;
  assign n37326 = ~n59275 & n59277;
  assign n37327 = x136 & x223;
  assign n37328 = n37326 & n37327;
  assign n37329 = n37326 | n37327;
  assign n37330 = ~n37328 & n37329;
  assign n59278 = n36879 & n37330;
  assign n59279 = (n37330 & n59042) | (n37330 & n59278) | (n59042 & n59278);
  assign n59280 = n36879 | n37330;
  assign n59281 = n59042 | n59280;
  assign n37333 = ~n59279 & n59281;
  assign n37334 = x135 & x224;
  assign n37335 = n37333 & n37334;
  assign n37336 = n37333 | n37334;
  assign n37337 = ~n37335 & n37336;
  assign n59282 = n36886 & n37337;
  assign n59283 = (n37337 & n59046) | (n37337 & n59282) | (n59046 & n59282);
  assign n59284 = n36886 | n37337;
  assign n59285 = n59046 | n59284;
  assign n37340 = ~n59283 & n59285;
  assign n37341 = x134 & x225;
  assign n37342 = n37340 & n37341;
  assign n37343 = n37340 | n37341;
  assign n37344 = ~n37342 & n37343;
  assign n59286 = n36893 & n37344;
  assign n59287 = (n37344 & n59050) | (n37344 & n59286) | (n59050 & n59286);
  assign n59288 = n36893 | n37344;
  assign n59289 = n59050 | n59288;
  assign n37347 = ~n59287 & n59289;
  assign n37348 = x133 & x226;
  assign n37349 = n37347 & n37348;
  assign n37350 = n37347 | n37348;
  assign n37351 = ~n37349 & n37350;
  assign n59290 = n36900 & n37351;
  assign n59291 = (n37351 & n59054) | (n37351 & n59290) | (n59054 & n59290);
  assign n59292 = n36900 | n37351;
  assign n59293 = n59054 | n59292;
  assign n37354 = ~n59291 & n59293;
  assign n37355 = x132 & x227;
  assign n37356 = n37354 & n37355;
  assign n37357 = n37354 | n37355;
  assign n37358 = ~n37356 & n37357;
  assign n59294 = n36907 & n37358;
  assign n59295 = (n37358 & n59058) | (n37358 & n59294) | (n59058 & n59294);
  assign n59296 = n36907 | n37358;
  assign n59297 = n59058 | n59296;
  assign n37361 = ~n59295 & n59297;
  assign n37362 = x131 & x228;
  assign n37363 = n37361 & n37362;
  assign n37364 = n37361 | n37362;
  assign n37365 = ~n37363 & n37364;
  assign n59298 = n36914 & n37365;
  assign n59299 = (n37365 & n59062) | (n37365 & n59298) | (n59062 & n59298);
  assign n59300 = n36914 | n37365;
  assign n59301 = n59062 | n59300;
  assign n37368 = ~n59299 & n59301;
  assign n37369 = x130 & x229;
  assign n37370 = n37368 & n37369;
  assign n37371 = n37368 | n37369;
  assign n37372 = ~n37370 & n37371;
  assign n59302 = n36921 & n37372;
  assign n59303 = (n37372 & n59067) | (n37372 & n59302) | (n59067 & n59302);
  assign n59304 = n36921 | n37372;
  assign n59305 = n59067 | n59304;
  assign n37375 = ~n59303 & n59305;
  assign n37376 = x129 & x230;
  assign n37377 = n37375 & n37376;
  assign n37378 = n37375 | n37376;
  assign n37379 = ~n37377 & n37378;
  assign n59083 = n36928 | n36930;
  assign n59306 = n37379 & n59083;
  assign n59307 = n36928 & n37379;
  assign n59308 = (n58846 & n59306) | (n58846 & n59307) | (n59306 & n59307);
  assign n59309 = n37379 | n59083;
  assign n59310 = n36928 | n37379;
  assign n59311 = (n58846 & n59309) | (n58846 & n59310) | (n59309 & n59310);
  assign n37382 = ~n59308 & n59311;
  assign n37383 = x128 & x231;
  assign n37384 = n37382 & n37383;
  assign n37385 = n37382 | n37383;
  assign n37386 = ~n37384 & n37385;
  assign n59081 = n36935 | n36937;
  assign n71998 = n37386 & n59081;
  assign n71999 = n36935 & n37386;
  assign n72000 = (n58844 & n71998) | (n58844 & n71999) | (n71998 & n71999);
  assign n72001 = n37386 | n59081;
  assign n72002 = n36935 | n37386;
  assign n72003 = (n58844 & n72001) | (n58844 & n72002) | (n72001 & n72002);
  assign n37389 = ~n72000 & n72003;
  assign n37390 = x127 & x232;
  assign n37391 = n37389 & n37390;
  assign n37392 = n37389 | n37390;
  assign n37393 = ~n37391 & n37392;
  assign n59079 = n36942 | n36944;
  assign n72004 = n37393 & n59079;
  assign n72005 = n36942 & n37393;
  assign n72006 = (n58842 & n72004) | (n58842 & n72005) | (n72004 & n72005);
  assign n72007 = n37393 | n59079;
  assign n72008 = n36942 | n37393;
  assign n72009 = (n58842 & n72007) | (n58842 & n72008) | (n72007 & n72008);
  assign n37396 = ~n72006 & n72009;
  assign n37397 = x126 & x233;
  assign n37398 = n37396 & n37397;
  assign n37399 = n37396 | n37397;
  assign n37400 = ~n37398 & n37399;
  assign n37401 = n59078 & n37400;
  assign n37402 = n59078 | n37400;
  assign n37403 = ~n37401 & n37402;
  assign n37404 = x125 & x234;
  assign n37405 = n37403 & n37404;
  assign n37406 = n37403 | n37404;
  assign n37407 = ~n37405 & n37406;
  assign n37408 = n59076 & n37407;
  assign n37409 = n59076 | n37407;
  assign n37410 = ~n37408 & n37409;
  assign n37411 = x124 & x235;
  assign n37412 = n37410 & n37411;
  assign n37413 = n37410 | n37411;
  assign n37414 = ~n37412 & n37413;
  assign n37415 = n37001 & n37414;
  assign n37416 = n37001 | n37414;
  assign n37417 = ~n37415 & n37416;
  assign n37418 = x123 & x236;
  assign n37419 = n37417 & n37418;
  assign n37420 = n37417 | n37418;
  assign n37421 = ~n37419 & n37420;
  assign n37422 = n37000 & n37421;
  assign n37423 = n37000 | n37421;
  assign n37424 = ~n37422 & n37423;
  assign n37425 = x122 & x237;
  assign n37426 = n37424 & n37425;
  assign n37427 = n37424 | n37425;
  assign n37428 = ~n37426 & n37427;
  assign n37429 = n71880 & n37428;
  assign n37430 = n71880 | n37428;
  assign n37431 = ~n37429 & n37430;
  assign n37432 = x121 & x238;
  assign n37433 = n37431 & n37432;
  assign n37434 = n37431 | n37432;
  assign n37435 = ~n37433 & n37434;
  assign n37436 = n59074 & n37435;
  assign n37437 = n59074 | n37435;
  assign n37438 = ~n37436 & n37437;
  assign n37439 = x120 & x239;
  assign n37440 = n37438 & n37439;
  assign n37441 = n37438 | n37439;
  assign n37442 = ~n37440 & n37441;
  assign n37443 = n59072 & n37442;
  assign n37444 = n59072 | n37442;
  assign n37445 = ~n37443 & n37444;
  assign n59312 = n37440 | n59072;
  assign n59313 = (n37440 & n37442) | (n37440 & n59312) | (n37442 & n59312);
  assign n59314 = n37433 | n59074;
  assign n59315 = (n37433 & n37435) | (n37433 & n59314) | (n37435 & n59314);
  assign n72010 = n37426 | n71880;
  assign n72011 = (n37426 & n37428) | (n37426 & n72010) | (n37428 & n72010);
  assign n37449 = n37419 | n37422;
  assign n59316 = n37412 | n37414;
  assign n59317 = (n37001 & n37412) | (n37001 & n59316) | (n37412 & n59316);
  assign n59318 = n37405 | n37407;
  assign n59319 = (n37405 & n59076) | (n37405 & n59318) | (n59076 & n59318);
  assign n59080 = (n36942 & n58842) | (n36942 & n59079) | (n58842 & n59079);
  assign n59082 = (n36935 & n58844) | (n36935 & n59081) | (n58844 & n59081);
  assign n59332 = n37195 | n37197;
  assign n72014 = n36746 | n37195;
  assign n72015 = (n37195 & n37197) | (n37195 & n72014) | (n37197 & n72014);
  assign n72016 = (n58968 & n59332) | (n58968 & n72015) | (n59332 & n72015);
  assign n72017 = (n58967 & n59332) | (n58967 & n72015) | (n59332 & n72015);
  assign n72018 = (n71647 & n72016) | (n71647 & n72017) | (n72016 & n72017);
  assign n59337 = n37174 | n37176;
  assign n72019 = n36725 | n37174;
  assign n72020 = (n37174 & n37176) | (n37174 & n72019) | (n37176 & n72019);
  assign n72021 = (n58958 & n59337) | (n58958 & n72020) | (n59337 & n72020);
  assign n72022 = (n58957 & n59337) | (n58957 & n72020) | (n59337 & n72020);
  assign n72023 = (n71652 & n72021) | (n71652 & n72022) | (n72021 & n72022);
  assign n59099 = (n58717 & n71892) | (n58717 & n59098) | (n71892 & n59098);
  assign n59342 = n37153 | n37155;
  assign n72024 = n36704 | n37153;
  assign n72025 = (n37153 & n37155) | (n37153 & n72024) | (n37155 & n72024);
  assign n72026 = (n58948 & n59342) | (n58948 & n72025) | (n59342 & n72025);
  assign n72027 = (n58947 & n59342) | (n58947 & n72025) | (n59342 & n72025);
  assign n72028 = (n58619 & n72026) | (n58619 & n72027) | (n72026 & n72027);
  assign n59104 = (n58707 & n71894) | (n58707 & n59103) | (n71894 & n59103);
  assign n59347 = n37132 | n37134;
  assign n72029 = n36683 | n37132;
  assign n72030 = (n37132 & n37134) | (n37132 & n72029) | (n37134 & n72029);
  assign n72031 = (n58938 & n59347) | (n58938 & n72030) | (n59347 & n72030);
  assign n72032 = (n58937 & n59347) | (n58937 & n72030) | (n59347 & n72030);
  assign n72033 = (n58624 & n72031) | (n58624 & n72032) | (n72031 & n72032);
  assign n59109 = (n58697 & n71896) | (n58697 & n59108) | (n71896 & n59108);
  assign n59352 = n37111 | n37113;
  assign n72034 = n36662 | n37111;
  assign n72035 = (n37111 & n37113) | (n37111 & n72034) | (n37113 & n72034);
  assign n72036 = (n58928 & n59352) | (n58928 & n72035) | (n59352 & n72035);
  assign n72037 = (n58927 & n59352) | (n58927 & n72035) | (n59352 & n72035);
  assign n72038 = (n58629 & n72036) | (n58629 & n72037) | (n72036 & n72037);
  assign n58879 = (n58399 & n71799) | (n58399 & n71801) | (n71799 & n71801);
  assign n72041 = n36627 | n37076;
  assign n72042 = (n37076 & n37078) | (n37076 & n72041) | (n37078 & n72041);
  assign n72043 = n37076 | n37078;
  assign n72044 = (n37076 & n59120) | (n37076 & n72043) | (n59120 & n72043);
  assign n72045 = (n58883 & n72042) | (n58883 & n72044) | (n72042 & n72044);
  assign n72046 = (n71803 & n72042) | (n71803 & n72044) | (n72042 & n72044);
  assign n72047 = (n71569 & n72045) | (n71569 & n72046) | (n72045 & n72046);
  assign n37502 = x175 & x185;
  assign n59370 = n71913 | n71923;
  assign n72054 = n37502 & n59370;
  assign n72052 = n37057 | n71913;
  assign n72053 = (n71913 & n71921) | (n71913 & n72052) | (n71921 & n72052);
  assign n72055 = n37502 & n72053;
  assign n72056 = (n71693 & n72054) | (n71693 & n72055) | (n72054 & n72055);
  assign n72057 = n37502 | n59370;
  assign n72058 = n37502 | n72053;
  assign n72059 = (n71693 & n72057) | (n71693 & n72058) | (n72057 & n72058);
  assign n37505 = ~n72056 & n72059;
  assign n72048 = n37062 | n37064;
  assign n72049 = (n37062 & n59125) | (n37062 & n72048) | (n59125 & n72048);
  assign n72060 = n37505 & n72049;
  assign n72050 = n36613 | n37062;
  assign n72051 = (n37062 & n37064) | (n37062 & n72050) | (n37064 & n72050);
  assign n72061 = n37505 & n72051;
  assign n72062 = (n71810 & n72060) | (n71810 & n72061) | (n72060 & n72061);
  assign n72063 = n37505 | n72049;
  assign n72064 = n37505 | n72051;
  assign n72065 = (n71810 & n72063) | (n71810 & n72064) | (n72063 & n72064);
  assign n37508 = ~n72062 & n72065;
  assign n37509 = x174 & x186;
  assign n37510 = n37508 & n37509;
  assign n37511 = n37508 | n37509;
  assign n37512 = ~n37510 & n37511;
  assign n59364 = n37069 | n37071;
  assign n59372 = n37512 & n59364;
  assign n59373 = n37069 & n37512;
  assign n72066 = (n59123 & n59372) | (n59123 & n59373) | (n59372 & n59373);
  assign n72067 = (n59372 & n59373) | (n59372 & n71907) | (n59373 & n71907);
  assign n72068 = (n71667 & n72066) | (n71667 & n72067) | (n72066 & n72067);
  assign n59375 = n37512 | n59364;
  assign n59376 = n37069 | n37512;
  assign n72069 = (n59123 & n59375) | (n59123 & n59376) | (n59375 & n59376);
  assign n72070 = (n59375 & n59376) | (n59375 & n71907) | (n59376 & n71907);
  assign n72071 = (n71667 & n72069) | (n71667 & n72070) | (n72069 & n72070);
  assign n37515 = ~n72068 & n72071;
  assign n37516 = x173 & x187;
  assign n37517 = n37515 & n37516;
  assign n37518 = n37515 | n37516;
  assign n37519 = ~n37517 & n37518;
  assign n37520 = n72047 & n37519;
  assign n37521 = n72047 | n37519;
  assign n37522 = ~n37520 & n37521;
  assign n37523 = x172 & x188;
  assign n37524 = n37522 & n37523;
  assign n37525 = n37522 | n37523;
  assign n37526 = ~n37524 & n37525;
  assign n59359 = n37083 | n37085;
  assign n59378 = n37526 & n59359;
  assign n59379 = n37083 & n37526;
  assign n59380 = (n71905 & n59378) | (n71905 & n59379) | (n59378 & n59379);
  assign n59381 = n37526 | n59359;
  assign n59382 = n37083 | n37526;
  assign n59383 = (n71905 & n59381) | (n71905 & n59382) | (n59381 & n59382);
  assign n37529 = ~n59380 & n59383;
  assign n37530 = x171 & x189;
  assign n37531 = n37529 & n37530;
  assign n37532 = n37529 | n37530;
  assign n37533 = ~n37531 & n37532;
  assign n59357 = n37090 | n59152;
  assign n72072 = n37533 & n59357;
  assign n72039 = n36641 | n37090;
  assign n72040 = (n37090 & n37092) | (n37090 & n72039) | (n37092 & n72039);
  assign n72073 = n37533 & n72040;
  assign n72074 = (n58879 & n72072) | (n58879 & n72073) | (n72072 & n72073);
  assign n72075 = n37533 | n59357;
  assign n72076 = n37533 | n72040;
  assign n72077 = (n58879 & n72075) | (n58879 & n72076) | (n72075 & n72076);
  assign n37536 = ~n72074 & n72077;
  assign n37537 = x170 & x190;
  assign n37538 = n37536 & n37537;
  assign n37539 = n37536 | n37537;
  assign n37540 = ~n37538 & n37539;
  assign n59354 = n37097 | n37099;
  assign n59384 = n37540 & n59354;
  assign n59385 = n37097 & n37540;
  assign n72078 = (n59113 & n59384) | (n59113 & n59385) | (n59384 & n59385);
  assign n72079 = (n59384 & n59385) | (n59384 & n71898) | (n59385 & n71898);
  assign n72080 = (n58687 & n72078) | (n58687 & n72079) | (n72078 & n72079);
  assign n59387 = n37540 | n59354;
  assign n59388 = n37097 | n37540;
  assign n72081 = (n59113 & n59387) | (n59113 & n59388) | (n59387 & n59388);
  assign n72082 = (n59387 & n59388) | (n59387 & n71898) | (n59388 & n71898);
  assign n72083 = (n58687 & n72081) | (n58687 & n72082) | (n72081 & n72082);
  assign n37543 = ~n72080 & n72083;
  assign n37544 = x169 & x191;
  assign n37545 = n37543 & n37544;
  assign n37546 = n37543 | n37544;
  assign n37547 = ~n37545 & n37546;
  assign n59390 = n37104 & n37547;
  assign n59391 = (n37547 & n59160) | (n37547 & n59390) | (n59160 & n59390);
  assign n59392 = n37104 | n37547;
  assign n59393 = n59160 | n59392;
  assign n37550 = ~n59391 & n59393;
  assign n37551 = x168 & x192;
  assign n37552 = n37550 & n37551;
  assign n37553 = n37550 | n37551;
  assign n37554 = ~n37552 & n37553;
  assign n37555 = n72038 & n37554;
  assign n37556 = n72038 | n37554;
  assign n37557 = ~n37555 & n37556;
  assign n37558 = x167 & x193;
  assign n37559 = n37557 & n37558;
  assign n37560 = n37557 | n37558;
  assign n37561 = ~n37559 & n37560;
  assign n59349 = n37118 | n37120;
  assign n59394 = n37561 & n59349;
  assign n59395 = n37118 & n37561;
  assign n59396 = (n59109 & n59394) | (n59109 & n59395) | (n59394 & n59395);
  assign n59397 = n37561 | n59349;
  assign n59398 = n37118 | n37561;
  assign n59399 = (n59109 & n59397) | (n59109 & n59398) | (n59397 & n59398);
  assign n37564 = ~n59396 & n59399;
  assign n37565 = x166 & x194;
  assign n37566 = n37564 & n37565;
  assign n37567 = n37564 | n37565;
  assign n37568 = ~n37566 & n37567;
  assign n59400 = n37125 & n37568;
  assign n59401 = (n37568 & n59170) | (n37568 & n59400) | (n59170 & n59400);
  assign n59402 = n37125 | n37568;
  assign n59403 = n59170 | n59402;
  assign n37571 = ~n59401 & n59403;
  assign n37572 = x165 & x195;
  assign n37573 = n37571 & n37572;
  assign n37574 = n37571 | n37572;
  assign n37575 = ~n37573 & n37574;
  assign n37576 = n72033 & n37575;
  assign n37577 = n72033 | n37575;
  assign n37578 = ~n37576 & n37577;
  assign n37579 = x164 & x196;
  assign n37580 = n37578 & n37579;
  assign n37581 = n37578 | n37579;
  assign n37582 = ~n37580 & n37581;
  assign n59344 = n37139 | n37141;
  assign n59404 = n37582 & n59344;
  assign n59405 = n37139 & n37582;
  assign n59406 = (n59104 & n59404) | (n59104 & n59405) | (n59404 & n59405);
  assign n59407 = n37582 | n59344;
  assign n59408 = n37139 | n37582;
  assign n59409 = (n59104 & n59407) | (n59104 & n59408) | (n59407 & n59408);
  assign n37585 = ~n59406 & n59409;
  assign n37586 = x163 & x197;
  assign n37587 = n37585 & n37586;
  assign n37588 = n37585 | n37586;
  assign n37589 = ~n37587 & n37588;
  assign n59410 = n37146 & n37589;
  assign n59411 = (n37589 & n59180) | (n37589 & n59410) | (n59180 & n59410);
  assign n59412 = n37146 | n37589;
  assign n59413 = n59180 | n59412;
  assign n37592 = ~n59411 & n59413;
  assign n37593 = x162 & x198;
  assign n37594 = n37592 & n37593;
  assign n37595 = n37592 | n37593;
  assign n37596 = ~n37594 & n37595;
  assign n37597 = n72028 & n37596;
  assign n37598 = n72028 | n37596;
  assign n37599 = ~n37597 & n37598;
  assign n37600 = x161 & x199;
  assign n37601 = n37599 & n37600;
  assign n37602 = n37599 | n37600;
  assign n37603 = ~n37601 & n37602;
  assign n59339 = n37160 | n37162;
  assign n59414 = n37603 & n59339;
  assign n59415 = n37160 & n37603;
  assign n59416 = (n59099 & n59414) | (n59099 & n59415) | (n59414 & n59415);
  assign n59417 = n37603 | n59339;
  assign n59418 = n37160 | n37603;
  assign n59419 = (n59099 & n59417) | (n59099 & n59418) | (n59417 & n59418);
  assign n37606 = ~n59416 & n59419;
  assign n37607 = x160 & x200;
  assign n37608 = n37606 & n37607;
  assign n37609 = n37606 | n37607;
  assign n37610 = ~n37608 & n37609;
  assign n59420 = n37167 & n37610;
  assign n59421 = (n37610 & n59190) | (n37610 & n59420) | (n59190 & n59420);
  assign n59422 = n37167 | n37610;
  assign n59423 = n59190 | n59422;
  assign n37613 = ~n59421 & n59423;
  assign n37614 = x159 & x201;
  assign n37615 = n37613 & n37614;
  assign n37616 = n37613 | n37614;
  assign n37617 = ~n37615 & n37616;
  assign n37618 = n72023 & n37617;
  assign n37619 = n72023 | n37617;
  assign n37620 = ~n37618 & n37619;
  assign n37621 = x158 & x202;
  assign n37622 = n37620 & n37621;
  assign n37623 = n37620 | n37621;
  assign n37624 = ~n37622 & n37623;
  assign n59334 = n37181 | n37183;
  assign n59424 = n37624 & n59334;
  assign n59425 = n37181 & n37624;
  assign n59426 = (n71890 & n59424) | (n71890 & n59425) | (n59424 & n59425);
  assign n59427 = n37624 | n59334;
  assign n59428 = n37181 | n37624;
  assign n59429 = (n71890 & n59427) | (n71890 & n59428) | (n59427 & n59428);
  assign n37627 = ~n59426 & n59429;
  assign n37628 = x157 & x203;
  assign n37629 = n37627 & n37628;
  assign n37630 = n37627 | n37628;
  assign n37631 = ~n37629 & n37630;
  assign n59430 = n37188 & n37631;
  assign n72084 = (n37631 & n59199) | (n37631 & n59430) | (n59199 & n59430);
  assign n72085 = (n37631 & n59198) | (n37631 & n59430) | (n59198 & n59430);
  assign n72086 = (n71777 & n72084) | (n71777 & n72085) | (n72084 & n72085);
  assign n59432 = n37188 | n37631;
  assign n72087 = n59199 | n59432;
  assign n72088 = n59198 | n59432;
  assign n72089 = (n71777 & n72087) | (n71777 & n72088) | (n72087 & n72088);
  assign n37634 = ~n72086 & n72089;
  assign n37635 = x156 & x204;
  assign n37636 = n37634 & n37635;
  assign n37637 = n37634 | n37635;
  assign n37638 = ~n37636 & n37637;
  assign n37639 = n72018 & n37638;
  assign n37640 = n72018 | n37638;
  assign n37641 = ~n37639 & n37640;
  assign n37642 = x155 & x205;
  assign n37643 = n37641 & n37642;
  assign n37644 = n37641 | n37642;
  assign n37645 = ~n37643 & n37644;
  assign n59329 = n37202 | n37204;
  assign n59434 = n37645 & n59329;
  assign n59435 = n37202 & n37645;
  assign n59436 = (n71885 & n59434) | (n71885 & n59435) | (n59434 & n59435);
  assign n59437 = n37645 | n59329;
  assign n59438 = n37202 | n37645;
  assign n59439 = (n71885 & n59437) | (n71885 & n59438) | (n59437 & n59438);
  assign n37648 = ~n59436 & n59439;
  assign n37649 = x154 & x206;
  assign n37650 = n37648 & n37649;
  assign n37651 = n37648 | n37649;
  assign n37652 = ~n37650 & n37651;
  assign n59440 = n37209 & n37652;
  assign n72090 = (n37652 & n59209) | (n37652 & n59440) | (n59209 & n59440);
  assign n72091 = (n37652 & n59208) | (n37652 & n59440) | (n59208 & n59440);
  assign n72092 = (n58851 & n72090) | (n58851 & n72091) | (n72090 & n72091);
  assign n59442 = n37209 | n37652;
  assign n72093 = n59209 | n59442;
  assign n72094 = n59208 | n59442;
  assign n72095 = (n58851 & n72093) | (n58851 & n72094) | (n72093 & n72094);
  assign n37655 = ~n72092 & n72095;
  assign n37656 = x153 & x207;
  assign n37657 = n37655 & n37656;
  assign n37658 = n37655 | n37656;
  assign n37659 = ~n37657 & n37658;
  assign n59327 = n37216 | n37218;
  assign n72096 = n37659 & n59327;
  assign n72012 = n36767 | n37216;
  assign n72013 = (n37216 & n37218) | (n37216 & n72012) | (n37218 & n72012);
  assign n72097 = n37659 & n72013;
  assign n72098 = (n71863 & n72096) | (n71863 & n72097) | (n72096 & n72097);
  assign n72099 = n37659 | n59327;
  assign n72100 = n37659 | n72013;
  assign n72101 = (n71863 & n72099) | (n71863 & n72100) | (n72099 & n72100);
  assign n37662 = ~n72098 & n72101;
  assign n37663 = x152 & x208;
  assign n37664 = n37662 & n37663;
  assign n37665 = n37662 | n37663;
  assign n37666 = ~n37664 & n37665;
  assign n59444 = n37223 & n37666;
  assign n72102 = (n37666 & n59218) | (n37666 & n59444) | (n59218 & n59444);
  assign n72103 = (n37225 & n37666) | (n37225 & n59444) | (n37666 & n59444);
  assign n72104 = (n58982 & n72102) | (n58982 & n72103) | (n72102 & n72103);
  assign n59446 = n37223 | n37666;
  assign n72105 = n59218 | n59446;
  assign n72106 = n37225 | n59446;
  assign n72107 = (n58982 & n72105) | (n58982 & n72106) | (n72105 & n72106);
  assign n37669 = ~n72104 & n72107;
  assign n37670 = x151 & x209;
  assign n37671 = n37669 & n37670;
  assign n37672 = n37669 | n37670;
  assign n37673 = ~n37671 & n37672;
  assign n59448 = n37230 & n37673;
  assign n59449 = (n37673 & n59223) | (n37673 & n59448) | (n59223 & n59448);
  assign n59450 = n37230 | n37673;
  assign n59451 = n59223 | n59450;
  assign n37676 = ~n59449 & n59451;
  assign n37677 = x150 & x210;
  assign n37678 = n37676 & n37677;
  assign n37679 = n37676 | n37677;
  assign n37680 = ~n37678 & n37679;
  assign n59452 = n37237 & n37680;
  assign n59453 = (n37680 & n59227) | (n37680 & n59452) | (n59227 & n59452);
  assign n59454 = n37237 | n37680;
  assign n59455 = n59227 | n59454;
  assign n37683 = ~n59453 & n59455;
  assign n37684 = x149 & x211;
  assign n37685 = n37683 & n37684;
  assign n37686 = n37683 | n37684;
  assign n37687 = ~n37685 & n37686;
  assign n59456 = n37244 & n37687;
  assign n59457 = (n37687 & n59231) | (n37687 & n59456) | (n59231 & n59456);
  assign n59458 = n37244 | n37687;
  assign n59459 = n59231 | n59458;
  assign n37690 = ~n59457 & n59459;
  assign n37691 = x148 & x212;
  assign n37692 = n37690 & n37691;
  assign n37693 = n37690 | n37691;
  assign n37694 = ~n37692 & n37693;
  assign n59460 = n37251 & n37694;
  assign n59461 = (n37694 & n59235) | (n37694 & n59460) | (n59235 & n59460);
  assign n59462 = n37251 | n37694;
  assign n59463 = n59235 | n59462;
  assign n37697 = ~n59461 & n59463;
  assign n37698 = x147 & x213;
  assign n37699 = n37697 & n37698;
  assign n37700 = n37697 | n37698;
  assign n37701 = ~n37699 & n37700;
  assign n59464 = n37258 & n37701;
  assign n59465 = (n37701 & n59239) | (n37701 & n59464) | (n59239 & n59464);
  assign n59466 = n37258 | n37701;
  assign n59467 = n59239 | n59466;
  assign n37704 = ~n59465 & n59467;
  assign n37705 = x146 & x214;
  assign n37706 = n37704 & n37705;
  assign n37707 = n37704 | n37705;
  assign n37708 = ~n37706 & n37707;
  assign n59468 = n37265 & n37708;
  assign n59469 = (n37708 & n59243) | (n37708 & n59468) | (n59243 & n59468);
  assign n59470 = n37265 | n37708;
  assign n59471 = n59243 | n59470;
  assign n37711 = ~n59469 & n59471;
  assign n37712 = x145 & x215;
  assign n37713 = n37711 & n37712;
  assign n37714 = n37711 | n37712;
  assign n37715 = ~n37713 & n37714;
  assign n59472 = n37272 & n37715;
  assign n59473 = (n37715 & n59247) | (n37715 & n59472) | (n59247 & n59472);
  assign n59474 = n37272 | n37715;
  assign n59475 = n59247 | n59474;
  assign n37718 = ~n59473 & n59475;
  assign n37719 = x144 & x216;
  assign n37720 = n37718 & n37719;
  assign n37721 = n37718 | n37719;
  assign n37722 = ~n37720 & n37721;
  assign n59476 = n37279 & n37722;
  assign n59477 = (n37722 & n59251) | (n37722 & n59476) | (n59251 & n59476);
  assign n59478 = n37279 | n37722;
  assign n59479 = n59251 | n59478;
  assign n37725 = ~n59477 & n59479;
  assign n37726 = x143 & x217;
  assign n37727 = n37725 & n37726;
  assign n37728 = n37725 | n37726;
  assign n37729 = ~n37727 & n37728;
  assign n59480 = n37286 & n37729;
  assign n59481 = (n37729 & n59255) | (n37729 & n59480) | (n59255 & n59480);
  assign n59482 = n37286 | n37729;
  assign n59483 = n59255 | n59482;
  assign n37732 = ~n59481 & n59483;
  assign n37733 = x142 & x218;
  assign n37734 = n37732 & n37733;
  assign n37735 = n37732 | n37733;
  assign n37736 = ~n37734 & n37735;
  assign n59484 = n37293 & n37736;
  assign n59485 = (n37736 & n59259) | (n37736 & n59484) | (n59259 & n59484);
  assign n59486 = n37293 | n37736;
  assign n59487 = n59259 | n59486;
  assign n37739 = ~n59485 & n59487;
  assign n37740 = x141 & x219;
  assign n37741 = n37739 & n37740;
  assign n37742 = n37739 | n37740;
  assign n37743 = ~n37741 & n37742;
  assign n59488 = n37300 & n37743;
  assign n59489 = (n37743 & n59263) | (n37743 & n59488) | (n59263 & n59488);
  assign n59490 = n37300 | n37743;
  assign n59491 = n59263 | n59490;
  assign n37746 = ~n59489 & n59491;
  assign n37747 = x140 & x220;
  assign n37748 = n37746 & n37747;
  assign n37749 = n37746 | n37747;
  assign n37750 = ~n37748 & n37749;
  assign n59492 = n37307 & n37750;
  assign n59493 = (n37750 & n59267) | (n37750 & n59492) | (n59267 & n59492);
  assign n59494 = n37307 | n37750;
  assign n59495 = n59267 | n59494;
  assign n37753 = ~n59493 & n59495;
  assign n37754 = x139 & x221;
  assign n37755 = n37753 & n37754;
  assign n37756 = n37753 | n37754;
  assign n37757 = ~n37755 & n37756;
  assign n59496 = n37314 & n37757;
  assign n59497 = (n37757 & n59271) | (n37757 & n59496) | (n59271 & n59496);
  assign n59498 = n37314 | n37757;
  assign n59499 = n59271 | n59498;
  assign n37760 = ~n59497 & n59499;
  assign n37761 = x138 & x222;
  assign n37762 = n37760 & n37761;
  assign n37763 = n37760 | n37761;
  assign n37764 = ~n37762 & n37763;
  assign n59500 = n37321 & n37764;
  assign n59501 = (n37764 & n59275) | (n37764 & n59500) | (n59275 & n59500);
  assign n59502 = n37321 | n37764;
  assign n59503 = n59275 | n59502;
  assign n37767 = ~n59501 & n59503;
  assign n37768 = x137 & x223;
  assign n37769 = n37767 & n37768;
  assign n37770 = n37767 | n37768;
  assign n37771 = ~n37769 & n37770;
  assign n59504 = n37328 & n37771;
  assign n59505 = (n37771 & n59279) | (n37771 & n59504) | (n59279 & n59504);
  assign n59506 = n37328 | n37771;
  assign n59507 = n59279 | n59506;
  assign n37774 = ~n59505 & n59507;
  assign n37775 = x136 & x224;
  assign n37776 = n37774 & n37775;
  assign n37777 = n37774 | n37775;
  assign n37778 = ~n37776 & n37777;
  assign n59508 = n37335 & n37778;
  assign n59509 = (n37778 & n59283) | (n37778 & n59508) | (n59283 & n59508);
  assign n59510 = n37335 | n37778;
  assign n59511 = n59283 | n59510;
  assign n37781 = ~n59509 & n59511;
  assign n37782 = x135 & x225;
  assign n37783 = n37781 & n37782;
  assign n37784 = n37781 | n37782;
  assign n37785 = ~n37783 & n37784;
  assign n59512 = n37342 & n37785;
  assign n59513 = (n37785 & n59287) | (n37785 & n59512) | (n59287 & n59512);
  assign n59514 = n37342 | n37785;
  assign n59515 = n59287 | n59514;
  assign n37788 = ~n59513 & n59515;
  assign n37789 = x134 & x226;
  assign n37790 = n37788 & n37789;
  assign n37791 = n37788 | n37789;
  assign n37792 = ~n37790 & n37791;
  assign n59516 = n37349 & n37792;
  assign n59517 = (n37792 & n59291) | (n37792 & n59516) | (n59291 & n59516);
  assign n59518 = n37349 | n37792;
  assign n59519 = n59291 | n59518;
  assign n37795 = ~n59517 & n59519;
  assign n37796 = x133 & x227;
  assign n37797 = n37795 & n37796;
  assign n37798 = n37795 | n37796;
  assign n37799 = ~n37797 & n37798;
  assign n59520 = n37356 & n37799;
  assign n59521 = (n37799 & n59295) | (n37799 & n59520) | (n59295 & n59520);
  assign n59522 = n37356 | n37799;
  assign n59523 = n59295 | n59522;
  assign n37802 = ~n59521 & n59523;
  assign n37803 = x132 & x228;
  assign n37804 = n37802 & n37803;
  assign n37805 = n37802 | n37803;
  assign n37806 = ~n37804 & n37805;
  assign n59524 = n37363 & n37806;
  assign n59525 = (n37806 & n59299) | (n37806 & n59524) | (n59299 & n59524);
  assign n59526 = n37363 | n37806;
  assign n59527 = n59299 | n59526;
  assign n37809 = ~n59525 & n59527;
  assign n37810 = x131 & x229;
  assign n37811 = n37809 & n37810;
  assign n37812 = n37809 | n37810;
  assign n37813 = ~n37811 & n37812;
  assign n59528 = n37370 & n37813;
  assign n59529 = (n37813 & n59303) | (n37813 & n59528) | (n59303 & n59528);
  assign n59530 = n37370 | n37813;
  assign n59531 = n59303 | n59530;
  assign n37816 = ~n59529 & n59531;
  assign n37817 = x130 & x230;
  assign n37818 = n37816 & n37817;
  assign n37819 = n37816 | n37817;
  assign n37820 = ~n37818 & n37819;
  assign n59532 = n37377 & n37820;
  assign n59533 = (n37820 & n59308) | (n37820 & n59532) | (n59308 & n59532);
  assign n59534 = n37377 | n37820;
  assign n59535 = n59308 | n59534;
  assign n37823 = ~n59533 & n59535;
  assign n37824 = x129 & x231;
  assign n37825 = n37823 & n37824;
  assign n37826 = n37823 | n37824;
  assign n37827 = ~n37825 & n37826;
  assign n59324 = n37384 | n37386;
  assign n59536 = n37827 & n59324;
  assign n59537 = n37384 & n37827;
  assign n59538 = (n59082 & n59536) | (n59082 & n59537) | (n59536 & n59537);
  assign n59539 = n37827 | n59324;
  assign n59540 = n37384 | n37827;
  assign n59541 = (n59082 & n59539) | (n59082 & n59540) | (n59539 & n59540);
  assign n37830 = ~n59538 & n59541;
  assign n37831 = x128 & x232;
  assign n37832 = n37830 & n37831;
  assign n37833 = n37830 | n37831;
  assign n37834 = ~n37832 & n37833;
  assign n59322 = n37391 | n37393;
  assign n72108 = n37834 & n59322;
  assign n72109 = n37391 & n37834;
  assign n72110 = (n59080 & n72108) | (n59080 & n72109) | (n72108 & n72109);
  assign n72111 = n37834 | n59322;
  assign n72112 = n37391 | n37834;
  assign n72113 = (n59080 & n72111) | (n59080 & n72112) | (n72111 & n72112);
  assign n37837 = ~n72110 & n72113;
  assign n37838 = x127 & x233;
  assign n37839 = n37837 & n37838;
  assign n37840 = n37837 | n37838;
  assign n37841 = ~n37839 & n37840;
  assign n59320 = n37398 | n37400;
  assign n72114 = n37841 & n59320;
  assign n72115 = n37398 & n37841;
  assign n72116 = (n59078 & n72114) | (n59078 & n72115) | (n72114 & n72115);
  assign n72117 = n37841 | n59320;
  assign n72118 = n37398 | n37841;
  assign n72119 = (n59078 & n72117) | (n59078 & n72118) | (n72117 & n72118);
  assign n37844 = ~n72116 & n72119;
  assign n37845 = x126 & x234;
  assign n37846 = n37844 & n37845;
  assign n37847 = n37844 | n37845;
  assign n37848 = ~n37846 & n37847;
  assign n37849 = n59319 & n37848;
  assign n37850 = n59319 | n37848;
  assign n37851 = ~n37849 & n37850;
  assign n37852 = x125 & x235;
  assign n37853 = n37851 & n37852;
  assign n37854 = n37851 | n37852;
  assign n37855 = ~n37853 & n37854;
  assign n37856 = n59317 & n37855;
  assign n37857 = n59317 | n37855;
  assign n37858 = ~n37856 & n37857;
  assign n37859 = x124 & x236;
  assign n37860 = n37858 & n37859;
  assign n37861 = n37858 | n37859;
  assign n37862 = ~n37860 & n37861;
  assign n37863 = n37449 & n37862;
  assign n37864 = n37449 | n37862;
  assign n37865 = ~n37863 & n37864;
  assign n37866 = x123 & x237;
  assign n37867 = n37865 & n37866;
  assign n37868 = n37865 | n37866;
  assign n37869 = ~n37867 & n37868;
  assign n37870 = n72011 & n37869;
  assign n37871 = n72011 | n37869;
  assign n37872 = ~n37870 & n37871;
  assign n37873 = x122 & x238;
  assign n37874 = n37872 & n37873;
  assign n37875 = n37872 | n37873;
  assign n37876 = ~n37874 & n37875;
  assign n37877 = n59315 & n37876;
  assign n37878 = n59315 | n37876;
  assign n37879 = ~n37877 & n37878;
  assign n37880 = x121 & x239;
  assign n37881 = n37879 & n37880;
  assign n37882 = n37879 | n37880;
  assign n37883 = ~n37881 & n37882;
  assign n37884 = n59313 & n37883;
  assign n37885 = n59313 | n37883;
  assign n37886 = ~n37884 & n37885;
  assign n59542 = n37881 | n59313;
  assign n59543 = (n37881 & n37883) | (n37881 & n59542) | (n37883 & n59542);
  assign n59544 = n37874 | n59315;
  assign n59545 = (n37874 & n37876) | (n37874 & n59544) | (n37876 & n59544);
  assign n72120 = n37867 | n72011;
  assign n72121 = (n37867 & n37869) | (n37867 & n72120) | (n37869 & n72120);
  assign n59546 = n37860 | n37862;
  assign n59547 = (n37449 & n37860) | (n37449 & n59546) | (n37860 & n59546);
  assign n59548 = n37853 | n37855;
  assign n59549 = (n37853 & n59317) | (n37853 & n59548) | (n59317 & n59548);
  assign n59321 = (n37398 & n59078) | (n37398 & n59320) | (n59078 & n59320);
  assign n59323 = (n37391 & n59080) | (n37391 & n59322) | (n59080 & n59322);
  assign n59328 = (n71863 & n72013) | (n71863 & n59327) | (n72013 & n59327);
  assign n59559 = n37650 | n37652;
  assign n72122 = n37209 | n37650;
  assign n72123 = (n37650 & n37652) | (n37650 & n72122) | (n37652 & n72122);
  assign n72124 = (n59209 & n59559) | (n59209 & n72123) | (n59559 & n72123);
  assign n72125 = (n59208 & n59559) | (n59208 & n72123) | (n59559 & n72123);
  assign n72126 = (n58851 & n72124) | (n58851 & n72125) | (n72124 & n72125);
  assign n59564 = n37629 | n37631;
  assign n72127 = n37188 | n37629;
  assign n72128 = (n37629 & n37631) | (n37629 & n72127) | (n37631 & n72127);
  assign n72129 = (n59199 & n59564) | (n59199 & n72128) | (n59564 & n72128);
  assign n72130 = (n59198 & n59564) | (n59198 & n72128) | (n59564 & n72128);
  assign n72131 = (n71777 & n72129) | (n71777 & n72130) | (n72129 & n72130);
  assign n59114 = (n58687 & n71898) | (n58687 & n59113) | (n71898 & n59113);
  assign n72144 = n37069 | n37510;
  assign n72145 = (n37510 & n37512) | (n37510 & n72144) | (n37512 & n72144);
  assign n72146 = n37510 | n37512;
  assign n72147 = (n37510 & n59364) | (n37510 & n72146) | (n59364 & n72146);
  assign n72148 = (n59123 & n72145) | (n59123 & n72147) | (n72145 & n72147);
  assign n72149 = (n71907 & n72145) | (n71907 & n72147) | (n72145 & n72147);
  assign n72150 = (n71667 & n72148) | (n71667 & n72149) | (n72148 & n72149);
  assign n37942 = x175 & x186;
  assign n72151 = n37942 & n72056;
  assign n72152 = (n37505 & n37942) | (n37505 & n72151) | (n37942 & n72151);
  assign n72153 = n37942 & n72055;
  assign n72154 = n37942 & n72054;
  assign n72155 = (n71693 & n72153) | (n71693 & n72154) | (n72153 & n72154);
  assign n72156 = (n72049 & n72152) | (n72049 & n72155) | (n72152 & n72155);
  assign n72157 = (n72051 & n72152) | (n72051 & n72155) | (n72152 & n72155);
  assign n72158 = (n71810 & n72156) | (n71810 & n72157) | (n72156 & n72157);
  assign n72159 = n37942 | n72056;
  assign n72160 = n37505 | n72159;
  assign n72161 = n37942 | n72055;
  assign n72162 = n37942 | n72054;
  assign n72163 = (n71693 & n72161) | (n71693 & n72162) | (n72161 & n72162);
  assign n72164 = (n72049 & n72160) | (n72049 & n72163) | (n72160 & n72163);
  assign n72165 = (n72051 & n72160) | (n72051 & n72163) | (n72160 & n72163);
  assign n72166 = (n71810 & n72164) | (n71810 & n72165) | (n72164 & n72165);
  assign n37945 = ~n72158 & n72166;
  assign n37946 = n72150 & n37945;
  assign n37947 = n72150 | n37945;
  assign n37948 = ~n37946 & n37947;
  assign n37949 = x174 & x187;
  assign n37950 = n37948 & n37949;
  assign n37951 = n37948 | n37949;
  assign n37952 = ~n37950 & n37951;
  assign n59594 = n37517 | n37519;
  assign n59607 = n37952 & n59594;
  assign n59608 = n37517 & n37952;
  assign n59609 = (n72047 & n59607) | (n72047 & n59608) | (n59607 & n59608);
  assign n59610 = n37952 | n59594;
  assign n59611 = n37517 | n37952;
  assign n59612 = (n72047 & n59610) | (n72047 & n59611) | (n59610 & n59611);
  assign n37955 = ~n59609 & n59612;
  assign n37956 = x173 & x188;
  assign n37957 = n37955 & n37956;
  assign n37958 = n37955 | n37956;
  assign n37959 = ~n37957 & n37958;
  assign n59592 = n37524 | n59378;
  assign n72167 = n37959 & n59592;
  assign n72142 = n37083 | n37524;
  assign n72143 = (n37524 & n37526) | (n37524 & n72142) | (n37526 & n72142);
  assign n72168 = n37959 & n72143;
  assign n72169 = (n71905 & n72167) | (n71905 & n72168) | (n72167 & n72168);
  assign n72170 = n37959 | n59592;
  assign n72171 = n37959 | n72143;
  assign n72172 = (n71905 & n72170) | (n71905 & n72171) | (n72170 & n72171);
  assign n37962 = ~n72169 & n72172;
  assign n37963 = x172 & x189;
  assign n37964 = n37962 & n37963;
  assign n37965 = n37962 | n37963;
  assign n37966 = ~n37964 & n37965;
  assign n59589 = n37531 | n37533;
  assign n59613 = n37966 & n59589;
  assign n59614 = n37531 & n37966;
  assign n72173 = (n59357 & n59613) | (n59357 & n59614) | (n59613 & n59614);
  assign n72174 = (n59613 & n59614) | (n59613 & n72040) | (n59614 & n72040);
  assign n72175 = (n58879 & n72173) | (n58879 & n72174) | (n72173 & n72174);
  assign n59616 = n37966 | n59589;
  assign n59617 = n37531 | n37966;
  assign n72176 = (n59357 & n59616) | (n59357 & n59617) | (n59616 & n59617);
  assign n72177 = (n59616 & n59617) | (n59616 & n72040) | (n59617 & n72040);
  assign n72178 = (n58879 & n72176) | (n58879 & n72177) | (n72176 & n72177);
  assign n37969 = ~n72175 & n72178;
  assign n37970 = x171 & x190;
  assign n37971 = n37969 & n37970;
  assign n37972 = n37969 | n37970;
  assign n37973 = ~n37971 & n37972;
  assign n59587 = n37538 | n59384;
  assign n72179 = n37973 & n59587;
  assign n72140 = n37097 | n37538;
  assign n72141 = (n37538 & n37540) | (n37538 & n72140) | (n37540 & n72140);
  assign n72180 = n37973 & n72141;
  assign n72181 = (n59114 & n72179) | (n59114 & n72180) | (n72179 & n72180);
  assign n72182 = n37973 | n59587;
  assign n72183 = n37973 | n72141;
  assign n72184 = (n59114 & n72182) | (n59114 & n72183) | (n72182 & n72183);
  assign n37976 = ~n72181 & n72184;
  assign n37977 = x170 & x191;
  assign n37978 = n37976 & n37977;
  assign n37979 = n37976 | n37977;
  assign n37980 = ~n37978 & n37979;
  assign n59584 = n37545 | n37547;
  assign n72185 = n37980 & n59584;
  assign n72138 = n37104 | n37545;
  assign n72139 = (n37545 & n37547) | (n37545 & n72138) | (n37547 & n72138);
  assign n72186 = n37980 & n72139;
  assign n72187 = (n59160 & n72185) | (n59160 & n72186) | (n72185 & n72186);
  assign n72188 = n37980 | n59584;
  assign n72189 = n37980 | n72139;
  assign n72190 = (n59160 & n72188) | (n59160 & n72189) | (n72188 & n72189);
  assign n37983 = ~n72187 & n72190;
  assign n37984 = x169 & x192;
  assign n37985 = n37983 & n37984;
  assign n37986 = n37983 | n37984;
  assign n37987 = ~n37985 & n37986;
  assign n59581 = n37552 | n37554;
  assign n59619 = n37987 & n59581;
  assign n59620 = n37552 & n37987;
  assign n59621 = (n72038 & n59619) | (n72038 & n59620) | (n59619 & n59620);
  assign n59622 = n37987 | n59581;
  assign n59623 = n37552 | n37987;
  assign n59624 = (n72038 & n59622) | (n72038 & n59623) | (n59622 & n59623);
  assign n37990 = ~n59621 & n59624;
  assign n37991 = x168 & x193;
  assign n37992 = n37990 & n37991;
  assign n37993 = n37990 | n37991;
  assign n37994 = ~n37992 & n37993;
  assign n59625 = n37559 & n37994;
  assign n72191 = (n37994 & n59395) | (n37994 & n59625) | (n59395 & n59625);
  assign n72192 = (n37994 & n59394) | (n37994 & n59625) | (n59394 & n59625);
  assign n72193 = (n59109 & n72191) | (n59109 & n72192) | (n72191 & n72192);
  assign n59627 = n37559 | n37994;
  assign n72194 = n59395 | n59627;
  assign n72195 = n59394 | n59627;
  assign n72196 = (n59109 & n72194) | (n59109 & n72195) | (n72194 & n72195);
  assign n37997 = ~n72193 & n72196;
  assign n37998 = x167 & x194;
  assign n37999 = n37997 & n37998;
  assign n38000 = n37997 | n37998;
  assign n38001 = ~n37999 & n38000;
  assign n59579 = n37566 | n37568;
  assign n72197 = n38001 & n59579;
  assign n72136 = n37125 | n37566;
  assign n72137 = (n37566 & n37568) | (n37566 & n72136) | (n37568 & n72136);
  assign n72198 = n38001 & n72137;
  assign n72199 = (n59170 & n72197) | (n59170 & n72198) | (n72197 & n72198);
  assign n72200 = n38001 | n59579;
  assign n72201 = n38001 | n72137;
  assign n72202 = (n59170 & n72200) | (n59170 & n72201) | (n72200 & n72201);
  assign n38004 = ~n72199 & n72202;
  assign n38005 = x166 & x195;
  assign n38006 = n38004 & n38005;
  assign n38007 = n38004 | n38005;
  assign n38008 = ~n38006 & n38007;
  assign n59576 = n37573 | n37575;
  assign n59629 = n38008 & n59576;
  assign n59630 = n37573 & n38008;
  assign n59631 = (n72033 & n59629) | (n72033 & n59630) | (n59629 & n59630);
  assign n59632 = n38008 | n59576;
  assign n59633 = n37573 | n38008;
  assign n59634 = (n72033 & n59632) | (n72033 & n59633) | (n59632 & n59633);
  assign n38011 = ~n59631 & n59634;
  assign n38012 = x165 & x196;
  assign n38013 = n38011 & n38012;
  assign n38014 = n38011 | n38012;
  assign n38015 = ~n38013 & n38014;
  assign n59635 = n37580 & n38015;
  assign n72203 = (n38015 & n59405) | (n38015 & n59635) | (n59405 & n59635);
  assign n72204 = (n38015 & n59404) | (n38015 & n59635) | (n59404 & n59635);
  assign n72205 = (n59104 & n72203) | (n59104 & n72204) | (n72203 & n72204);
  assign n59637 = n37580 | n38015;
  assign n72206 = n59405 | n59637;
  assign n72207 = n59404 | n59637;
  assign n72208 = (n59104 & n72206) | (n59104 & n72207) | (n72206 & n72207);
  assign n38018 = ~n72205 & n72208;
  assign n38019 = x164 & x197;
  assign n38020 = n38018 & n38019;
  assign n38021 = n38018 | n38019;
  assign n38022 = ~n38020 & n38021;
  assign n59574 = n37587 | n37589;
  assign n72209 = n38022 & n59574;
  assign n72134 = n37146 | n37587;
  assign n72135 = (n37587 & n37589) | (n37587 & n72134) | (n37589 & n72134);
  assign n72210 = n38022 & n72135;
  assign n72211 = (n59180 & n72209) | (n59180 & n72210) | (n72209 & n72210);
  assign n72212 = n38022 | n59574;
  assign n72213 = n38022 | n72135;
  assign n72214 = (n59180 & n72212) | (n59180 & n72213) | (n72212 & n72213);
  assign n38025 = ~n72211 & n72214;
  assign n38026 = x163 & x198;
  assign n38027 = n38025 & n38026;
  assign n38028 = n38025 | n38026;
  assign n38029 = ~n38027 & n38028;
  assign n59571 = n37594 | n37596;
  assign n59639 = n38029 & n59571;
  assign n59640 = n37594 & n38029;
  assign n59641 = (n72028 & n59639) | (n72028 & n59640) | (n59639 & n59640);
  assign n59642 = n38029 | n59571;
  assign n59643 = n37594 | n38029;
  assign n59644 = (n72028 & n59642) | (n72028 & n59643) | (n59642 & n59643);
  assign n38032 = ~n59641 & n59644;
  assign n38033 = x162 & x199;
  assign n38034 = n38032 & n38033;
  assign n38035 = n38032 | n38033;
  assign n38036 = ~n38034 & n38035;
  assign n59645 = n37601 & n38036;
  assign n72215 = (n38036 & n59415) | (n38036 & n59645) | (n59415 & n59645);
  assign n72216 = (n38036 & n59414) | (n38036 & n59645) | (n59414 & n59645);
  assign n72217 = (n59099 & n72215) | (n59099 & n72216) | (n72215 & n72216);
  assign n59647 = n37601 | n38036;
  assign n72218 = n59415 | n59647;
  assign n72219 = n59414 | n59647;
  assign n72220 = (n59099 & n72218) | (n59099 & n72219) | (n72218 & n72219);
  assign n38039 = ~n72217 & n72220;
  assign n38040 = x161 & x200;
  assign n38041 = n38039 & n38040;
  assign n38042 = n38039 | n38040;
  assign n38043 = ~n38041 & n38042;
  assign n59569 = n37608 | n37610;
  assign n72221 = n38043 & n59569;
  assign n72132 = n37167 | n37608;
  assign n72133 = (n37608 & n37610) | (n37608 & n72132) | (n37610 & n72132);
  assign n72222 = n38043 & n72133;
  assign n72223 = (n59190 & n72221) | (n59190 & n72222) | (n72221 & n72222);
  assign n72224 = n38043 | n59569;
  assign n72225 = n38043 | n72133;
  assign n72226 = (n59190 & n72224) | (n59190 & n72225) | (n72224 & n72225);
  assign n38046 = ~n72223 & n72226;
  assign n38047 = x160 & x201;
  assign n38048 = n38046 & n38047;
  assign n38049 = n38046 | n38047;
  assign n38050 = ~n38048 & n38049;
  assign n59566 = n37615 | n37617;
  assign n59649 = n38050 & n59566;
  assign n59650 = n37615 & n38050;
  assign n59651 = (n72023 & n59649) | (n72023 & n59650) | (n59649 & n59650);
  assign n59652 = n38050 | n59566;
  assign n59653 = n37615 | n38050;
  assign n59654 = (n72023 & n59652) | (n72023 & n59653) | (n59652 & n59653);
  assign n38053 = ~n59651 & n59654;
  assign n38054 = x159 & x202;
  assign n38055 = n38053 & n38054;
  assign n38056 = n38053 | n38054;
  assign n38057 = ~n38055 & n38056;
  assign n59655 = n37622 & n38057;
  assign n72227 = (n38057 & n59425) | (n38057 & n59655) | (n59425 & n59655);
  assign n72228 = (n38057 & n59424) | (n38057 & n59655) | (n59424 & n59655);
  assign n72229 = (n71890 & n72227) | (n71890 & n72228) | (n72227 & n72228);
  assign n59657 = n37622 | n38057;
  assign n72230 = n59425 | n59657;
  assign n72231 = n59424 | n59657;
  assign n72232 = (n71890 & n72230) | (n71890 & n72231) | (n72230 & n72231);
  assign n38060 = ~n72229 & n72232;
  assign n38061 = x158 & x203;
  assign n38062 = n38060 & n38061;
  assign n38063 = n38060 | n38061;
  assign n38064 = ~n38062 & n38063;
  assign n38065 = n72131 & n38064;
  assign n38066 = n72131 | n38064;
  assign n38067 = ~n38065 & n38066;
  assign n38068 = x157 & x204;
  assign n38069 = n38067 & n38068;
  assign n38070 = n38067 | n38068;
  assign n38071 = ~n38069 & n38070;
  assign n59561 = n37636 | n37638;
  assign n59659 = n38071 & n59561;
  assign n59660 = n37636 & n38071;
  assign n59661 = (n72018 & n59659) | (n72018 & n59660) | (n59659 & n59660);
  assign n59662 = n38071 | n59561;
  assign n59663 = n37636 | n38071;
  assign n59664 = (n72018 & n59662) | (n72018 & n59663) | (n59662 & n59663);
  assign n38074 = ~n59661 & n59664;
  assign n38075 = x156 & x205;
  assign n38076 = n38074 & n38075;
  assign n38077 = n38074 | n38075;
  assign n38078 = ~n38076 & n38077;
  assign n59665 = n37643 & n38078;
  assign n72233 = (n38078 & n59435) | (n38078 & n59665) | (n59435 & n59665);
  assign n72234 = (n38078 & n59434) | (n38078 & n59665) | (n59434 & n59665);
  assign n72235 = (n71885 & n72233) | (n71885 & n72234) | (n72233 & n72234);
  assign n59667 = n37643 | n38078;
  assign n72236 = n59435 | n59667;
  assign n72237 = n59434 | n59667;
  assign n72238 = (n71885 & n72236) | (n71885 & n72237) | (n72236 & n72237);
  assign n38081 = ~n72235 & n72238;
  assign n38082 = x155 & x206;
  assign n38083 = n38081 & n38082;
  assign n38084 = n38081 | n38082;
  assign n38085 = ~n38083 & n38084;
  assign n38086 = n72126 & n38085;
  assign n38087 = n72126 | n38085;
  assign n38088 = ~n38086 & n38087;
  assign n38089 = x154 & x207;
  assign n38090 = n38088 & n38089;
  assign n38091 = n38088 | n38089;
  assign n38092 = ~n38090 & n38091;
  assign n59556 = n37657 | n37659;
  assign n59669 = n38092 & n59556;
  assign n59670 = n37657 & n38092;
  assign n59671 = (n59328 & n59669) | (n59328 & n59670) | (n59669 & n59670);
  assign n59672 = n38092 | n59556;
  assign n59673 = n37657 | n38092;
  assign n59674 = (n59328 & n59672) | (n59328 & n59673) | (n59672 & n59673);
  assign n38095 = ~n59671 & n59674;
  assign n38096 = x153 & x208;
  assign n38097 = n38095 & n38096;
  assign n38098 = n38095 | n38096;
  assign n38099 = ~n38097 & n38098;
  assign n59675 = n37664 & n38099;
  assign n59676 = (n38099 & n72104) | (n38099 & n59675) | (n72104 & n59675);
  assign n59677 = n37664 | n38099;
  assign n59678 = n72104 | n59677;
  assign n38102 = ~n59676 & n59678;
  assign n38103 = x152 & x209;
  assign n38104 = n38102 & n38103;
  assign n38105 = n38102 | n38103;
  assign n38106 = ~n38104 & n38105;
  assign n59679 = n37671 & n38106;
  assign n59680 = (n38106 & n59449) | (n38106 & n59679) | (n59449 & n59679);
  assign n59681 = n37671 | n38106;
  assign n59682 = n59449 | n59681;
  assign n38109 = ~n59680 & n59682;
  assign n38110 = x151 & x210;
  assign n38111 = n38109 & n38110;
  assign n38112 = n38109 | n38110;
  assign n38113 = ~n38111 & n38112;
  assign n59683 = n37678 & n38113;
  assign n59684 = (n38113 & n59453) | (n38113 & n59683) | (n59453 & n59683);
  assign n59685 = n37678 | n38113;
  assign n59686 = n59453 | n59685;
  assign n38116 = ~n59684 & n59686;
  assign n38117 = x150 & x211;
  assign n38118 = n38116 & n38117;
  assign n38119 = n38116 | n38117;
  assign n38120 = ~n38118 & n38119;
  assign n59687 = n37685 & n38120;
  assign n59688 = (n38120 & n59457) | (n38120 & n59687) | (n59457 & n59687);
  assign n59689 = n37685 | n38120;
  assign n59690 = n59457 | n59689;
  assign n38123 = ~n59688 & n59690;
  assign n38124 = x149 & x212;
  assign n38125 = n38123 & n38124;
  assign n38126 = n38123 | n38124;
  assign n38127 = ~n38125 & n38126;
  assign n59691 = n37692 & n38127;
  assign n59692 = (n38127 & n59461) | (n38127 & n59691) | (n59461 & n59691);
  assign n59693 = n37692 | n38127;
  assign n59694 = n59461 | n59693;
  assign n38130 = ~n59692 & n59694;
  assign n38131 = x148 & x213;
  assign n38132 = n38130 & n38131;
  assign n38133 = n38130 | n38131;
  assign n38134 = ~n38132 & n38133;
  assign n59695 = n37699 & n38134;
  assign n59696 = (n38134 & n59465) | (n38134 & n59695) | (n59465 & n59695);
  assign n59697 = n37699 | n38134;
  assign n59698 = n59465 | n59697;
  assign n38137 = ~n59696 & n59698;
  assign n38138 = x147 & x214;
  assign n38139 = n38137 & n38138;
  assign n38140 = n38137 | n38138;
  assign n38141 = ~n38139 & n38140;
  assign n59699 = n37706 & n38141;
  assign n59700 = (n38141 & n59469) | (n38141 & n59699) | (n59469 & n59699);
  assign n59701 = n37706 | n38141;
  assign n59702 = n59469 | n59701;
  assign n38144 = ~n59700 & n59702;
  assign n38145 = x146 & x215;
  assign n38146 = n38144 & n38145;
  assign n38147 = n38144 | n38145;
  assign n38148 = ~n38146 & n38147;
  assign n59703 = n37713 & n38148;
  assign n59704 = (n38148 & n59473) | (n38148 & n59703) | (n59473 & n59703);
  assign n59705 = n37713 | n38148;
  assign n59706 = n59473 | n59705;
  assign n38151 = ~n59704 & n59706;
  assign n38152 = x145 & x216;
  assign n38153 = n38151 & n38152;
  assign n38154 = n38151 | n38152;
  assign n38155 = ~n38153 & n38154;
  assign n59707 = n37720 & n38155;
  assign n59708 = (n38155 & n59477) | (n38155 & n59707) | (n59477 & n59707);
  assign n59709 = n37720 | n38155;
  assign n59710 = n59477 | n59709;
  assign n38158 = ~n59708 & n59710;
  assign n38159 = x144 & x217;
  assign n38160 = n38158 & n38159;
  assign n38161 = n38158 | n38159;
  assign n38162 = ~n38160 & n38161;
  assign n59711 = n37727 & n38162;
  assign n59712 = (n38162 & n59481) | (n38162 & n59711) | (n59481 & n59711);
  assign n59713 = n37727 | n38162;
  assign n59714 = n59481 | n59713;
  assign n38165 = ~n59712 & n59714;
  assign n38166 = x143 & x218;
  assign n38167 = n38165 & n38166;
  assign n38168 = n38165 | n38166;
  assign n38169 = ~n38167 & n38168;
  assign n59715 = n37734 & n38169;
  assign n59716 = (n38169 & n59485) | (n38169 & n59715) | (n59485 & n59715);
  assign n59717 = n37734 | n38169;
  assign n59718 = n59485 | n59717;
  assign n38172 = ~n59716 & n59718;
  assign n38173 = x142 & x219;
  assign n38174 = n38172 & n38173;
  assign n38175 = n38172 | n38173;
  assign n38176 = ~n38174 & n38175;
  assign n59719 = n37741 & n38176;
  assign n59720 = (n38176 & n59489) | (n38176 & n59719) | (n59489 & n59719);
  assign n59721 = n37741 | n38176;
  assign n59722 = n59489 | n59721;
  assign n38179 = ~n59720 & n59722;
  assign n38180 = x141 & x220;
  assign n38181 = n38179 & n38180;
  assign n38182 = n38179 | n38180;
  assign n38183 = ~n38181 & n38182;
  assign n59723 = n37748 & n38183;
  assign n59724 = (n38183 & n59493) | (n38183 & n59723) | (n59493 & n59723);
  assign n59725 = n37748 | n38183;
  assign n59726 = n59493 | n59725;
  assign n38186 = ~n59724 & n59726;
  assign n38187 = x140 & x221;
  assign n38188 = n38186 & n38187;
  assign n38189 = n38186 | n38187;
  assign n38190 = ~n38188 & n38189;
  assign n59727 = n37755 & n38190;
  assign n59728 = (n38190 & n59497) | (n38190 & n59727) | (n59497 & n59727);
  assign n59729 = n37755 | n38190;
  assign n59730 = n59497 | n59729;
  assign n38193 = ~n59728 & n59730;
  assign n38194 = x139 & x222;
  assign n38195 = n38193 & n38194;
  assign n38196 = n38193 | n38194;
  assign n38197 = ~n38195 & n38196;
  assign n59731 = n37762 & n38197;
  assign n59732 = (n38197 & n59501) | (n38197 & n59731) | (n59501 & n59731);
  assign n59733 = n37762 | n38197;
  assign n59734 = n59501 | n59733;
  assign n38200 = ~n59732 & n59734;
  assign n38201 = x138 & x223;
  assign n38202 = n38200 & n38201;
  assign n38203 = n38200 | n38201;
  assign n38204 = ~n38202 & n38203;
  assign n59735 = n37769 & n38204;
  assign n59736 = (n38204 & n59505) | (n38204 & n59735) | (n59505 & n59735);
  assign n59737 = n37769 | n38204;
  assign n59738 = n59505 | n59737;
  assign n38207 = ~n59736 & n59738;
  assign n38208 = x137 & x224;
  assign n38209 = n38207 & n38208;
  assign n38210 = n38207 | n38208;
  assign n38211 = ~n38209 & n38210;
  assign n59739 = n37776 & n38211;
  assign n59740 = (n38211 & n59509) | (n38211 & n59739) | (n59509 & n59739);
  assign n59741 = n37776 | n38211;
  assign n59742 = n59509 | n59741;
  assign n38214 = ~n59740 & n59742;
  assign n38215 = x136 & x225;
  assign n38216 = n38214 & n38215;
  assign n38217 = n38214 | n38215;
  assign n38218 = ~n38216 & n38217;
  assign n59743 = n37783 & n38218;
  assign n59744 = (n38218 & n59513) | (n38218 & n59743) | (n59513 & n59743);
  assign n59745 = n37783 | n38218;
  assign n59746 = n59513 | n59745;
  assign n38221 = ~n59744 & n59746;
  assign n38222 = x135 & x226;
  assign n38223 = n38221 & n38222;
  assign n38224 = n38221 | n38222;
  assign n38225 = ~n38223 & n38224;
  assign n59747 = n37790 & n38225;
  assign n59748 = (n38225 & n59517) | (n38225 & n59747) | (n59517 & n59747);
  assign n59749 = n37790 | n38225;
  assign n59750 = n59517 | n59749;
  assign n38228 = ~n59748 & n59750;
  assign n38229 = x134 & x227;
  assign n38230 = n38228 & n38229;
  assign n38231 = n38228 | n38229;
  assign n38232 = ~n38230 & n38231;
  assign n59751 = n37797 & n38232;
  assign n59752 = (n38232 & n59521) | (n38232 & n59751) | (n59521 & n59751);
  assign n59753 = n37797 | n38232;
  assign n59754 = n59521 | n59753;
  assign n38235 = ~n59752 & n59754;
  assign n38236 = x133 & x228;
  assign n38237 = n38235 & n38236;
  assign n38238 = n38235 | n38236;
  assign n38239 = ~n38237 & n38238;
  assign n59755 = n37804 & n38239;
  assign n59756 = (n38239 & n59525) | (n38239 & n59755) | (n59525 & n59755);
  assign n59757 = n37804 | n38239;
  assign n59758 = n59525 | n59757;
  assign n38242 = ~n59756 & n59758;
  assign n38243 = x132 & x229;
  assign n38244 = n38242 & n38243;
  assign n38245 = n38242 | n38243;
  assign n38246 = ~n38244 & n38245;
  assign n59759 = n37811 & n38246;
  assign n59760 = (n38246 & n59529) | (n38246 & n59759) | (n59529 & n59759);
  assign n59761 = n37811 | n38246;
  assign n59762 = n59529 | n59761;
  assign n38249 = ~n59760 & n59762;
  assign n38250 = x131 & x230;
  assign n38251 = n38249 & n38250;
  assign n38252 = n38249 | n38250;
  assign n38253 = ~n38251 & n38252;
  assign n59763 = n37818 & n38253;
  assign n59764 = (n38253 & n59533) | (n38253 & n59763) | (n59533 & n59763);
  assign n59765 = n37818 | n38253;
  assign n59766 = n59533 | n59765;
  assign n38256 = ~n59764 & n59766;
  assign n38257 = x130 & x231;
  assign n38258 = n38256 & n38257;
  assign n38259 = n38256 | n38257;
  assign n38260 = ~n38258 & n38259;
  assign n59767 = n37825 & n38260;
  assign n59768 = (n38260 & n59538) | (n38260 & n59767) | (n59538 & n59767);
  assign n59769 = n37825 | n38260;
  assign n59770 = n59538 | n59769;
  assign n38263 = ~n59768 & n59770;
  assign n38264 = x129 & x232;
  assign n38265 = n38263 & n38264;
  assign n38266 = n38263 | n38264;
  assign n38267 = ~n38265 & n38266;
  assign n59554 = n37832 | n37834;
  assign n59771 = n38267 & n59554;
  assign n59772 = n37832 & n38267;
  assign n59773 = (n59323 & n59771) | (n59323 & n59772) | (n59771 & n59772);
  assign n59774 = n38267 | n59554;
  assign n59775 = n37832 | n38267;
  assign n59776 = (n59323 & n59774) | (n59323 & n59775) | (n59774 & n59775);
  assign n38270 = ~n59773 & n59776;
  assign n38271 = x128 & x233;
  assign n38272 = n38270 & n38271;
  assign n38273 = n38270 | n38271;
  assign n38274 = ~n38272 & n38273;
  assign n59552 = n37839 | n37841;
  assign n72239 = n38274 & n59552;
  assign n72240 = n37839 & n38274;
  assign n72241 = (n59321 & n72239) | (n59321 & n72240) | (n72239 & n72240);
  assign n72242 = n38274 | n59552;
  assign n72243 = n37839 | n38274;
  assign n72244 = (n59321 & n72242) | (n59321 & n72243) | (n72242 & n72243);
  assign n38277 = ~n72241 & n72244;
  assign n38278 = x127 & x234;
  assign n38279 = n38277 & n38278;
  assign n38280 = n38277 | n38278;
  assign n38281 = ~n38279 & n38280;
  assign n59550 = n37846 | n37848;
  assign n72245 = n38281 & n59550;
  assign n72246 = n37846 & n38281;
  assign n72247 = (n59319 & n72245) | (n59319 & n72246) | (n72245 & n72246);
  assign n72248 = n38281 | n59550;
  assign n72249 = n37846 | n38281;
  assign n72250 = (n59319 & n72248) | (n59319 & n72249) | (n72248 & n72249);
  assign n38284 = ~n72247 & n72250;
  assign n38285 = x126 & x235;
  assign n38286 = n38284 & n38285;
  assign n38287 = n38284 | n38285;
  assign n38288 = ~n38286 & n38287;
  assign n38289 = n59549 & n38288;
  assign n38290 = n59549 | n38288;
  assign n38291 = ~n38289 & n38290;
  assign n38292 = x125 & x236;
  assign n38293 = n38291 & n38292;
  assign n38294 = n38291 | n38292;
  assign n38295 = ~n38293 & n38294;
  assign n38296 = n59547 & n38295;
  assign n38297 = n59547 | n38295;
  assign n38298 = ~n38296 & n38297;
  assign n38299 = x124 & x237;
  assign n38300 = n38298 & n38299;
  assign n38301 = n38298 | n38299;
  assign n38302 = ~n38300 & n38301;
  assign n38303 = n72121 & n38302;
  assign n38304 = n72121 | n38302;
  assign n38305 = ~n38303 & n38304;
  assign n38306 = x123 & x238;
  assign n38307 = n38305 & n38306;
  assign n38308 = n38305 | n38306;
  assign n38309 = ~n38307 & n38308;
  assign n38310 = n59545 & n38309;
  assign n38311 = n59545 | n38309;
  assign n38312 = ~n38310 & n38311;
  assign n38313 = x122 & x239;
  assign n38314 = n38312 & n38313;
  assign n38315 = n38312 | n38313;
  assign n38316 = ~n38314 & n38315;
  assign n38317 = n59543 & n38316;
  assign n38318 = n59543 | n38316;
  assign n38319 = ~n38317 & n38318;
  assign n59777 = n38314 | n59543;
  assign n59778 = (n38314 & n38316) | (n38314 & n59777) | (n38316 & n59777);
  assign n59779 = n38307 | n59545;
  assign n59780 = (n38307 & n38309) | (n38307 & n59779) | (n38309 & n59779);
  assign n59781 = n38300 | n38302;
  assign n59782 = (n72121 & n38300) | (n72121 & n59781) | (n38300 & n59781);
  assign n59783 = n38293 | n38295;
  assign n59784 = (n38293 & n59547) | (n38293 & n59783) | (n59547 & n59783);
  assign n59551 = (n37846 & n59319) | (n37846 & n59550) | (n59319 & n59550);
  assign n59553 = (n37839 & n59321) | (n37839 & n59552) | (n59321 & n59552);
  assign n59797 = n38076 | n38078;
  assign n72253 = n37643 | n38076;
  assign n72254 = (n38076 & n38078) | (n38076 & n72253) | (n38078 & n72253);
  assign n72255 = (n59435 & n59797) | (n59435 & n72254) | (n59797 & n72254);
  assign n72256 = (n59434 & n59797) | (n59434 & n72254) | (n59797 & n72254);
  assign n72257 = (n71885 & n72255) | (n71885 & n72256) | (n72255 & n72256);
  assign n59802 = n38055 | n38057;
  assign n72258 = n37622 | n38055;
  assign n72259 = (n38055 & n38057) | (n38055 & n72258) | (n38057 & n72258);
  assign n72260 = (n59425 & n59802) | (n59425 & n72259) | (n59802 & n72259);
  assign n72261 = (n59424 & n59802) | (n59424 & n72259) | (n59802 & n72259);
  assign n72262 = (n71890 & n72260) | (n71890 & n72261) | (n72260 & n72261);
  assign n59570 = (n59190 & n72133) | (n59190 & n59569) | (n72133 & n59569);
  assign n59807 = n38034 | n38036;
  assign n72263 = n37601 | n38034;
  assign n72264 = (n38034 & n38036) | (n38034 & n72263) | (n38036 & n72263);
  assign n72265 = (n59415 & n59807) | (n59415 & n72264) | (n59807 & n72264);
  assign n72266 = (n59414 & n59807) | (n59414 & n72264) | (n59807 & n72264);
  assign n72267 = (n59099 & n72265) | (n59099 & n72266) | (n72265 & n72266);
  assign n59575 = (n59180 & n72135) | (n59180 & n59574) | (n72135 & n59574);
  assign n59812 = n38013 | n38015;
  assign n72268 = n37580 | n38013;
  assign n72269 = (n38013 & n38015) | (n38013 & n72268) | (n38015 & n72268);
  assign n72270 = (n59405 & n59812) | (n59405 & n72269) | (n59812 & n72269);
  assign n72271 = (n59404 & n59812) | (n59404 & n72269) | (n59812 & n72269);
  assign n72272 = (n59104 & n72270) | (n59104 & n72271) | (n72270 & n72271);
  assign n59580 = (n59170 & n72137) | (n59170 & n59579) | (n72137 & n59579);
  assign n59817 = n37992 | n37994;
  assign n72273 = n37559 | n37992;
  assign n72274 = (n37992 & n37994) | (n37992 & n72273) | (n37994 & n72273);
  assign n72275 = (n59395 & n59817) | (n59395 & n72274) | (n59817 & n72274);
  assign n72276 = (n59394 & n59817) | (n59394 & n72274) | (n59817 & n72274);
  assign n72277 = (n59109 & n72275) | (n59109 & n72276) | (n72275 & n72276);
  assign n59585 = (n59160 & n72139) | (n59160 & n59584) | (n72139 & n59584);
  assign n72278 = n37531 | n37964;
  assign n72279 = (n37964 & n37966) | (n37964 & n72278) | (n37966 & n72278);
  assign n72280 = n37964 | n37966;
  assign n72281 = (n37964 & n59589) | (n37964 & n72280) | (n59589 & n72280);
  assign n72282 = (n59357 & n72279) | (n59357 & n72281) | (n72279 & n72281);
  assign n72283 = (n72040 & n72279) | (n72040 & n72281) | (n72279 & n72281);
  assign n72284 = (n58879 & n72282) | (n58879 & n72283) | (n72282 & n72283);
  assign n38374 = x175 & x187;
  assign n72287 = n38374 & n72158;
  assign n72288 = (n37945 & n38374) | (n37945 & n72287) | (n38374 & n72287);
  assign n59834 = n38374 & n72158;
  assign n59835 = (n72150 & n72288) | (n72150 & n59834) | (n72288 & n59834);
  assign n72289 = n38374 | n72158;
  assign n72290 = n37945 | n72289;
  assign n59837 = n38374 | n72158;
  assign n59838 = (n72150 & n72290) | (n72150 & n59837) | (n72290 & n59837);
  assign n38377 = ~n59835 & n59838;
  assign n59829 = n37950 | n59607;
  assign n72291 = n38377 & n59829;
  assign n72285 = n37517 | n37950;
  assign n72286 = (n37950 & n37952) | (n37950 & n72285) | (n37952 & n72285);
  assign n72292 = n38377 & n72286;
  assign n72293 = (n72047 & n72291) | (n72047 & n72292) | (n72291 & n72292);
  assign n72294 = n38377 | n59829;
  assign n72295 = n38377 | n72286;
  assign n72296 = (n72047 & n72294) | (n72047 & n72295) | (n72294 & n72295);
  assign n38380 = ~n72293 & n72296;
  assign n38381 = x174 & x188;
  assign n38382 = n38380 & n38381;
  assign n38383 = n38380 | n38381;
  assign n38384 = ~n38382 & n38383;
  assign n59826 = n37957 | n37959;
  assign n59839 = n38384 & n59826;
  assign n59840 = n37957 & n38384;
  assign n72297 = (n59592 & n59839) | (n59592 & n59840) | (n59839 & n59840);
  assign n72298 = (n59839 & n59840) | (n59839 & n72143) | (n59840 & n72143);
  assign n72299 = (n71905 & n72297) | (n71905 & n72298) | (n72297 & n72298);
  assign n59842 = n38384 | n59826;
  assign n59843 = n37957 | n38384;
  assign n72300 = (n59592 & n59842) | (n59592 & n59843) | (n59842 & n59843);
  assign n72301 = (n59842 & n59843) | (n59842 & n72143) | (n59843 & n72143);
  assign n72302 = (n71905 & n72300) | (n71905 & n72301) | (n72300 & n72301);
  assign n38387 = ~n72299 & n72302;
  assign n38388 = x173 & x189;
  assign n38389 = n38387 & n38388;
  assign n38390 = n38387 | n38388;
  assign n38391 = ~n38389 & n38390;
  assign n38392 = n72284 & n38391;
  assign n38393 = n72284 | n38391;
  assign n38394 = ~n38392 & n38393;
  assign n38395 = x172 & x190;
  assign n38396 = n38394 & n38395;
  assign n38397 = n38394 | n38395;
  assign n38398 = ~n38396 & n38397;
  assign n59821 = n37971 | n37973;
  assign n59845 = n38398 & n59821;
  assign n59846 = n37971 & n38398;
  assign n72303 = (n59587 & n59845) | (n59587 & n59846) | (n59845 & n59846);
  assign n72304 = (n59845 & n59846) | (n59845 & n72141) | (n59846 & n72141);
  assign n72305 = (n59114 & n72303) | (n59114 & n72304) | (n72303 & n72304);
  assign n59848 = n38398 | n59821;
  assign n59849 = n37971 | n38398;
  assign n72306 = (n59587 & n59848) | (n59587 & n59849) | (n59848 & n59849);
  assign n72307 = (n59848 & n59849) | (n59848 & n72141) | (n59849 & n72141);
  assign n72308 = (n59114 & n72306) | (n59114 & n72307) | (n72306 & n72307);
  assign n38401 = ~n72305 & n72308;
  assign n38402 = x171 & x191;
  assign n38403 = n38401 & n38402;
  assign n38404 = n38401 | n38402;
  assign n38405 = ~n38403 & n38404;
  assign n59819 = n37978 | n37980;
  assign n59851 = n38405 & n59819;
  assign n59852 = n37978 & n38405;
  assign n59853 = (n59585 & n59851) | (n59585 & n59852) | (n59851 & n59852);
  assign n59854 = n38405 | n59819;
  assign n59855 = n37978 | n38405;
  assign n59856 = (n59585 & n59854) | (n59585 & n59855) | (n59854 & n59855);
  assign n38408 = ~n59853 & n59856;
  assign n38409 = x170 & x192;
  assign n38410 = n38408 & n38409;
  assign n38411 = n38408 | n38409;
  assign n38412 = ~n38410 & n38411;
  assign n59857 = n37985 & n38412;
  assign n59858 = (n38412 & n59621) | (n38412 & n59857) | (n59621 & n59857);
  assign n59859 = n37985 | n38412;
  assign n59860 = n59621 | n59859;
  assign n38415 = ~n59858 & n59860;
  assign n38416 = x169 & x193;
  assign n38417 = n38415 & n38416;
  assign n38418 = n38415 | n38416;
  assign n38419 = ~n38417 & n38418;
  assign n38420 = n72277 & n38419;
  assign n38421 = n72277 | n38419;
  assign n38422 = ~n38420 & n38421;
  assign n38423 = x168 & x194;
  assign n38424 = n38422 & n38423;
  assign n38425 = n38422 | n38423;
  assign n38426 = ~n38424 & n38425;
  assign n59814 = n37999 | n38001;
  assign n59861 = n38426 & n59814;
  assign n59862 = n37999 & n38426;
  assign n59863 = (n59580 & n59861) | (n59580 & n59862) | (n59861 & n59862);
  assign n59864 = n38426 | n59814;
  assign n59865 = n37999 | n38426;
  assign n59866 = (n59580 & n59864) | (n59580 & n59865) | (n59864 & n59865);
  assign n38429 = ~n59863 & n59866;
  assign n38430 = x167 & x195;
  assign n38431 = n38429 & n38430;
  assign n38432 = n38429 | n38430;
  assign n38433 = ~n38431 & n38432;
  assign n59867 = n38006 & n38433;
  assign n59868 = (n38433 & n59631) | (n38433 & n59867) | (n59631 & n59867);
  assign n59869 = n38006 | n38433;
  assign n59870 = n59631 | n59869;
  assign n38436 = ~n59868 & n59870;
  assign n38437 = x166 & x196;
  assign n38438 = n38436 & n38437;
  assign n38439 = n38436 | n38437;
  assign n38440 = ~n38438 & n38439;
  assign n38441 = n72272 & n38440;
  assign n38442 = n72272 | n38440;
  assign n38443 = ~n38441 & n38442;
  assign n38444 = x165 & x197;
  assign n38445 = n38443 & n38444;
  assign n38446 = n38443 | n38444;
  assign n38447 = ~n38445 & n38446;
  assign n59809 = n38020 | n38022;
  assign n59871 = n38447 & n59809;
  assign n59872 = n38020 & n38447;
  assign n59873 = (n59575 & n59871) | (n59575 & n59872) | (n59871 & n59872);
  assign n59874 = n38447 | n59809;
  assign n59875 = n38020 | n38447;
  assign n59876 = (n59575 & n59874) | (n59575 & n59875) | (n59874 & n59875);
  assign n38450 = ~n59873 & n59876;
  assign n38451 = x164 & x198;
  assign n38452 = n38450 & n38451;
  assign n38453 = n38450 | n38451;
  assign n38454 = ~n38452 & n38453;
  assign n59877 = n38027 & n38454;
  assign n59878 = (n38454 & n59641) | (n38454 & n59877) | (n59641 & n59877);
  assign n59879 = n38027 | n38454;
  assign n59880 = n59641 | n59879;
  assign n38457 = ~n59878 & n59880;
  assign n38458 = x163 & x199;
  assign n38459 = n38457 & n38458;
  assign n38460 = n38457 | n38458;
  assign n38461 = ~n38459 & n38460;
  assign n38462 = n72267 & n38461;
  assign n38463 = n72267 | n38461;
  assign n38464 = ~n38462 & n38463;
  assign n38465 = x162 & x200;
  assign n38466 = n38464 & n38465;
  assign n38467 = n38464 | n38465;
  assign n38468 = ~n38466 & n38467;
  assign n59804 = n38041 | n38043;
  assign n59881 = n38468 & n59804;
  assign n59882 = n38041 & n38468;
  assign n59883 = (n59570 & n59881) | (n59570 & n59882) | (n59881 & n59882);
  assign n59884 = n38468 | n59804;
  assign n59885 = n38041 | n38468;
  assign n59886 = (n59570 & n59884) | (n59570 & n59885) | (n59884 & n59885);
  assign n38471 = ~n59883 & n59886;
  assign n38472 = x161 & x201;
  assign n38473 = n38471 & n38472;
  assign n38474 = n38471 | n38472;
  assign n38475 = ~n38473 & n38474;
  assign n59887 = n38048 & n38475;
  assign n59888 = (n38475 & n59651) | (n38475 & n59887) | (n59651 & n59887);
  assign n59889 = n38048 | n38475;
  assign n59890 = n59651 | n59889;
  assign n38478 = ~n59888 & n59890;
  assign n38479 = x160 & x202;
  assign n38480 = n38478 & n38479;
  assign n38481 = n38478 | n38479;
  assign n38482 = ~n38480 & n38481;
  assign n38483 = n72262 & n38482;
  assign n38484 = n72262 | n38482;
  assign n38485 = ~n38483 & n38484;
  assign n38486 = x159 & x203;
  assign n38487 = n38485 & n38486;
  assign n38488 = n38485 | n38486;
  assign n38489 = ~n38487 & n38488;
  assign n59799 = n38062 | n38064;
  assign n59891 = n38489 & n59799;
  assign n59892 = n38062 & n38489;
  assign n59893 = (n72131 & n59891) | (n72131 & n59892) | (n59891 & n59892);
  assign n59894 = n38489 | n59799;
  assign n59895 = n38062 | n38489;
  assign n59896 = (n72131 & n59894) | (n72131 & n59895) | (n59894 & n59895);
  assign n38492 = ~n59893 & n59896;
  assign n38493 = x158 & x204;
  assign n38494 = n38492 & n38493;
  assign n38495 = n38492 | n38493;
  assign n38496 = ~n38494 & n38495;
  assign n59897 = n38069 & n38496;
  assign n72309 = (n38496 & n59660) | (n38496 & n59897) | (n59660 & n59897);
  assign n72310 = (n38496 & n59659) | (n38496 & n59897) | (n59659 & n59897);
  assign n72311 = (n72018 & n72309) | (n72018 & n72310) | (n72309 & n72310);
  assign n59899 = n38069 | n38496;
  assign n72312 = n59660 | n59899;
  assign n72313 = n59659 | n59899;
  assign n72314 = (n72018 & n72312) | (n72018 & n72313) | (n72312 & n72313);
  assign n38499 = ~n72311 & n72314;
  assign n38500 = x157 & x205;
  assign n38501 = n38499 & n38500;
  assign n38502 = n38499 | n38500;
  assign n38503 = ~n38501 & n38502;
  assign n38504 = n72257 & n38503;
  assign n38505 = n72257 | n38503;
  assign n38506 = ~n38504 & n38505;
  assign n38507 = x156 & x206;
  assign n38508 = n38506 & n38507;
  assign n38509 = n38506 | n38507;
  assign n38510 = ~n38508 & n38509;
  assign n59794 = n38083 | n38085;
  assign n59901 = n38510 & n59794;
  assign n59902 = n38083 & n38510;
  assign n59903 = (n72126 & n59901) | (n72126 & n59902) | (n59901 & n59902);
  assign n59904 = n38510 | n59794;
  assign n59905 = n38083 | n38510;
  assign n59906 = (n72126 & n59904) | (n72126 & n59905) | (n59904 & n59905);
  assign n38513 = ~n59903 & n59906;
  assign n38514 = x155 & x207;
  assign n38515 = n38513 & n38514;
  assign n38516 = n38513 | n38514;
  assign n38517 = ~n38515 & n38516;
  assign n59907 = n38090 & n38517;
  assign n72315 = (n38517 & n59670) | (n38517 & n59907) | (n59670 & n59907);
  assign n72316 = (n38517 & n59669) | (n38517 & n59907) | (n59669 & n59907);
  assign n72317 = (n59328 & n72315) | (n59328 & n72316) | (n72315 & n72316);
  assign n59909 = n38090 | n38517;
  assign n72318 = n59670 | n59909;
  assign n72319 = n59669 | n59909;
  assign n72320 = (n59328 & n72318) | (n59328 & n72319) | (n72318 & n72319);
  assign n38520 = ~n72317 & n72320;
  assign n38521 = x154 & x208;
  assign n38522 = n38520 & n38521;
  assign n38523 = n38520 | n38521;
  assign n38524 = ~n38522 & n38523;
  assign n59792 = n38097 | n38099;
  assign n72321 = n38524 & n59792;
  assign n72251 = n37664 | n38097;
  assign n72252 = (n38097 & n38099) | (n38097 & n72251) | (n38099 & n72251);
  assign n72322 = n38524 & n72252;
  assign n72323 = (n72104 & n72321) | (n72104 & n72322) | (n72321 & n72322);
  assign n72324 = n38524 | n59792;
  assign n72325 = n38524 | n72252;
  assign n72326 = (n72104 & n72324) | (n72104 & n72325) | (n72324 & n72325);
  assign n38527 = ~n72323 & n72326;
  assign n38528 = x153 & x209;
  assign n38529 = n38527 & n38528;
  assign n38530 = n38527 | n38528;
  assign n38531 = ~n38529 & n38530;
  assign n59911 = n38104 & n38531;
  assign n72327 = (n38531 & n59679) | (n38531 & n59911) | (n59679 & n59911);
  assign n72328 = (n38106 & n38531) | (n38106 & n59911) | (n38531 & n59911);
  assign n72329 = (n59449 & n72327) | (n59449 & n72328) | (n72327 & n72328);
  assign n59913 = n38104 | n38531;
  assign n72330 = n59679 | n59913;
  assign n72331 = n38106 | n59913;
  assign n72332 = (n59449 & n72330) | (n59449 & n72331) | (n72330 & n72331);
  assign n38534 = ~n72329 & n72332;
  assign n38535 = x152 & x210;
  assign n38536 = n38534 & n38535;
  assign n38537 = n38534 | n38535;
  assign n38538 = ~n38536 & n38537;
  assign n59915 = n38111 & n38538;
  assign n59916 = (n38538 & n59684) | (n38538 & n59915) | (n59684 & n59915);
  assign n59917 = n38111 | n38538;
  assign n59918 = n59684 | n59917;
  assign n38541 = ~n59916 & n59918;
  assign n38542 = x151 & x211;
  assign n38543 = n38541 & n38542;
  assign n38544 = n38541 | n38542;
  assign n38545 = ~n38543 & n38544;
  assign n59919 = n38118 & n38545;
  assign n59920 = (n38545 & n59688) | (n38545 & n59919) | (n59688 & n59919);
  assign n59921 = n38118 | n38545;
  assign n59922 = n59688 | n59921;
  assign n38548 = ~n59920 & n59922;
  assign n38549 = x150 & x212;
  assign n38550 = n38548 & n38549;
  assign n38551 = n38548 | n38549;
  assign n38552 = ~n38550 & n38551;
  assign n59923 = n38125 & n38552;
  assign n59924 = (n38552 & n59692) | (n38552 & n59923) | (n59692 & n59923);
  assign n59925 = n38125 | n38552;
  assign n59926 = n59692 | n59925;
  assign n38555 = ~n59924 & n59926;
  assign n38556 = x149 & x213;
  assign n38557 = n38555 & n38556;
  assign n38558 = n38555 | n38556;
  assign n38559 = ~n38557 & n38558;
  assign n59927 = n38132 & n38559;
  assign n59928 = (n38559 & n59696) | (n38559 & n59927) | (n59696 & n59927);
  assign n59929 = n38132 | n38559;
  assign n59930 = n59696 | n59929;
  assign n38562 = ~n59928 & n59930;
  assign n38563 = x148 & x214;
  assign n38564 = n38562 & n38563;
  assign n38565 = n38562 | n38563;
  assign n38566 = ~n38564 & n38565;
  assign n59931 = n38139 & n38566;
  assign n59932 = (n38566 & n59700) | (n38566 & n59931) | (n59700 & n59931);
  assign n59933 = n38139 | n38566;
  assign n59934 = n59700 | n59933;
  assign n38569 = ~n59932 & n59934;
  assign n38570 = x147 & x215;
  assign n38571 = n38569 & n38570;
  assign n38572 = n38569 | n38570;
  assign n38573 = ~n38571 & n38572;
  assign n59935 = n38146 & n38573;
  assign n59936 = (n38573 & n59704) | (n38573 & n59935) | (n59704 & n59935);
  assign n59937 = n38146 | n38573;
  assign n59938 = n59704 | n59937;
  assign n38576 = ~n59936 & n59938;
  assign n38577 = x146 & x216;
  assign n38578 = n38576 & n38577;
  assign n38579 = n38576 | n38577;
  assign n38580 = ~n38578 & n38579;
  assign n59939 = n38153 & n38580;
  assign n59940 = (n38580 & n59708) | (n38580 & n59939) | (n59708 & n59939);
  assign n59941 = n38153 | n38580;
  assign n59942 = n59708 | n59941;
  assign n38583 = ~n59940 & n59942;
  assign n38584 = x145 & x217;
  assign n38585 = n38583 & n38584;
  assign n38586 = n38583 | n38584;
  assign n38587 = ~n38585 & n38586;
  assign n59943 = n38160 & n38587;
  assign n59944 = (n38587 & n59712) | (n38587 & n59943) | (n59712 & n59943);
  assign n59945 = n38160 | n38587;
  assign n59946 = n59712 | n59945;
  assign n38590 = ~n59944 & n59946;
  assign n38591 = x144 & x218;
  assign n38592 = n38590 & n38591;
  assign n38593 = n38590 | n38591;
  assign n38594 = ~n38592 & n38593;
  assign n59947 = n38167 & n38594;
  assign n59948 = (n38594 & n59716) | (n38594 & n59947) | (n59716 & n59947);
  assign n59949 = n38167 | n38594;
  assign n59950 = n59716 | n59949;
  assign n38597 = ~n59948 & n59950;
  assign n38598 = x143 & x219;
  assign n38599 = n38597 & n38598;
  assign n38600 = n38597 | n38598;
  assign n38601 = ~n38599 & n38600;
  assign n59951 = n38174 & n38601;
  assign n59952 = (n38601 & n59720) | (n38601 & n59951) | (n59720 & n59951);
  assign n59953 = n38174 | n38601;
  assign n59954 = n59720 | n59953;
  assign n38604 = ~n59952 & n59954;
  assign n38605 = x142 & x220;
  assign n38606 = n38604 & n38605;
  assign n38607 = n38604 | n38605;
  assign n38608 = ~n38606 & n38607;
  assign n59955 = n38181 & n38608;
  assign n59956 = (n38608 & n59724) | (n38608 & n59955) | (n59724 & n59955);
  assign n59957 = n38181 | n38608;
  assign n59958 = n59724 | n59957;
  assign n38611 = ~n59956 & n59958;
  assign n38612 = x141 & x221;
  assign n38613 = n38611 & n38612;
  assign n38614 = n38611 | n38612;
  assign n38615 = ~n38613 & n38614;
  assign n59959 = n38188 & n38615;
  assign n59960 = (n38615 & n59728) | (n38615 & n59959) | (n59728 & n59959);
  assign n59961 = n38188 | n38615;
  assign n59962 = n59728 | n59961;
  assign n38618 = ~n59960 & n59962;
  assign n38619 = x140 & x222;
  assign n38620 = n38618 & n38619;
  assign n38621 = n38618 | n38619;
  assign n38622 = ~n38620 & n38621;
  assign n59963 = n38195 & n38622;
  assign n59964 = (n38622 & n59732) | (n38622 & n59963) | (n59732 & n59963);
  assign n59965 = n38195 | n38622;
  assign n59966 = n59732 | n59965;
  assign n38625 = ~n59964 & n59966;
  assign n38626 = x139 & x223;
  assign n38627 = n38625 & n38626;
  assign n38628 = n38625 | n38626;
  assign n38629 = ~n38627 & n38628;
  assign n59967 = n38202 & n38629;
  assign n59968 = (n38629 & n59736) | (n38629 & n59967) | (n59736 & n59967);
  assign n59969 = n38202 | n38629;
  assign n59970 = n59736 | n59969;
  assign n38632 = ~n59968 & n59970;
  assign n38633 = x138 & x224;
  assign n38634 = n38632 & n38633;
  assign n38635 = n38632 | n38633;
  assign n38636 = ~n38634 & n38635;
  assign n59971 = n38209 & n38636;
  assign n59972 = (n38636 & n59740) | (n38636 & n59971) | (n59740 & n59971);
  assign n59973 = n38209 | n38636;
  assign n59974 = n59740 | n59973;
  assign n38639 = ~n59972 & n59974;
  assign n38640 = x137 & x225;
  assign n38641 = n38639 & n38640;
  assign n38642 = n38639 | n38640;
  assign n38643 = ~n38641 & n38642;
  assign n59975 = n38216 & n38643;
  assign n59976 = (n38643 & n59744) | (n38643 & n59975) | (n59744 & n59975);
  assign n59977 = n38216 | n38643;
  assign n59978 = n59744 | n59977;
  assign n38646 = ~n59976 & n59978;
  assign n38647 = x136 & x226;
  assign n38648 = n38646 & n38647;
  assign n38649 = n38646 | n38647;
  assign n38650 = ~n38648 & n38649;
  assign n59979 = n38223 & n38650;
  assign n59980 = (n38650 & n59748) | (n38650 & n59979) | (n59748 & n59979);
  assign n59981 = n38223 | n38650;
  assign n59982 = n59748 | n59981;
  assign n38653 = ~n59980 & n59982;
  assign n38654 = x135 & x227;
  assign n38655 = n38653 & n38654;
  assign n38656 = n38653 | n38654;
  assign n38657 = ~n38655 & n38656;
  assign n59983 = n38230 & n38657;
  assign n59984 = (n38657 & n59752) | (n38657 & n59983) | (n59752 & n59983);
  assign n59985 = n38230 | n38657;
  assign n59986 = n59752 | n59985;
  assign n38660 = ~n59984 & n59986;
  assign n38661 = x134 & x228;
  assign n38662 = n38660 & n38661;
  assign n38663 = n38660 | n38661;
  assign n38664 = ~n38662 & n38663;
  assign n59987 = n38237 & n38664;
  assign n59988 = (n38664 & n59756) | (n38664 & n59987) | (n59756 & n59987);
  assign n59989 = n38237 | n38664;
  assign n59990 = n59756 | n59989;
  assign n38667 = ~n59988 & n59990;
  assign n38668 = x133 & x229;
  assign n38669 = n38667 & n38668;
  assign n38670 = n38667 | n38668;
  assign n38671 = ~n38669 & n38670;
  assign n59991 = n38244 & n38671;
  assign n59992 = (n38671 & n59760) | (n38671 & n59991) | (n59760 & n59991);
  assign n59993 = n38244 | n38671;
  assign n59994 = n59760 | n59993;
  assign n38674 = ~n59992 & n59994;
  assign n38675 = x132 & x230;
  assign n38676 = n38674 & n38675;
  assign n38677 = n38674 | n38675;
  assign n38678 = ~n38676 & n38677;
  assign n59995 = n38251 & n38678;
  assign n59996 = (n38678 & n59764) | (n38678 & n59995) | (n59764 & n59995);
  assign n59997 = n38251 | n38678;
  assign n59998 = n59764 | n59997;
  assign n38681 = ~n59996 & n59998;
  assign n38682 = x131 & x231;
  assign n38683 = n38681 & n38682;
  assign n38684 = n38681 | n38682;
  assign n38685 = ~n38683 & n38684;
  assign n59999 = n38258 & n38685;
  assign n60000 = (n38685 & n59768) | (n38685 & n59999) | (n59768 & n59999);
  assign n60001 = n38258 | n38685;
  assign n60002 = n59768 | n60001;
  assign n38688 = ~n60000 & n60002;
  assign n38689 = x130 & x232;
  assign n38690 = n38688 & n38689;
  assign n38691 = n38688 | n38689;
  assign n38692 = ~n38690 & n38691;
  assign n60003 = n38265 & n38692;
  assign n60004 = (n38692 & n59773) | (n38692 & n60003) | (n59773 & n60003);
  assign n60005 = n38265 | n38692;
  assign n60006 = n59773 | n60005;
  assign n38695 = ~n60004 & n60006;
  assign n38696 = x129 & x233;
  assign n38697 = n38695 & n38696;
  assign n38698 = n38695 | n38696;
  assign n38699 = ~n38697 & n38698;
  assign n59789 = n38272 | n38274;
  assign n60007 = n38699 & n59789;
  assign n60008 = n38272 & n38699;
  assign n60009 = (n59553 & n60007) | (n59553 & n60008) | (n60007 & n60008);
  assign n60010 = n38699 | n59789;
  assign n60011 = n38272 | n38699;
  assign n60012 = (n59553 & n60010) | (n59553 & n60011) | (n60010 & n60011);
  assign n38702 = ~n60009 & n60012;
  assign n38703 = x128 & x234;
  assign n38704 = n38702 & n38703;
  assign n38705 = n38702 | n38703;
  assign n38706 = ~n38704 & n38705;
  assign n59787 = n38279 | n38281;
  assign n72333 = n38706 & n59787;
  assign n72334 = n38279 & n38706;
  assign n72335 = (n59551 & n72333) | (n59551 & n72334) | (n72333 & n72334);
  assign n72336 = n38706 | n59787;
  assign n72337 = n38279 | n38706;
  assign n72338 = (n59551 & n72336) | (n59551 & n72337) | (n72336 & n72337);
  assign n38709 = ~n72335 & n72338;
  assign n38710 = x127 & x235;
  assign n38711 = n38709 & n38710;
  assign n38712 = n38709 | n38710;
  assign n38713 = ~n38711 & n38712;
  assign n59785 = n38286 | n38288;
  assign n72339 = n38713 & n59785;
  assign n72340 = n38286 & n38713;
  assign n72341 = (n59549 & n72339) | (n59549 & n72340) | (n72339 & n72340);
  assign n72342 = n38713 | n59785;
  assign n72343 = n38286 | n38713;
  assign n72344 = (n59549 & n72342) | (n59549 & n72343) | (n72342 & n72343);
  assign n38716 = ~n72341 & n72344;
  assign n38717 = x126 & x236;
  assign n38718 = n38716 & n38717;
  assign n38719 = n38716 | n38717;
  assign n38720 = ~n38718 & n38719;
  assign n38721 = n59784 & n38720;
  assign n38722 = n59784 | n38720;
  assign n38723 = ~n38721 & n38722;
  assign n38724 = x125 & x237;
  assign n38725 = n38723 & n38724;
  assign n38726 = n38723 | n38724;
  assign n38727 = ~n38725 & n38726;
  assign n38728 = n59782 & n38727;
  assign n38729 = n59782 | n38727;
  assign n38730 = ~n38728 & n38729;
  assign n38731 = x124 & x238;
  assign n38732 = n38730 & n38731;
  assign n38733 = n38730 | n38731;
  assign n38734 = ~n38732 & n38733;
  assign n38735 = n59780 & n38734;
  assign n38736 = n59780 | n38734;
  assign n38737 = ~n38735 & n38736;
  assign n38738 = x123 & x239;
  assign n38739 = n38737 & n38738;
  assign n38740 = n38737 | n38738;
  assign n38741 = ~n38739 & n38740;
  assign n38742 = n59778 & n38741;
  assign n38743 = n59778 | n38741;
  assign n38744 = ~n38742 & n38743;
  assign n38745 = n38739 | n38742;
  assign n38746 = n38732 | n38735;
  assign n60013 = n38725 | n38727;
  assign n60014 = (n38725 & n59782) | (n38725 & n60013) | (n59782 & n60013);
  assign n59786 = (n38286 & n59549) | (n38286 & n59785) | (n59549 & n59785);
  assign n59788 = (n38279 & n59551) | (n38279 & n59787) | (n59551 & n59787);
  assign n59793 = (n72104 & n72252) | (n72104 & n59792) | (n72252 & n59792);
  assign n60024 = n38515 | n38517;
  assign n72345 = n38090 | n38515;
  assign n72346 = (n38515 & n38517) | (n38515 & n72345) | (n38517 & n72345);
  assign n72347 = (n59670 & n60024) | (n59670 & n72346) | (n60024 & n72346);
  assign n72348 = (n59669 & n60024) | (n59669 & n72346) | (n60024 & n72346);
  assign n72349 = (n59328 & n72347) | (n59328 & n72348) | (n72347 & n72348);
  assign n60029 = n38494 | n38496;
  assign n72350 = n38069 | n38494;
  assign n72351 = (n38494 & n38496) | (n38494 & n72350) | (n38496 & n72350);
  assign n72352 = (n59660 & n60029) | (n59660 & n72351) | (n60029 & n72351);
  assign n72353 = (n59659 & n60029) | (n59659 & n72351) | (n60029 & n72351);
  assign n72354 = (n72018 & n72352) | (n72018 & n72353) | (n72352 & n72353);
  assign n59588 = (n59114 & n72141) | (n59114 & n59587) | (n72141 & n59587);
  assign n72365 = n37957 | n38382;
  assign n72366 = (n38382 & n38384) | (n38382 & n72365) | (n38384 & n72365);
  assign n72367 = n38382 | n38384;
  assign n72368 = (n38382 & n59826) | (n38382 & n72367) | (n59826 & n72367);
  assign n72369 = (n59592 & n72366) | (n59592 & n72368) | (n72366 & n72368);
  assign n72370 = (n72143 & n72366) | (n72143 & n72368) | (n72366 & n72368);
  assign n72371 = (n71905 & n72369) | (n71905 & n72370) | (n72369 & n72370);
  assign n38798 = x175 & x188;
  assign n72373 = n38798 & n72288;
  assign n72374 = n38798 & n59834;
  assign n72375 = (n72150 & n72373) | (n72150 & n72374) | (n72373 & n72374);
  assign n72372 = (n38377 & n38798) | (n38377 & n72375) | (n38798 & n72375);
  assign n72376 = (n59829 & n72372) | (n59829 & n72375) | (n72372 & n72375);
  assign n72377 = (n72286 & n72372) | (n72286 & n72375) | (n72372 & n72375);
  assign n72378 = (n72047 & n72376) | (n72047 & n72377) | (n72376 & n72377);
  assign n72380 = n38798 | n72288;
  assign n72381 = n38798 | n59834;
  assign n72382 = (n72150 & n72380) | (n72150 & n72381) | (n72380 & n72381);
  assign n72379 = n38377 | n72382;
  assign n72383 = (n59829 & n72379) | (n59829 & n72382) | (n72379 & n72382);
  assign n72384 = (n72286 & n72379) | (n72286 & n72382) | (n72379 & n72382);
  assign n72385 = (n72047 & n72383) | (n72047 & n72384) | (n72383 & n72384);
  assign n38801 = ~n72378 & n72385;
  assign n38802 = n72371 & n38801;
  assign n38803 = n72371 | n38801;
  assign n38804 = ~n38802 & n38803;
  assign n38805 = x174 & x189;
  assign n38806 = n38804 & n38805;
  assign n38807 = n38804 | n38805;
  assign n38808 = ~n38806 & n38807;
  assign n60054 = n38389 | n38391;
  assign n60067 = n38808 & n60054;
  assign n60068 = n38389 & n38808;
  assign n60069 = (n72284 & n60067) | (n72284 & n60068) | (n60067 & n60068);
  assign n60070 = n38808 | n60054;
  assign n60071 = n38389 | n38808;
  assign n60072 = (n72284 & n60070) | (n72284 & n60071) | (n60070 & n60071);
  assign n38811 = ~n60069 & n60072;
  assign n38812 = x173 & x190;
  assign n38813 = n38811 & n38812;
  assign n38814 = n38811 | n38812;
  assign n38815 = ~n38813 & n38814;
  assign n60052 = n38396 | n59845;
  assign n72386 = n38815 & n60052;
  assign n72363 = n37971 | n38396;
  assign n72364 = (n38396 & n38398) | (n38396 & n72363) | (n38398 & n72363);
  assign n72387 = n38815 & n72364;
  assign n72388 = (n59588 & n72386) | (n59588 & n72387) | (n72386 & n72387);
  assign n72389 = n38815 | n60052;
  assign n72390 = n38815 | n72364;
  assign n72391 = (n59588 & n72389) | (n59588 & n72390) | (n72389 & n72390);
  assign n38818 = ~n72388 & n72391;
  assign n38819 = x172 & x191;
  assign n38820 = n38818 & n38819;
  assign n38821 = n38818 | n38819;
  assign n38822 = ~n38820 & n38821;
  assign n60073 = n38403 & n38822;
  assign n72392 = (n38822 & n59851) | (n38822 & n60073) | (n59851 & n60073);
  assign n72393 = (n38822 & n59852) | (n38822 & n60073) | (n59852 & n60073);
  assign n72394 = (n59585 & n72392) | (n59585 & n72393) | (n72392 & n72393);
  assign n60075 = n38403 | n38822;
  assign n72395 = n59851 | n60075;
  assign n72396 = n59852 | n60075;
  assign n72397 = (n59585 & n72395) | (n59585 & n72396) | (n72395 & n72396);
  assign n38825 = ~n72394 & n72397;
  assign n38826 = x171 & x192;
  assign n38827 = n38825 & n38826;
  assign n38828 = n38825 | n38826;
  assign n38829 = ~n38827 & n38828;
  assign n60049 = n38410 | n38412;
  assign n72398 = n38829 & n60049;
  assign n72361 = n37985 | n38410;
  assign n72362 = (n38410 & n38412) | (n38410 & n72361) | (n38412 & n72361);
  assign n72399 = n38829 & n72362;
  assign n72400 = (n59621 & n72398) | (n59621 & n72399) | (n72398 & n72399);
  assign n72401 = n38829 | n60049;
  assign n72402 = n38829 | n72362;
  assign n72403 = (n59621 & n72401) | (n59621 & n72402) | (n72401 & n72402);
  assign n38832 = ~n72400 & n72403;
  assign n38833 = x170 & x193;
  assign n38834 = n38832 & n38833;
  assign n38835 = n38832 | n38833;
  assign n38836 = ~n38834 & n38835;
  assign n60046 = n38417 | n38419;
  assign n60077 = n38836 & n60046;
  assign n60078 = n38417 & n38836;
  assign n60079 = (n72277 & n60077) | (n72277 & n60078) | (n60077 & n60078);
  assign n60080 = n38836 | n60046;
  assign n60081 = n38417 | n38836;
  assign n60082 = (n72277 & n60080) | (n72277 & n60081) | (n60080 & n60081);
  assign n38839 = ~n60079 & n60082;
  assign n38840 = x169 & x194;
  assign n38841 = n38839 & n38840;
  assign n38842 = n38839 | n38840;
  assign n38843 = ~n38841 & n38842;
  assign n60083 = n38424 & n38843;
  assign n72404 = (n38843 & n59862) | (n38843 & n60083) | (n59862 & n60083);
  assign n72405 = (n38843 & n59861) | (n38843 & n60083) | (n59861 & n60083);
  assign n72406 = (n59580 & n72404) | (n59580 & n72405) | (n72404 & n72405);
  assign n60085 = n38424 | n38843;
  assign n72407 = n59862 | n60085;
  assign n72408 = n59861 | n60085;
  assign n72409 = (n59580 & n72407) | (n59580 & n72408) | (n72407 & n72408);
  assign n38846 = ~n72406 & n72409;
  assign n38847 = x168 & x195;
  assign n38848 = n38846 & n38847;
  assign n38849 = n38846 | n38847;
  assign n38850 = ~n38848 & n38849;
  assign n60044 = n38431 | n38433;
  assign n72410 = n38850 & n60044;
  assign n72359 = n38006 | n38431;
  assign n72360 = (n38431 & n38433) | (n38431 & n72359) | (n38433 & n72359);
  assign n72411 = n38850 & n72360;
  assign n72412 = (n59631 & n72410) | (n59631 & n72411) | (n72410 & n72411);
  assign n72413 = n38850 | n60044;
  assign n72414 = n38850 | n72360;
  assign n72415 = (n59631 & n72413) | (n59631 & n72414) | (n72413 & n72414);
  assign n38853 = ~n72412 & n72415;
  assign n38854 = x167 & x196;
  assign n38855 = n38853 & n38854;
  assign n38856 = n38853 | n38854;
  assign n38857 = ~n38855 & n38856;
  assign n60041 = n38438 | n38440;
  assign n60087 = n38857 & n60041;
  assign n60088 = n38438 & n38857;
  assign n60089 = (n72272 & n60087) | (n72272 & n60088) | (n60087 & n60088);
  assign n60090 = n38857 | n60041;
  assign n60091 = n38438 | n38857;
  assign n60092 = (n72272 & n60090) | (n72272 & n60091) | (n60090 & n60091);
  assign n38860 = ~n60089 & n60092;
  assign n38861 = x166 & x197;
  assign n38862 = n38860 & n38861;
  assign n38863 = n38860 | n38861;
  assign n38864 = ~n38862 & n38863;
  assign n60093 = n38445 & n38864;
  assign n72416 = (n38864 & n59872) | (n38864 & n60093) | (n59872 & n60093);
  assign n72417 = (n38864 & n59871) | (n38864 & n60093) | (n59871 & n60093);
  assign n72418 = (n59575 & n72416) | (n59575 & n72417) | (n72416 & n72417);
  assign n60095 = n38445 | n38864;
  assign n72419 = n59872 | n60095;
  assign n72420 = n59871 | n60095;
  assign n72421 = (n59575 & n72419) | (n59575 & n72420) | (n72419 & n72420);
  assign n38867 = ~n72418 & n72421;
  assign n38868 = x165 & x198;
  assign n38869 = n38867 & n38868;
  assign n38870 = n38867 | n38868;
  assign n38871 = ~n38869 & n38870;
  assign n60039 = n38452 | n38454;
  assign n72422 = n38871 & n60039;
  assign n72357 = n38027 | n38452;
  assign n72358 = (n38452 & n38454) | (n38452 & n72357) | (n38454 & n72357);
  assign n72423 = n38871 & n72358;
  assign n72424 = (n59641 & n72422) | (n59641 & n72423) | (n72422 & n72423);
  assign n72425 = n38871 | n60039;
  assign n72426 = n38871 | n72358;
  assign n72427 = (n59641 & n72425) | (n59641 & n72426) | (n72425 & n72426);
  assign n38874 = ~n72424 & n72427;
  assign n38875 = x164 & x199;
  assign n38876 = n38874 & n38875;
  assign n38877 = n38874 | n38875;
  assign n38878 = ~n38876 & n38877;
  assign n60036 = n38459 | n38461;
  assign n60097 = n38878 & n60036;
  assign n60098 = n38459 & n38878;
  assign n60099 = (n72267 & n60097) | (n72267 & n60098) | (n60097 & n60098);
  assign n60100 = n38878 | n60036;
  assign n60101 = n38459 | n38878;
  assign n60102 = (n72267 & n60100) | (n72267 & n60101) | (n60100 & n60101);
  assign n38881 = ~n60099 & n60102;
  assign n38882 = x163 & x200;
  assign n38883 = n38881 & n38882;
  assign n38884 = n38881 | n38882;
  assign n38885 = ~n38883 & n38884;
  assign n60103 = n38466 & n38885;
  assign n72428 = (n38885 & n59882) | (n38885 & n60103) | (n59882 & n60103);
  assign n72429 = (n38885 & n59881) | (n38885 & n60103) | (n59881 & n60103);
  assign n72430 = (n59570 & n72428) | (n59570 & n72429) | (n72428 & n72429);
  assign n60105 = n38466 | n38885;
  assign n72431 = n59882 | n60105;
  assign n72432 = n59881 | n60105;
  assign n72433 = (n59570 & n72431) | (n59570 & n72432) | (n72431 & n72432);
  assign n38888 = ~n72430 & n72433;
  assign n38889 = x162 & x201;
  assign n38890 = n38888 & n38889;
  assign n38891 = n38888 | n38889;
  assign n38892 = ~n38890 & n38891;
  assign n60034 = n38473 | n38475;
  assign n72434 = n38892 & n60034;
  assign n72355 = n38048 | n38473;
  assign n72356 = (n38473 & n38475) | (n38473 & n72355) | (n38475 & n72355);
  assign n72435 = n38892 & n72356;
  assign n72436 = (n59651 & n72434) | (n59651 & n72435) | (n72434 & n72435);
  assign n72437 = n38892 | n60034;
  assign n72438 = n38892 | n72356;
  assign n72439 = (n59651 & n72437) | (n59651 & n72438) | (n72437 & n72438);
  assign n38895 = ~n72436 & n72439;
  assign n38896 = x161 & x202;
  assign n38897 = n38895 & n38896;
  assign n38898 = n38895 | n38896;
  assign n38899 = ~n38897 & n38898;
  assign n60031 = n38480 | n38482;
  assign n60107 = n38899 & n60031;
  assign n60108 = n38480 & n38899;
  assign n60109 = (n72262 & n60107) | (n72262 & n60108) | (n60107 & n60108);
  assign n60110 = n38899 | n60031;
  assign n60111 = n38480 | n38899;
  assign n60112 = (n72262 & n60110) | (n72262 & n60111) | (n60110 & n60111);
  assign n38902 = ~n60109 & n60112;
  assign n38903 = x160 & x203;
  assign n38904 = n38902 & n38903;
  assign n38905 = n38902 | n38903;
  assign n38906 = ~n38904 & n38905;
  assign n60113 = n38487 & n38906;
  assign n72440 = (n38906 & n59892) | (n38906 & n60113) | (n59892 & n60113);
  assign n72441 = (n38906 & n59891) | (n38906 & n60113) | (n59891 & n60113);
  assign n72442 = (n72131 & n72440) | (n72131 & n72441) | (n72440 & n72441);
  assign n60115 = n38487 | n38906;
  assign n72443 = n59892 | n60115;
  assign n72444 = n59891 | n60115;
  assign n72445 = (n72131 & n72443) | (n72131 & n72444) | (n72443 & n72444);
  assign n38909 = ~n72442 & n72445;
  assign n38910 = x159 & x204;
  assign n38911 = n38909 & n38910;
  assign n38912 = n38909 | n38910;
  assign n38913 = ~n38911 & n38912;
  assign n38914 = n72354 & n38913;
  assign n38915 = n72354 | n38913;
  assign n38916 = ~n38914 & n38915;
  assign n38917 = x158 & x205;
  assign n38918 = n38916 & n38917;
  assign n38919 = n38916 | n38917;
  assign n38920 = ~n38918 & n38919;
  assign n60026 = n38501 | n38503;
  assign n60117 = n38920 & n60026;
  assign n60118 = n38501 & n38920;
  assign n60119 = (n72257 & n60117) | (n72257 & n60118) | (n60117 & n60118);
  assign n60120 = n38920 | n60026;
  assign n60121 = n38501 | n38920;
  assign n60122 = (n72257 & n60120) | (n72257 & n60121) | (n60120 & n60121);
  assign n38923 = ~n60119 & n60122;
  assign n38924 = x157 & x206;
  assign n38925 = n38923 & n38924;
  assign n38926 = n38923 | n38924;
  assign n38927 = ~n38925 & n38926;
  assign n60123 = n38508 & n38927;
  assign n72446 = (n38927 & n59902) | (n38927 & n60123) | (n59902 & n60123);
  assign n72447 = (n38927 & n59901) | (n38927 & n60123) | (n59901 & n60123);
  assign n72448 = (n72126 & n72446) | (n72126 & n72447) | (n72446 & n72447);
  assign n60125 = n38508 | n38927;
  assign n72449 = n59902 | n60125;
  assign n72450 = n59901 | n60125;
  assign n72451 = (n72126 & n72449) | (n72126 & n72450) | (n72449 & n72450);
  assign n38930 = ~n72448 & n72451;
  assign n38931 = x156 & x207;
  assign n38932 = n38930 & n38931;
  assign n38933 = n38930 | n38931;
  assign n38934 = ~n38932 & n38933;
  assign n38935 = n72349 & n38934;
  assign n38936 = n72349 | n38934;
  assign n38937 = ~n38935 & n38936;
  assign n38938 = x155 & x208;
  assign n38939 = n38937 & n38938;
  assign n38940 = n38937 | n38938;
  assign n38941 = ~n38939 & n38940;
  assign n60021 = n38522 | n38524;
  assign n60127 = n38941 & n60021;
  assign n60128 = n38522 & n38941;
  assign n60129 = (n59793 & n60127) | (n59793 & n60128) | (n60127 & n60128);
  assign n60130 = n38941 | n60021;
  assign n60131 = n38522 | n38941;
  assign n60132 = (n59793 & n60130) | (n59793 & n60131) | (n60130 & n60131);
  assign n38944 = ~n60129 & n60132;
  assign n38945 = x154 & x209;
  assign n38946 = n38944 & n38945;
  assign n38947 = n38944 | n38945;
  assign n38948 = ~n38946 & n38947;
  assign n60133 = n38529 & n38948;
  assign n60134 = (n38948 & n72329) | (n38948 & n60133) | (n72329 & n60133);
  assign n60135 = n38529 | n38948;
  assign n60136 = n72329 | n60135;
  assign n38951 = ~n60134 & n60136;
  assign n38952 = x153 & x210;
  assign n38953 = n38951 & n38952;
  assign n38954 = n38951 | n38952;
  assign n38955 = ~n38953 & n38954;
  assign n60137 = n38536 & n38955;
  assign n60138 = (n38955 & n59916) | (n38955 & n60137) | (n59916 & n60137);
  assign n60139 = n38536 | n38955;
  assign n60140 = n59916 | n60139;
  assign n38958 = ~n60138 & n60140;
  assign n38959 = x152 & x211;
  assign n38960 = n38958 & n38959;
  assign n38961 = n38958 | n38959;
  assign n38962 = ~n38960 & n38961;
  assign n60141 = n38543 & n38962;
  assign n60142 = (n38962 & n59920) | (n38962 & n60141) | (n59920 & n60141);
  assign n60143 = n38543 | n38962;
  assign n60144 = n59920 | n60143;
  assign n38965 = ~n60142 & n60144;
  assign n38966 = x151 & x212;
  assign n38967 = n38965 & n38966;
  assign n38968 = n38965 | n38966;
  assign n38969 = ~n38967 & n38968;
  assign n60145 = n38550 & n38969;
  assign n60146 = (n38969 & n59924) | (n38969 & n60145) | (n59924 & n60145);
  assign n60147 = n38550 | n38969;
  assign n60148 = n59924 | n60147;
  assign n38972 = ~n60146 & n60148;
  assign n38973 = x150 & x213;
  assign n38974 = n38972 & n38973;
  assign n38975 = n38972 | n38973;
  assign n38976 = ~n38974 & n38975;
  assign n60149 = n38557 & n38976;
  assign n60150 = (n38976 & n59928) | (n38976 & n60149) | (n59928 & n60149);
  assign n60151 = n38557 | n38976;
  assign n60152 = n59928 | n60151;
  assign n38979 = ~n60150 & n60152;
  assign n38980 = x149 & x214;
  assign n38981 = n38979 & n38980;
  assign n38982 = n38979 | n38980;
  assign n38983 = ~n38981 & n38982;
  assign n60153 = n38564 & n38983;
  assign n60154 = (n38983 & n59932) | (n38983 & n60153) | (n59932 & n60153);
  assign n60155 = n38564 | n38983;
  assign n60156 = n59932 | n60155;
  assign n38986 = ~n60154 & n60156;
  assign n38987 = x148 & x215;
  assign n38988 = n38986 & n38987;
  assign n38989 = n38986 | n38987;
  assign n38990 = ~n38988 & n38989;
  assign n60157 = n38571 & n38990;
  assign n60158 = (n38990 & n59936) | (n38990 & n60157) | (n59936 & n60157);
  assign n60159 = n38571 | n38990;
  assign n60160 = n59936 | n60159;
  assign n38993 = ~n60158 & n60160;
  assign n38994 = x147 & x216;
  assign n38995 = n38993 & n38994;
  assign n38996 = n38993 | n38994;
  assign n38997 = ~n38995 & n38996;
  assign n60161 = n38578 & n38997;
  assign n60162 = (n38997 & n59940) | (n38997 & n60161) | (n59940 & n60161);
  assign n60163 = n38578 | n38997;
  assign n60164 = n59940 | n60163;
  assign n39000 = ~n60162 & n60164;
  assign n39001 = x146 & x217;
  assign n39002 = n39000 & n39001;
  assign n39003 = n39000 | n39001;
  assign n39004 = ~n39002 & n39003;
  assign n60165 = n38585 & n39004;
  assign n60166 = (n39004 & n59944) | (n39004 & n60165) | (n59944 & n60165);
  assign n60167 = n38585 | n39004;
  assign n60168 = n59944 | n60167;
  assign n39007 = ~n60166 & n60168;
  assign n39008 = x145 & x218;
  assign n39009 = n39007 & n39008;
  assign n39010 = n39007 | n39008;
  assign n39011 = ~n39009 & n39010;
  assign n60169 = n38592 & n39011;
  assign n60170 = (n39011 & n59948) | (n39011 & n60169) | (n59948 & n60169);
  assign n60171 = n38592 | n39011;
  assign n60172 = n59948 | n60171;
  assign n39014 = ~n60170 & n60172;
  assign n39015 = x144 & x219;
  assign n39016 = n39014 & n39015;
  assign n39017 = n39014 | n39015;
  assign n39018 = ~n39016 & n39017;
  assign n60173 = n38599 & n39018;
  assign n60174 = (n39018 & n59952) | (n39018 & n60173) | (n59952 & n60173);
  assign n60175 = n38599 | n39018;
  assign n60176 = n59952 | n60175;
  assign n39021 = ~n60174 & n60176;
  assign n39022 = x143 & x220;
  assign n39023 = n39021 & n39022;
  assign n39024 = n39021 | n39022;
  assign n39025 = ~n39023 & n39024;
  assign n60177 = n38606 & n39025;
  assign n60178 = (n39025 & n59956) | (n39025 & n60177) | (n59956 & n60177);
  assign n60179 = n38606 | n39025;
  assign n60180 = n59956 | n60179;
  assign n39028 = ~n60178 & n60180;
  assign n39029 = x142 & x221;
  assign n39030 = n39028 & n39029;
  assign n39031 = n39028 | n39029;
  assign n39032 = ~n39030 & n39031;
  assign n60181 = n38613 & n39032;
  assign n60182 = (n39032 & n59960) | (n39032 & n60181) | (n59960 & n60181);
  assign n60183 = n38613 | n39032;
  assign n60184 = n59960 | n60183;
  assign n39035 = ~n60182 & n60184;
  assign n39036 = x141 & x222;
  assign n39037 = n39035 & n39036;
  assign n39038 = n39035 | n39036;
  assign n39039 = ~n39037 & n39038;
  assign n60185 = n38620 & n39039;
  assign n60186 = (n39039 & n59964) | (n39039 & n60185) | (n59964 & n60185);
  assign n60187 = n38620 | n39039;
  assign n60188 = n59964 | n60187;
  assign n39042 = ~n60186 & n60188;
  assign n39043 = x140 & x223;
  assign n39044 = n39042 & n39043;
  assign n39045 = n39042 | n39043;
  assign n39046 = ~n39044 & n39045;
  assign n60189 = n38627 & n39046;
  assign n60190 = (n39046 & n59968) | (n39046 & n60189) | (n59968 & n60189);
  assign n60191 = n38627 | n39046;
  assign n60192 = n59968 | n60191;
  assign n39049 = ~n60190 & n60192;
  assign n39050 = x139 & x224;
  assign n39051 = n39049 & n39050;
  assign n39052 = n39049 | n39050;
  assign n39053 = ~n39051 & n39052;
  assign n60193 = n38634 & n39053;
  assign n60194 = (n39053 & n59972) | (n39053 & n60193) | (n59972 & n60193);
  assign n60195 = n38634 | n39053;
  assign n60196 = n59972 | n60195;
  assign n39056 = ~n60194 & n60196;
  assign n39057 = x138 & x225;
  assign n39058 = n39056 & n39057;
  assign n39059 = n39056 | n39057;
  assign n39060 = ~n39058 & n39059;
  assign n60197 = n38641 & n39060;
  assign n60198 = (n39060 & n59976) | (n39060 & n60197) | (n59976 & n60197);
  assign n60199 = n38641 | n39060;
  assign n60200 = n59976 | n60199;
  assign n39063 = ~n60198 & n60200;
  assign n39064 = x137 & x226;
  assign n39065 = n39063 & n39064;
  assign n39066 = n39063 | n39064;
  assign n39067 = ~n39065 & n39066;
  assign n60201 = n38648 & n39067;
  assign n60202 = (n39067 & n59980) | (n39067 & n60201) | (n59980 & n60201);
  assign n60203 = n38648 | n39067;
  assign n60204 = n59980 | n60203;
  assign n39070 = ~n60202 & n60204;
  assign n39071 = x136 & x227;
  assign n39072 = n39070 & n39071;
  assign n39073 = n39070 | n39071;
  assign n39074 = ~n39072 & n39073;
  assign n60205 = n38655 & n39074;
  assign n60206 = (n39074 & n59984) | (n39074 & n60205) | (n59984 & n60205);
  assign n60207 = n38655 | n39074;
  assign n60208 = n59984 | n60207;
  assign n39077 = ~n60206 & n60208;
  assign n39078 = x135 & x228;
  assign n39079 = n39077 & n39078;
  assign n39080 = n39077 | n39078;
  assign n39081 = ~n39079 & n39080;
  assign n60209 = n38662 & n39081;
  assign n60210 = (n39081 & n59988) | (n39081 & n60209) | (n59988 & n60209);
  assign n60211 = n38662 | n39081;
  assign n60212 = n59988 | n60211;
  assign n39084 = ~n60210 & n60212;
  assign n39085 = x134 & x229;
  assign n39086 = n39084 & n39085;
  assign n39087 = n39084 | n39085;
  assign n39088 = ~n39086 & n39087;
  assign n60213 = n38669 & n39088;
  assign n60214 = (n39088 & n59992) | (n39088 & n60213) | (n59992 & n60213);
  assign n60215 = n38669 | n39088;
  assign n60216 = n59992 | n60215;
  assign n39091 = ~n60214 & n60216;
  assign n39092 = x133 & x230;
  assign n39093 = n39091 & n39092;
  assign n39094 = n39091 | n39092;
  assign n39095 = ~n39093 & n39094;
  assign n60217 = n38676 & n39095;
  assign n60218 = (n39095 & n59996) | (n39095 & n60217) | (n59996 & n60217);
  assign n60219 = n38676 | n39095;
  assign n60220 = n59996 | n60219;
  assign n39098 = ~n60218 & n60220;
  assign n39099 = x132 & x231;
  assign n39100 = n39098 & n39099;
  assign n39101 = n39098 | n39099;
  assign n39102 = ~n39100 & n39101;
  assign n60221 = n38683 & n39102;
  assign n60222 = (n39102 & n60000) | (n39102 & n60221) | (n60000 & n60221);
  assign n60223 = n38683 | n39102;
  assign n60224 = n60000 | n60223;
  assign n39105 = ~n60222 & n60224;
  assign n39106 = x131 & x232;
  assign n39107 = n39105 & n39106;
  assign n39108 = n39105 | n39106;
  assign n39109 = ~n39107 & n39108;
  assign n60225 = n38690 & n39109;
  assign n60226 = (n39109 & n60004) | (n39109 & n60225) | (n60004 & n60225);
  assign n60227 = n38690 | n39109;
  assign n60228 = n60004 | n60227;
  assign n39112 = ~n60226 & n60228;
  assign n39113 = x130 & x233;
  assign n39114 = n39112 & n39113;
  assign n39115 = n39112 | n39113;
  assign n39116 = ~n39114 & n39115;
  assign n60229 = n38697 & n39116;
  assign n60230 = (n39116 & n60009) | (n39116 & n60229) | (n60009 & n60229);
  assign n60231 = n38697 | n39116;
  assign n60232 = n60009 | n60231;
  assign n39119 = ~n60230 & n60232;
  assign n39120 = x129 & x234;
  assign n39121 = n39119 & n39120;
  assign n39122 = n39119 | n39120;
  assign n39123 = ~n39121 & n39122;
  assign n60019 = n38704 | n38706;
  assign n60233 = n39123 & n60019;
  assign n60234 = n38704 & n39123;
  assign n60235 = (n59788 & n60233) | (n59788 & n60234) | (n60233 & n60234);
  assign n60236 = n39123 | n60019;
  assign n60237 = n38704 | n39123;
  assign n60238 = (n59788 & n60236) | (n59788 & n60237) | (n60236 & n60237);
  assign n39126 = ~n60235 & n60238;
  assign n39127 = x128 & x235;
  assign n39128 = n39126 & n39127;
  assign n39129 = n39126 | n39127;
  assign n39130 = ~n39128 & n39129;
  assign n60017 = n38711 | n38713;
  assign n72452 = n39130 & n60017;
  assign n72453 = n38711 & n39130;
  assign n72454 = (n59786 & n72452) | (n59786 & n72453) | (n72452 & n72453);
  assign n72455 = n39130 | n60017;
  assign n72456 = n38711 | n39130;
  assign n72457 = (n59786 & n72455) | (n59786 & n72456) | (n72455 & n72456);
  assign n39133 = ~n72454 & n72457;
  assign n39134 = x127 & x236;
  assign n39135 = n39133 & n39134;
  assign n39136 = n39133 | n39134;
  assign n39137 = ~n39135 & n39136;
  assign n60015 = n38718 | n38720;
  assign n72458 = n39137 & n60015;
  assign n72459 = n38718 & n39137;
  assign n72460 = (n59784 & n72458) | (n59784 & n72459) | (n72458 & n72459);
  assign n72461 = n39137 | n60015;
  assign n72462 = n38718 | n39137;
  assign n72463 = (n59784 & n72461) | (n59784 & n72462) | (n72461 & n72462);
  assign n39140 = ~n72460 & n72463;
  assign n39141 = x126 & x237;
  assign n39142 = n39140 & n39141;
  assign n39143 = n39140 | n39141;
  assign n39144 = ~n39142 & n39143;
  assign n39145 = n60014 & n39144;
  assign n39146 = n60014 | n39144;
  assign n39147 = ~n39145 & n39146;
  assign n39148 = x125 & x238;
  assign n39149 = n39147 & n39148;
  assign n39150 = n39147 | n39148;
  assign n39151 = ~n39149 & n39150;
  assign n39152 = n38746 & n39151;
  assign n39153 = n38746 | n39151;
  assign n39154 = ~n39152 & n39153;
  assign n39155 = x124 & x239;
  assign n39156 = n39154 & n39155;
  assign n39157 = n39154 | n39155;
  assign n39158 = ~n39156 & n39157;
  assign n39159 = n38745 & n39158;
  assign n39160 = n38745 | n39158;
  assign n39161 = ~n39159 & n39160;
  assign n39162 = n39156 | n39159;
  assign n60239 = n39149 | n39151;
  assign n60240 = (n38746 & n39149) | (n38746 & n60239) | (n39149 & n60239);
  assign n60016 = (n38718 & n59784) | (n38718 & n60015) | (n59784 & n60015);
  assign n60018 = (n38711 & n59786) | (n38711 & n60017) | (n59786 & n60017);
  assign n60253 = n38925 | n38927;
  assign n72466 = n38508 | n38925;
  assign n72467 = (n38925 & n38927) | (n38925 & n72466) | (n38927 & n72466);
  assign n72468 = (n59902 & n60253) | (n59902 & n72467) | (n60253 & n72467);
  assign n72469 = (n59901 & n60253) | (n59901 & n72467) | (n60253 & n72467);
  assign n72470 = (n72126 & n72468) | (n72126 & n72469) | (n72468 & n72469);
  assign n60258 = n38904 | n38906;
  assign n72471 = n38487 | n38904;
  assign n72472 = (n38904 & n38906) | (n38904 & n72471) | (n38906 & n72471);
  assign n72473 = (n59892 & n60258) | (n59892 & n72472) | (n60258 & n72472);
  assign n72474 = (n59891 & n60258) | (n59891 & n72472) | (n60258 & n72472);
  assign n72475 = (n72131 & n72473) | (n72131 & n72474) | (n72473 & n72474);
  assign n60035 = (n59651 & n72356) | (n59651 & n60034) | (n72356 & n60034);
  assign n60263 = n38883 | n38885;
  assign n72476 = n38466 | n38883;
  assign n72477 = (n38883 & n38885) | (n38883 & n72476) | (n38885 & n72476);
  assign n72478 = (n59882 & n60263) | (n59882 & n72477) | (n60263 & n72477);
  assign n72479 = (n59881 & n60263) | (n59881 & n72477) | (n60263 & n72477);
  assign n72480 = (n59570 & n72478) | (n59570 & n72479) | (n72478 & n72479);
  assign n60040 = (n59641 & n72358) | (n59641 & n60039) | (n72358 & n60039);
  assign n60268 = n38862 | n38864;
  assign n72481 = n38445 | n38862;
  assign n72482 = (n38862 & n38864) | (n38862 & n72481) | (n38864 & n72481);
  assign n72483 = (n59872 & n60268) | (n59872 & n72482) | (n60268 & n72482);
  assign n72484 = (n59871 & n60268) | (n59871 & n72482) | (n60268 & n72482);
  assign n72485 = (n59575 & n72483) | (n59575 & n72484) | (n72483 & n72484);
  assign n60045 = (n59631 & n72360) | (n59631 & n60044) | (n72360 & n60044);
  assign n60273 = n38841 | n38843;
  assign n72486 = n38424 | n38841;
  assign n72487 = (n38841 & n38843) | (n38841 & n72486) | (n38843 & n72486);
  assign n72488 = (n59862 & n60273) | (n59862 & n72487) | (n60273 & n72487);
  assign n72489 = (n59861 & n60273) | (n59861 & n72487) | (n60273 & n72487);
  assign n72490 = (n59580 & n72488) | (n59580 & n72489) | (n72488 & n72489);
  assign n60050 = (n59621 & n72362) | (n59621 & n60049) | (n72362 & n60049);
  assign n60278 = n38820 | n38822;
  assign n72491 = n38403 | n38820;
  assign n72492 = (n38820 & n38822) | (n38820 & n72491) | (n38822 & n72491);
  assign n72493 = (n59851 & n60278) | (n59851 & n72492) | (n60278 & n72492);
  assign n72494 = (n59852 & n60278) | (n59852 & n72492) | (n60278 & n72492);
  assign n72495 = (n59585 & n72493) | (n59585 & n72494) | (n72493 & n72494);
  assign n39214 = x175 & x189;
  assign n72498 = n39214 & n72378;
  assign n72499 = (n38801 & n39214) | (n38801 & n72498) | (n39214 & n72498);
  assign n60288 = n39214 & n72378;
  assign n60289 = (n72371 & n72499) | (n72371 & n60288) | (n72499 & n60288);
  assign n72500 = n39214 | n72378;
  assign n72501 = n38801 | n72500;
  assign n60291 = n39214 | n72378;
  assign n60292 = (n72371 & n72501) | (n72371 & n60291) | (n72501 & n60291);
  assign n39217 = ~n60289 & n60292;
  assign n60283 = n38806 | n60067;
  assign n72502 = n39217 & n60283;
  assign n72496 = n38389 | n38806;
  assign n72497 = (n38806 & n38808) | (n38806 & n72496) | (n38808 & n72496);
  assign n72503 = n39217 & n72497;
  assign n72504 = (n72284 & n72502) | (n72284 & n72503) | (n72502 & n72503);
  assign n72505 = n39217 | n60283;
  assign n72506 = n39217 | n72497;
  assign n72507 = (n72284 & n72505) | (n72284 & n72506) | (n72505 & n72506);
  assign n39220 = ~n72504 & n72507;
  assign n39221 = x174 & x190;
  assign n39222 = n39220 & n39221;
  assign n39223 = n39220 | n39221;
  assign n39224 = ~n39222 & n39223;
  assign n60280 = n38813 | n38815;
  assign n60293 = n39224 & n60280;
  assign n60294 = n38813 & n39224;
  assign n72508 = (n60052 & n60293) | (n60052 & n60294) | (n60293 & n60294);
  assign n72509 = (n60293 & n60294) | (n60293 & n72364) | (n60294 & n72364);
  assign n72510 = (n59588 & n72508) | (n59588 & n72509) | (n72508 & n72509);
  assign n60296 = n39224 | n60280;
  assign n60297 = n38813 | n39224;
  assign n72511 = (n60052 & n60296) | (n60052 & n60297) | (n60296 & n60297);
  assign n72512 = (n60296 & n60297) | (n60296 & n72364) | (n60297 & n72364);
  assign n72513 = (n59588 & n72511) | (n59588 & n72512) | (n72511 & n72512);
  assign n39227 = ~n72510 & n72513;
  assign n39228 = x173 & x191;
  assign n39229 = n39227 & n39228;
  assign n39230 = n39227 | n39228;
  assign n39231 = ~n39229 & n39230;
  assign n39232 = n72495 & n39231;
  assign n39233 = n72495 | n39231;
  assign n39234 = ~n39232 & n39233;
  assign n39235 = x172 & x192;
  assign n39236 = n39234 & n39235;
  assign n39237 = n39234 | n39235;
  assign n39238 = ~n39236 & n39237;
  assign n60275 = n38827 | n38829;
  assign n60299 = n39238 & n60275;
  assign n60300 = n38827 & n39238;
  assign n60301 = (n60050 & n60299) | (n60050 & n60300) | (n60299 & n60300);
  assign n60302 = n39238 | n60275;
  assign n60303 = n38827 | n39238;
  assign n60304 = (n60050 & n60302) | (n60050 & n60303) | (n60302 & n60303);
  assign n39241 = ~n60301 & n60304;
  assign n39242 = x171 & x193;
  assign n39243 = n39241 & n39242;
  assign n39244 = n39241 | n39242;
  assign n39245 = ~n39243 & n39244;
  assign n60305 = n38834 & n39245;
  assign n60306 = (n39245 & n60079) | (n39245 & n60305) | (n60079 & n60305);
  assign n60307 = n38834 | n39245;
  assign n60308 = n60079 | n60307;
  assign n39248 = ~n60306 & n60308;
  assign n39249 = x170 & x194;
  assign n39250 = n39248 & n39249;
  assign n39251 = n39248 | n39249;
  assign n39252 = ~n39250 & n39251;
  assign n39253 = n72490 & n39252;
  assign n39254 = n72490 | n39252;
  assign n39255 = ~n39253 & n39254;
  assign n39256 = x169 & x195;
  assign n39257 = n39255 & n39256;
  assign n39258 = n39255 | n39256;
  assign n39259 = ~n39257 & n39258;
  assign n60270 = n38848 | n38850;
  assign n60309 = n39259 & n60270;
  assign n60310 = n38848 & n39259;
  assign n60311 = (n60045 & n60309) | (n60045 & n60310) | (n60309 & n60310);
  assign n60312 = n39259 | n60270;
  assign n60313 = n38848 | n39259;
  assign n60314 = (n60045 & n60312) | (n60045 & n60313) | (n60312 & n60313);
  assign n39262 = ~n60311 & n60314;
  assign n39263 = x168 & x196;
  assign n39264 = n39262 & n39263;
  assign n39265 = n39262 | n39263;
  assign n39266 = ~n39264 & n39265;
  assign n60315 = n38855 & n39266;
  assign n60316 = (n39266 & n60089) | (n39266 & n60315) | (n60089 & n60315);
  assign n60317 = n38855 | n39266;
  assign n60318 = n60089 | n60317;
  assign n39269 = ~n60316 & n60318;
  assign n39270 = x167 & x197;
  assign n39271 = n39269 & n39270;
  assign n39272 = n39269 | n39270;
  assign n39273 = ~n39271 & n39272;
  assign n39274 = n72485 & n39273;
  assign n39275 = n72485 | n39273;
  assign n39276 = ~n39274 & n39275;
  assign n39277 = x166 & x198;
  assign n39278 = n39276 & n39277;
  assign n39279 = n39276 | n39277;
  assign n39280 = ~n39278 & n39279;
  assign n60265 = n38869 | n38871;
  assign n60319 = n39280 & n60265;
  assign n60320 = n38869 & n39280;
  assign n60321 = (n60040 & n60319) | (n60040 & n60320) | (n60319 & n60320);
  assign n60322 = n39280 | n60265;
  assign n60323 = n38869 | n39280;
  assign n60324 = (n60040 & n60322) | (n60040 & n60323) | (n60322 & n60323);
  assign n39283 = ~n60321 & n60324;
  assign n39284 = x165 & x199;
  assign n39285 = n39283 & n39284;
  assign n39286 = n39283 | n39284;
  assign n39287 = ~n39285 & n39286;
  assign n60325 = n38876 & n39287;
  assign n60326 = (n39287 & n60099) | (n39287 & n60325) | (n60099 & n60325);
  assign n60327 = n38876 | n39287;
  assign n60328 = n60099 | n60327;
  assign n39290 = ~n60326 & n60328;
  assign n39291 = x164 & x200;
  assign n39292 = n39290 & n39291;
  assign n39293 = n39290 | n39291;
  assign n39294 = ~n39292 & n39293;
  assign n39295 = n72480 & n39294;
  assign n39296 = n72480 | n39294;
  assign n39297 = ~n39295 & n39296;
  assign n39298 = x163 & x201;
  assign n39299 = n39297 & n39298;
  assign n39300 = n39297 | n39298;
  assign n39301 = ~n39299 & n39300;
  assign n60260 = n38890 | n38892;
  assign n60329 = n39301 & n60260;
  assign n60330 = n38890 & n39301;
  assign n60331 = (n60035 & n60329) | (n60035 & n60330) | (n60329 & n60330);
  assign n60332 = n39301 | n60260;
  assign n60333 = n38890 | n39301;
  assign n60334 = (n60035 & n60332) | (n60035 & n60333) | (n60332 & n60333);
  assign n39304 = ~n60331 & n60334;
  assign n39305 = x162 & x202;
  assign n39306 = n39304 & n39305;
  assign n39307 = n39304 | n39305;
  assign n39308 = ~n39306 & n39307;
  assign n60335 = n38897 & n39308;
  assign n60336 = (n39308 & n60109) | (n39308 & n60335) | (n60109 & n60335);
  assign n60337 = n38897 | n39308;
  assign n60338 = n60109 | n60337;
  assign n39311 = ~n60336 & n60338;
  assign n39312 = x161 & x203;
  assign n39313 = n39311 & n39312;
  assign n39314 = n39311 | n39312;
  assign n39315 = ~n39313 & n39314;
  assign n39316 = n72475 & n39315;
  assign n39317 = n72475 | n39315;
  assign n39318 = ~n39316 & n39317;
  assign n39319 = x160 & x204;
  assign n39320 = n39318 & n39319;
  assign n39321 = n39318 | n39319;
  assign n39322 = ~n39320 & n39321;
  assign n60255 = n38911 | n38913;
  assign n60339 = n39322 & n60255;
  assign n60340 = n38911 & n39322;
  assign n60341 = (n72354 & n60339) | (n72354 & n60340) | (n60339 & n60340);
  assign n60342 = n39322 | n60255;
  assign n60343 = n38911 | n39322;
  assign n60344 = (n72354 & n60342) | (n72354 & n60343) | (n60342 & n60343);
  assign n39325 = ~n60341 & n60344;
  assign n39326 = x159 & x205;
  assign n39327 = n39325 & n39326;
  assign n39328 = n39325 | n39326;
  assign n39329 = ~n39327 & n39328;
  assign n60345 = n38918 & n39329;
  assign n72514 = (n39329 & n60118) | (n39329 & n60345) | (n60118 & n60345);
  assign n72515 = (n39329 & n60117) | (n39329 & n60345) | (n60117 & n60345);
  assign n72516 = (n72257 & n72514) | (n72257 & n72515) | (n72514 & n72515);
  assign n60347 = n38918 | n39329;
  assign n72517 = n60118 | n60347;
  assign n72518 = n60117 | n60347;
  assign n72519 = (n72257 & n72517) | (n72257 & n72518) | (n72517 & n72518);
  assign n39332 = ~n72516 & n72519;
  assign n39333 = x158 & x206;
  assign n39334 = n39332 & n39333;
  assign n39335 = n39332 | n39333;
  assign n39336 = ~n39334 & n39335;
  assign n39337 = n72470 & n39336;
  assign n39338 = n72470 | n39336;
  assign n39339 = ~n39337 & n39338;
  assign n39340 = x157 & x207;
  assign n39341 = n39339 & n39340;
  assign n39342 = n39339 | n39340;
  assign n39343 = ~n39341 & n39342;
  assign n60250 = n38932 | n38934;
  assign n60349 = n39343 & n60250;
  assign n60350 = n38932 & n39343;
  assign n60351 = (n72349 & n60349) | (n72349 & n60350) | (n60349 & n60350);
  assign n60352 = n39343 | n60250;
  assign n60353 = n38932 | n39343;
  assign n60354 = (n72349 & n60352) | (n72349 & n60353) | (n60352 & n60353);
  assign n39346 = ~n60351 & n60354;
  assign n39347 = x156 & x208;
  assign n39348 = n39346 & n39347;
  assign n39349 = n39346 | n39347;
  assign n39350 = ~n39348 & n39349;
  assign n60355 = n38939 & n39350;
  assign n72520 = (n39350 & n60128) | (n39350 & n60355) | (n60128 & n60355);
  assign n72521 = (n39350 & n60127) | (n39350 & n60355) | (n60127 & n60355);
  assign n72522 = (n59793 & n72520) | (n59793 & n72521) | (n72520 & n72521);
  assign n60357 = n38939 | n39350;
  assign n72523 = n60128 | n60357;
  assign n72524 = n60127 | n60357;
  assign n72525 = (n59793 & n72523) | (n59793 & n72524) | (n72523 & n72524);
  assign n39353 = ~n72522 & n72525;
  assign n39354 = x155 & x209;
  assign n39355 = n39353 & n39354;
  assign n39356 = n39353 | n39354;
  assign n39357 = ~n39355 & n39356;
  assign n60248 = n38946 | n38948;
  assign n72526 = n39357 & n60248;
  assign n72464 = n38529 | n38946;
  assign n72465 = (n38946 & n38948) | (n38946 & n72464) | (n38948 & n72464);
  assign n72527 = n39357 & n72465;
  assign n72528 = (n72329 & n72526) | (n72329 & n72527) | (n72526 & n72527);
  assign n72529 = n39357 | n60248;
  assign n72530 = n39357 | n72465;
  assign n72531 = (n72329 & n72529) | (n72329 & n72530) | (n72529 & n72530);
  assign n39360 = ~n72528 & n72531;
  assign n39361 = x154 & x210;
  assign n39362 = n39360 & n39361;
  assign n39363 = n39360 | n39361;
  assign n39364 = ~n39362 & n39363;
  assign n60359 = n38953 & n39364;
  assign n72532 = (n39364 & n60137) | (n39364 & n60359) | (n60137 & n60359);
  assign n72533 = (n38955 & n39364) | (n38955 & n60359) | (n39364 & n60359);
  assign n72534 = (n59916 & n72532) | (n59916 & n72533) | (n72532 & n72533);
  assign n60361 = n38953 | n39364;
  assign n72535 = n60137 | n60361;
  assign n72536 = n38955 | n60361;
  assign n72537 = (n59916 & n72535) | (n59916 & n72536) | (n72535 & n72536);
  assign n39367 = ~n72534 & n72537;
  assign n39368 = x153 & x211;
  assign n39369 = n39367 & n39368;
  assign n39370 = n39367 | n39368;
  assign n39371 = ~n39369 & n39370;
  assign n60363 = n38960 & n39371;
  assign n60364 = (n39371 & n60142) | (n39371 & n60363) | (n60142 & n60363);
  assign n60365 = n38960 | n39371;
  assign n60366 = n60142 | n60365;
  assign n39374 = ~n60364 & n60366;
  assign n39375 = x152 & x212;
  assign n39376 = n39374 & n39375;
  assign n39377 = n39374 | n39375;
  assign n39378 = ~n39376 & n39377;
  assign n60367 = n38967 & n39378;
  assign n60368 = (n39378 & n60146) | (n39378 & n60367) | (n60146 & n60367);
  assign n60369 = n38967 | n39378;
  assign n60370 = n60146 | n60369;
  assign n39381 = ~n60368 & n60370;
  assign n39382 = x151 & x213;
  assign n39383 = n39381 & n39382;
  assign n39384 = n39381 | n39382;
  assign n39385 = ~n39383 & n39384;
  assign n60371 = n38974 & n39385;
  assign n60372 = (n39385 & n60150) | (n39385 & n60371) | (n60150 & n60371);
  assign n60373 = n38974 | n39385;
  assign n60374 = n60150 | n60373;
  assign n39388 = ~n60372 & n60374;
  assign n39389 = x150 & x214;
  assign n39390 = n39388 & n39389;
  assign n39391 = n39388 | n39389;
  assign n39392 = ~n39390 & n39391;
  assign n60375 = n38981 & n39392;
  assign n60376 = (n39392 & n60154) | (n39392 & n60375) | (n60154 & n60375);
  assign n60377 = n38981 | n39392;
  assign n60378 = n60154 | n60377;
  assign n39395 = ~n60376 & n60378;
  assign n39396 = x149 & x215;
  assign n39397 = n39395 & n39396;
  assign n39398 = n39395 | n39396;
  assign n39399 = ~n39397 & n39398;
  assign n60379 = n38988 & n39399;
  assign n60380 = (n39399 & n60158) | (n39399 & n60379) | (n60158 & n60379);
  assign n60381 = n38988 | n39399;
  assign n60382 = n60158 | n60381;
  assign n39402 = ~n60380 & n60382;
  assign n39403 = x148 & x216;
  assign n39404 = n39402 & n39403;
  assign n39405 = n39402 | n39403;
  assign n39406 = ~n39404 & n39405;
  assign n60383 = n38995 & n39406;
  assign n60384 = (n39406 & n60162) | (n39406 & n60383) | (n60162 & n60383);
  assign n60385 = n38995 | n39406;
  assign n60386 = n60162 | n60385;
  assign n39409 = ~n60384 & n60386;
  assign n39410 = x147 & x217;
  assign n39411 = n39409 & n39410;
  assign n39412 = n39409 | n39410;
  assign n39413 = ~n39411 & n39412;
  assign n60387 = n39002 & n39413;
  assign n60388 = (n39413 & n60166) | (n39413 & n60387) | (n60166 & n60387);
  assign n60389 = n39002 | n39413;
  assign n60390 = n60166 | n60389;
  assign n39416 = ~n60388 & n60390;
  assign n39417 = x146 & x218;
  assign n39418 = n39416 & n39417;
  assign n39419 = n39416 | n39417;
  assign n39420 = ~n39418 & n39419;
  assign n60391 = n39009 & n39420;
  assign n60392 = (n39420 & n60170) | (n39420 & n60391) | (n60170 & n60391);
  assign n60393 = n39009 | n39420;
  assign n60394 = n60170 | n60393;
  assign n39423 = ~n60392 & n60394;
  assign n39424 = x145 & x219;
  assign n39425 = n39423 & n39424;
  assign n39426 = n39423 | n39424;
  assign n39427 = ~n39425 & n39426;
  assign n60395 = n39016 & n39427;
  assign n60396 = (n39427 & n60174) | (n39427 & n60395) | (n60174 & n60395);
  assign n60397 = n39016 | n39427;
  assign n60398 = n60174 | n60397;
  assign n39430 = ~n60396 & n60398;
  assign n39431 = x144 & x220;
  assign n39432 = n39430 & n39431;
  assign n39433 = n39430 | n39431;
  assign n39434 = ~n39432 & n39433;
  assign n60399 = n39023 & n39434;
  assign n60400 = (n39434 & n60178) | (n39434 & n60399) | (n60178 & n60399);
  assign n60401 = n39023 | n39434;
  assign n60402 = n60178 | n60401;
  assign n39437 = ~n60400 & n60402;
  assign n39438 = x143 & x221;
  assign n39439 = n39437 & n39438;
  assign n39440 = n39437 | n39438;
  assign n39441 = ~n39439 & n39440;
  assign n60403 = n39030 & n39441;
  assign n60404 = (n39441 & n60182) | (n39441 & n60403) | (n60182 & n60403);
  assign n60405 = n39030 | n39441;
  assign n60406 = n60182 | n60405;
  assign n39444 = ~n60404 & n60406;
  assign n39445 = x142 & x222;
  assign n39446 = n39444 & n39445;
  assign n39447 = n39444 | n39445;
  assign n39448 = ~n39446 & n39447;
  assign n60407 = n39037 & n39448;
  assign n60408 = (n39448 & n60186) | (n39448 & n60407) | (n60186 & n60407);
  assign n60409 = n39037 | n39448;
  assign n60410 = n60186 | n60409;
  assign n39451 = ~n60408 & n60410;
  assign n39452 = x141 & x223;
  assign n39453 = n39451 & n39452;
  assign n39454 = n39451 | n39452;
  assign n39455 = ~n39453 & n39454;
  assign n60411 = n39044 & n39455;
  assign n60412 = (n39455 & n60190) | (n39455 & n60411) | (n60190 & n60411);
  assign n60413 = n39044 | n39455;
  assign n60414 = n60190 | n60413;
  assign n39458 = ~n60412 & n60414;
  assign n39459 = x140 & x224;
  assign n39460 = n39458 & n39459;
  assign n39461 = n39458 | n39459;
  assign n39462 = ~n39460 & n39461;
  assign n60415 = n39051 & n39462;
  assign n60416 = (n39462 & n60194) | (n39462 & n60415) | (n60194 & n60415);
  assign n60417 = n39051 | n39462;
  assign n60418 = n60194 | n60417;
  assign n39465 = ~n60416 & n60418;
  assign n39466 = x139 & x225;
  assign n39467 = n39465 & n39466;
  assign n39468 = n39465 | n39466;
  assign n39469 = ~n39467 & n39468;
  assign n60419 = n39058 & n39469;
  assign n60420 = (n39469 & n60198) | (n39469 & n60419) | (n60198 & n60419);
  assign n60421 = n39058 | n39469;
  assign n60422 = n60198 | n60421;
  assign n39472 = ~n60420 & n60422;
  assign n39473 = x138 & x226;
  assign n39474 = n39472 & n39473;
  assign n39475 = n39472 | n39473;
  assign n39476 = ~n39474 & n39475;
  assign n60423 = n39065 & n39476;
  assign n60424 = (n39476 & n60202) | (n39476 & n60423) | (n60202 & n60423);
  assign n60425 = n39065 | n39476;
  assign n60426 = n60202 | n60425;
  assign n39479 = ~n60424 & n60426;
  assign n39480 = x137 & x227;
  assign n39481 = n39479 & n39480;
  assign n39482 = n39479 | n39480;
  assign n39483 = ~n39481 & n39482;
  assign n60427 = n39072 & n39483;
  assign n60428 = (n39483 & n60206) | (n39483 & n60427) | (n60206 & n60427);
  assign n60429 = n39072 | n39483;
  assign n60430 = n60206 | n60429;
  assign n39486 = ~n60428 & n60430;
  assign n39487 = x136 & x228;
  assign n39488 = n39486 & n39487;
  assign n39489 = n39486 | n39487;
  assign n39490 = ~n39488 & n39489;
  assign n60431 = n39079 & n39490;
  assign n60432 = (n39490 & n60210) | (n39490 & n60431) | (n60210 & n60431);
  assign n60433 = n39079 | n39490;
  assign n60434 = n60210 | n60433;
  assign n39493 = ~n60432 & n60434;
  assign n39494 = x135 & x229;
  assign n39495 = n39493 & n39494;
  assign n39496 = n39493 | n39494;
  assign n39497 = ~n39495 & n39496;
  assign n60435 = n39086 & n39497;
  assign n60436 = (n39497 & n60214) | (n39497 & n60435) | (n60214 & n60435);
  assign n60437 = n39086 | n39497;
  assign n60438 = n60214 | n60437;
  assign n39500 = ~n60436 & n60438;
  assign n39501 = x134 & x230;
  assign n39502 = n39500 & n39501;
  assign n39503 = n39500 | n39501;
  assign n39504 = ~n39502 & n39503;
  assign n60439 = n39093 & n39504;
  assign n60440 = (n39504 & n60218) | (n39504 & n60439) | (n60218 & n60439);
  assign n60441 = n39093 | n39504;
  assign n60442 = n60218 | n60441;
  assign n39507 = ~n60440 & n60442;
  assign n39508 = x133 & x231;
  assign n39509 = n39507 & n39508;
  assign n39510 = n39507 | n39508;
  assign n39511 = ~n39509 & n39510;
  assign n60443 = n39100 & n39511;
  assign n60444 = (n39511 & n60222) | (n39511 & n60443) | (n60222 & n60443);
  assign n60445 = n39100 | n39511;
  assign n60446 = n60222 | n60445;
  assign n39514 = ~n60444 & n60446;
  assign n39515 = x132 & x232;
  assign n39516 = n39514 & n39515;
  assign n39517 = n39514 | n39515;
  assign n39518 = ~n39516 & n39517;
  assign n60447 = n39107 & n39518;
  assign n60448 = (n39518 & n60226) | (n39518 & n60447) | (n60226 & n60447);
  assign n60449 = n39107 | n39518;
  assign n60450 = n60226 | n60449;
  assign n39521 = ~n60448 & n60450;
  assign n39522 = x131 & x233;
  assign n39523 = n39521 & n39522;
  assign n39524 = n39521 | n39522;
  assign n39525 = ~n39523 & n39524;
  assign n60451 = n39114 & n39525;
  assign n60452 = (n39525 & n60230) | (n39525 & n60451) | (n60230 & n60451);
  assign n60453 = n39114 | n39525;
  assign n60454 = n60230 | n60453;
  assign n39528 = ~n60452 & n60454;
  assign n39529 = x130 & x234;
  assign n39530 = n39528 & n39529;
  assign n39531 = n39528 | n39529;
  assign n39532 = ~n39530 & n39531;
  assign n60455 = n39121 & n39532;
  assign n60456 = (n39532 & n60235) | (n39532 & n60455) | (n60235 & n60455);
  assign n60457 = n39121 | n39532;
  assign n60458 = n60235 | n60457;
  assign n39535 = ~n60456 & n60458;
  assign n39536 = x129 & x235;
  assign n39537 = n39535 & n39536;
  assign n39538 = n39535 | n39536;
  assign n39539 = ~n39537 & n39538;
  assign n60245 = n39128 | n39130;
  assign n60459 = n39539 & n60245;
  assign n60460 = n39128 & n39539;
  assign n60461 = (n60018 & n60459) | (n60018 & n60460) | (n60459 & n60460);
  assign n60462 = n39539 | n60245;
  assign n60463 = n39128 | n39539;
  assign n60464 = (n60018 & n60462) | (n60018 & n60463) | (n60462 & n60463);
  assign n39542 = ~n60461 & n60464;
  assign n39543 = x128 & x236;
  assign n39544 = n39542 & n39543;
  assign n39545 = n39542 | n39543;
  assign n39546 = ~n39544 & n39545;
  assign n60243 = n39135 | n39137;
  assign n72538 = n39546 & n60243;
  assign n72539 = n39135 & n39546;
  assign n72540 = (n60016 & n72538) | (n60016 & n72539) | (n72538 & n72539);
  assign n72541 = n39546 | n60243;
  assign n72542 = n39135 | n39546;
  assign n72543 = (n60016 & n72541) | (n60016 & n72542) | (n72541 & n72542);
  assign n39549 = ~n72540 & n72543;
  assign n39550 = x127 & x237;
  assign n39551 = n39549 & n39550;
  assign n39552 = n39549 | n39550;
  assign n39553 = ~n39551 & n39552;
  assign n60241 = n39142 | n39144;
  assign n72544 = n39553 & n60241;
  assign n72545 = n39142 & n39553;
  assign n72546 = (n60014 & n72544) | (n60014 & n72545) | (n72544 & n72545);
  assign n72547 = n39553 | n60241;
  assign n72548 = n39142 | n39553;
  assign n72549 = (n60014 & n72547) | (n60014 & n72548) | (n72547 & n72548);
  assign n39556 = ~n72546 & n72549;
  assign n39557 = x126 & x238;
  assign n39558 = n39556 & n39557;
  assign n39559 = n39556 | n39557;
  assign n39560 = ~n39558 & n39559;
  assign n39561 = n60240 & n39560;
  assign n39562 = n60240 | n39560;
  assign n39563 = ~n39561 & n39562;
  assign n39564 = x125 & x239;
  assign n39565 = n39563 & n39564;
  assign n39566 = n39563 | n39564;
  assign n39567 = ~n39565 & n39566;
  assign n39568 = n39162 & n39567;
  assign n39569 = n39162 | n39567;
  assign n39570 = ~n39568 & n39569;
  assign n60465 = n39565 | n39567;
  assign n60466 = (n39162 & n39565) | (n39162 & n60465) | (n39565 & n60465);
  assign n60242 = (n39142 & n60014) | (n39142 & n60241) | (n60014 & n60241);
  assign n60244 = (n39135 & n60016) | (n39135 & n60243) | (n60016 & n60243);
  assign n60249 = (n72329 & n72465) | (n72329 & n60248) | (n72465 & n60248);
  assign n60476 = n39348 | n39350;
  assign n72550 = n38939 | n39348;
  assign n72551 = (n39348 & n39350) | (n39348 & n72550) | (n39350 & n72550);
  assign n72552 = (n60128 & n60476) | (n60128 & n72551) | (n60476 & n72551);
  assign n72553 = (n60127 & n60476) | (n60127 & n72551) | (n60476 & n72551);
  assign n72554 = (n59793 & n72552) | (n59793 & n72553) | (n72552 & n72553);
  assign n60481 = n39327 | n39329;
  assign n72555 = n38918 | n39327;
  assign n72556 = (n39327 & n39329) | (n39327 & n72555) | (n39329 & n72555);
  assign n72557 = (n60118 & n60481) | (n60118 & n72556) | (n60481 & n72556);
  assign n72558 = (n60117 & n60481) | (n60117 & n72556) | (n60481 & n72556);
  assign n72559 = (n72257 & n72557) | (n72257 & n72558) | (n72557 & n72558);
  assign n72568 = n38813 | n39222;
  assign n72569 = (n39222 & n39224) | (n39222 & n72568) | (n39224 & n72568);
  assign n72570 = n39222 | n39224;
  assign n72571 = (n39222 & n60280) | (n39222 & n72570) | (n60280 & n72570);
  assign n72572 = (n60052 & n72569) | (n60052 & n72571) | (n72569 & n72571);
  assign n72573 = (n72364 & n72569) | (n72364 & n72571) | (n72569 & n72571);
  assign n72574 = (n59588 & n72572) | (n59588 & n72573) | (n72572 & n72573);
  assign n39622 = x175 & x190;
  assign n72576 = n39622 & n72499;
  assign n72577 = n39622 & n60288;
  assign n72578 = (n72371 & n72576) | (n72371 & n72577) | (n72576 & n72577);
  assign n72575 = (n39217 & n39622) | (n39217 & n72578) | (n39622 & n72578);
  assign n72579 = (n60283 & n72575) | (n60283 & n72578) | (n72575 & n72578);
  assign n72580 = (n72497 & n72575) | (n72497 & n72578) | (n72575 & n72578);
  assign n72581 = (n72284 & n72579) | (n72284 & n72580) | (n72579 & n72580);
  assign n72583 = n39622 | n72499;
  assign n72584 = n39622 | n60288;
  assign n72585 = (n72371 & n72583) | (n72371 & n72584) | (n72583 & n72584);
  assign n72582 = n39217 | n72585;
  assign n72586 = (n60283 & n72582) | (n60283 & n72585) | (n72582 & n72585);
  assign n72587 = (n72497 & n72582) | (n72497 & n72585) | (n72582 & n72585);
  assign n72588 = (n72284 & n72586) | (n72284 & n72587) | (n72586 & n72587);
  assign n39625 = ~n72581 & n72588;
  assign n39626 = n72574 & n39625;
  assign n39627 = n72574 | n39625;
  assign n39628 = ~n39626 & n39627;
  assign n39629 = x174 & x191;
  assign n39630 = n39628 & n39629;
  assign n39631 = n39628 | n39629;
  assign n39632 = ~n39630 & n39631;
  assign n60503 = n39229 | n39231;
  assign n60516 = n39632 & n60503;
  assign n60517 = n39229 & n39632;
  assign n60518 = (n72495 & n60516) | (n72495 & n60517) | (n60516 & n60517);
  assign n60519 = n39632 | n60503;
  assign n60520 = n39229 | n39632;
  assign n60521 = (n72495 & n60519) | (n72495 & n60520) | (n60519 & n60520);
  assign n39635 = ~n60518 & n60521;
  assign n39636 = x173 & x192;
  assign n39637 = n39635 & n39636;
  assign n39638 = n39635 | n39636;
  assign n39639 = ~n39637 & n39638;
  assign n60522 = n39236 & n39639;
  assign n72589 = (n39639 & n60300) | (n39639 & n60522) | (n60300 & n60522);
  assign n72590 = (n39639 & n60299) | (n39639 & n60522) | (n60299 & n60522);
  assign n72591 = (n60050 & n72589) | (n60050 & n72590) | (n72589 & n72590);
  assign n60524 = n39236 | n39639;
  assign n72592 = n60300 | n60524;
  assign n72593 = n60299 | n60524;
  assign n72594 = (n60050 & n72592) | (n60050 & n72593) | (n72592 & n72593);
  assign n39642 = ~n72591 & n72594;
  assign n39643 = x172 & x193;
  assign n39644 = n39642 & n39643;
  assign n39645 = n39642 | n39643;
  assign n39646 = ~n39644 & n39645;
  assign n60501 = n39243 | n39245;
  assign n72595 = n39646 & n60501;
  assign n72566 = n38834 | n39243;
  assign n72567 = (n39243 & n39245) | (n39243 & n72566) | (n39245 & n72566);
  assign n72596 = n39646 & n72567;
  assign n72597 = (n60079 & n72595) | (n60079 & n72596) | (n72595 & n72596);
  assign n72598 = n39646 | n60501;
  assign n72599 = n39646 | n72567;
  assign n72600 = (n60079 & n72598) | (n60079 & n72599) | (n72598 & n72599);
  assign n39649 = ~n72597 & n72600;
  assign n39650 = x171 & x194;
  assign n39651 = n39649 & n39650;
  assign n39652 = n39649 | n39650;
  assign n39653 = ~n39651 & n39652;
  assign n60498 = n39250 | n39252;
  assign n60526 = n39653 & n60498;
  assign n60527 = n39250 & n39653;
  assign n60528 = (n72490 & n60526) | (n72490 & n60527) | (n60526 & n60527);
  assign n60529 = n39653 | n60498;
  assign n60530 = n39250 | n39653;
  assign n60531 = (n72490 & n60529) | (n72490 & n60530) | (n60529 & n60530);
  assign n39656 = ~n60528 & n60531;
  assign n39657 = x170 & x195;
  assign n39658 = n39656 & n39657;
  assign n39659 = n39656 | n39657;
  assign n39660 = ~n39658 & n39659;
  assign n60532 = n39257 & n39660;
  assign n72601 = (n39660 & n60310) | (n39660 & n60532) | (n60310 & n60532);
  assign n72602 = (n39660 & n60309) | (n39660 & n60532) | (n60309 & n60532);
  assign n72603 = (n60045 & n72601) | (n60045 & n72602) | (n72601 & n72602);
  assign n60534 = n39257 | n39660;
  assign n72604 = n60310 | n60534;
  assign n72605 = n60309 | n60534;
  assign n72606 = (n60045 & n72604) | (n60045 & n72605) | (n72604 & n72605);
  assign n39663 = ~n72603 & n72606;
  assign n39664 = x169 & x196;
  assign n39665 = n39663 & n39664;
  assign n39666 = n39663 | n39664;
  assign n39667 = ~n39665 & n39666;
  assign n60496 = n39264 | n39266;
  assign n72607 = n39667 & n60496;
  assign n72564 = n38855 | n39264;
  assign n72565 = (n39264 & n39266) | (n39264 & n72564) | (n39266 & n72564);
  assign n72608 = n39667 & n72565;
  assign n72609 = (n60089 & n72607) | (n60089 & n72608) | (n72607 & n72608);
  assign n72610 = n39667 | n60496;
  assign n72611 = n39667 | n72565;
  assign n72612 = (n60089 & n72610) | (n60089 & n72611) | (n72610 & n72611);
  assign n39670 = ~n72609 & n72612;
  assign n39671 = x168 & x197;
  assign n39672 = n39670 & n39671;
  assign n39673 = n39670 | n39671;
  assign n39674 = ~n39672 & n39673;
  assign n60493 = n39271 | n39273;
  assign n60536 = n39674 & n60493;
  assign n60537 = n39271 & n39674;
  assign n60538 = (n72485 & n60536) | (n72485 & n60537) | (n60536 & n60537);
  assign n60539 = n39674 | n60493;
  assign n60540 = n39271 | n39674;
  assign n60541 = (n72485 & n60539) | (n72485 & n60540) | (n60539 & n60540);
  assign n39677 = ~n60538 & n60541;
  assign n39678 = x167 & x198;
  assign n39679 = n39677 & n39678;
  assign n39680 = n39677 | n39678;
  assign n39681 = ~n39679 & n39680;
  assign n60542 = n39278 & n39681;
  assign n72613 = (n39681 & n60320) | (n39681 & n60542) | (n60320 & n60542);
  assign n72614 = (n39681 & n60319) | (n39681 & n60542) | (n60319 & n60542);
  assign n72615 = (n60040 & n72613) | (n60040 & n72614) | (n72613 & n72614);
  assign n60544 = n39278 | n39681;
  assign n72616 = n60320 | n60544;
  assign n72617 = n60319 | n60544;
  assign n72618 = (n60040 & n72616) | (n60040 & n72617) | (n72616 & n72617);
  assign n39684 = ~n72615 & n72618;
  assign n39685 = x166 & x199;
  assign n39686 = n39684 & n39685;
  assign n39687 = n39684 | n39685;
  assign n39688 = ~n39686 & n39687;
  assign n60491 = n39285 | n39287;
  assign n72619 = n39688 & n60491;
  assign n72562 = n38876 | n39285;
  assign n72563 = (n39285 & n39287) | (n39285 & n72562) | (n39287 & n72562);
  assign n72620 = n39688 & n72563;
  assign n72621 = (n60099 & n72619) | (n60099 & n72620) | (n72619 & n72620);
  assign n72622 = n39688 | n60491;
  assign n72623 = n39688 | n72563;
  assign n72624 = (n60099 & n72622) | (n60099 & n72623) | (n72622 & n72623);
  assign n39691 = ~n72621 & n72624;
  assign n39692 = x165 & x200;
  assign n39693 = n39691 & n39692;
  assign n39694 = n39691 | n39692;
  assign n39695 = ~n39693 & n39694;
  assign n60488 = n39292 | n39294;
  assign n60546 = n39695 & n60488;
  assign n60547 = n39292 & n39695;
  assign n60548 = (n72480 & n60546) | (n72480 & n60547) | (n60546 & n60547);
  assign n60549 = n39695 | n60488;
  assign n60550 = n39292 | n39695;
  assign n60551 = (n72480 & n60549) | (n72480 & n60550) | (n60549 & n60550);
  assign n39698 = ~n60548 & n60551;
  assign n39699 = x164 & x201;
  assign n39700 = n39698 & n39699;
  assign n39701 = n39698 | n39699;
  assign n39702 = ~n39700 & n39701;
  assign n60552 = n39299 & n39702;
  assign n72625 = (n39702 & n60330) | (n39702 & n60552) | (n60330 & n60552);
  assign n72626 = (n39702 & n60329) | (n39702 & n60552) | (n60329 & n60552);
  assign n72627 = (n60035 & n72625) | (n60035 & n72626) | (n72625 & n72626);
  assign n60554 = n39299 | n39702;
  assign n72628 = n60330 | n60554;
  assign n72629 = n60329 | n60554;
  assign n72630 = (n60035 & n72628) | (n60035 & n72629) | (n72628 & n72629);
  assign n39705 = ~n72627 & n72630;
  assign n39706 = x163 & x202;
  assign n39707 = n39705 & n39706;
  assign n39708 = n39705 | n39706;
  assign n39709 = ~n39707 & n39708;
  assign n60486 = n39306 | n39308;
  assign n72631 = n39709 & n60486;
  assign n72560 = n38897 | n39306;
  assign n72561 = (n39306 & n39308) | (n39306 & n72560) | (n39308 & n72560);
  assign n72632 = n39709 & n72561;
  assign n72633 = (n60109 & n72631) | (n60109 & n72632) | (n72631 & n72632);
  assign n72634 = n39709 | n60486;
  assign n72635 = n39709 | n72561;
  assign n72636 = (n60109 & n72634) | (n60109 & n72635) | (n72634 & n72635);
  assign n39712 = ~n72633 & n72636;
  assign n39713 = x162 & x203;
  assign n39714 = n39712 & n39713;
  assign n39715 = n39712 | n39713;
  assign n39716 = ~n39714 & n39715;
  assign n60483 = n39313 | n39315;
  assign n60556 = n39716 & n60483;
  assign n60557 = n39313 & n39716;
  assign n60558 = (n72475 & n60556) | (n72475 & n60557) | (n60556 & n60557);
  assign n60559 = n39716 | n60483;
  assign n60560 = n39313 | n39716;
  assign n60561 = (n72475 & n60559) | (n72475 & n60560) | (n60559 & n60560);
  assign n39719 = ~n60558 & n60561;
  assign n39720 = x161 & x204;
  assign n39721 = n39719 & n39720;
  assign n39722 = n39719 | n39720;
  assign n39723 = ~n39721 & n39722;
  assign n60562 = n39320 & n39723;
  assign n72637 = (n39723 & n60340) | (n39723 & n60562) | (n60340 & n60562);
  assign n72638 = (n39723 & n60339) | (n39723 & n60562) | (n60339 & n60562);
  assign n72639 = (n72354 & n72637) | (n72354 & n72638) | (n72637 & n72638);
  assign n60564 = n39320 | n39723;
  assign n72640 = n60340 | n60564;
  assign n72641 = n60339 | n60564;
  assign n72642 = (n72354 & n72640) | (n72354 & n72641) | (n72640 & n72641);
  assign n39726 = ~n72639 & n72642;
  assign n39727 = x160 & x205;
  assign n39728 = n39726 & n39727;
  assign n39729 = n39726 | n39727;
  assign n39730 = ~n39728 & n39729;
  assign n39731 = n72559 & n39730;
  assign n39732 = n72559 | n39730;
  assign n39733 = ~n39731 & n39732;
  assign n39734 = x159 & x206;
  assign n39735 = n39733 & n39734;
  assign n39736 = n39733 | n39734;
  assign n39737 = ~n39735 & n39736;
  assign n60478 = n39334 | n39336;
  assign n60566 = n39737 & n60478;
  assign n60567 = n39334 & n39737;
  assign n60568 = (n72470 & n60566) | (n72470 & n60567) | (n60566 & n60567);
  assign n60569 = n39737 | n60478;
  assign n60570 = n39334 | n39737;
  assign n60571 = (n72470 & n60569) | (n72470 & n60570) | (n60569 & n60570);
  assign n39740 = ~n60568 & n60571;
  assign n39741 = x158 & x207;
  assign n39742 = n39740 & n39741;
  assign n39743 = n39740 | n39741;
  assign n39744 = ~n39742 & n39743;
  assign n60572 = n39341 & n39744;
  assign n72643 = (n39744 & n60350) | (n39744 & n60572) | (n60350 & n60572);
  assign n72644 = (n39744 & n60349) | (n39744 & n60572) | (n60349 & n60572);
  assign n72645 = (n72349 & n72643) | (n72349 & n72644) | (n72643 & n72644);
  assign n60574 = n39341 | n39744;
  assign n72646 = n60350 | n60574;
  assign n72647 = n60349 | n60574;
  assign n72648 = (n72349 & n72646) | (n72349 & n72647) | (n72646 & n72647);
  assign n39747 = ~n72645 & n72648;
  assign n39748 = x157 & x208;
  assign n39749 = n39747 & n39748;
  assign n39750 = n39747 | n39748;
  assign n39751 = ~n39749 & n39750;
  assign n39752 = n72554 & n39751;
  assign n39753 = n72554 | n39751;
  assign n39754 = ~n39752 & n39753;
  assign n39755 = x156 & x209;
  assign n39756 = n39754 & n39755;
  assign n39757 = n39754 | n39755;
  assign n39758 = ~n39756 & n39757;
  assign n60473 = n39355 | n39357;
  assign n60576 = n39758 & n60473;
  assign n60577 = n39355 & n39758;
  assign n60578 = (n60249 & n60576) | (n60249 & n60577) | (n60576 & n60577);
  assign n60579 = n39758 | n60473;
  assign n60580 = n39355 | n39758;
  assign n60581 = (n60249 & n60579) | (n60249 & n60580) | (n60579 & n60580);
  assign n39761 = ~n60578 & n60581;
  assign n39762 = x155 & x210;
  assign n39763 = n39761 & n39762;
  assign n39764 = n39761 | n39762;
  assign n39765 = ~n39763 & n39764;
  assign n60582 = n39362 & n39765;
  assign n60583 = (n39765 & n72534) | (n39765 & n60582) | (n72534 & n60582);
  assign n60584 = n39362 | n39765;
  assign n60585 = n72534 | n60584;
  assign n39768 = ~n60583 & n60585;
  assign n39769 = x154 & x211;
  assign n39770 = n39768 & n39769;
  assign n39771 = n39768 | n39769;
  assign n39772 = ~n39770 & n39771;
  assign n60586 = n39369 & n39772;
  assign n60587 = (n39772 & n60364) | (n39772 & n60586) | (n60364 & n60586);
  assign n60588 = n39369 | n39772;
  assign n60589 = n60364 | n60588;
  assign n39775 = ~n60587 & n60589;
  assign n39776 = x153 & x212;
  assign n39777 = n39775 & n39776;
  assign n39778 = n39775 | n39776;
  assign n39779 = ~n39777 & n39778;
  assign n60590 = n39376 & n39779;
  assign n60591 = (n39779 & n60368) | (n39779 & n60590) | (n60368 & n60590);
  assign n60592 = n39376 | n39779;
  assign n60593 = n60368 | n60592;
  assign n39782 = ~n60591 & n60593;
  assign n39783 = x152 & x213;
  assign n39784 = n39782 & n39783;
  assign n39785 = n39782 | n39783;
  assign n39786 = ~n39784 & n39785;
  assign n60594 = n39383 & n39786;
  assign n60595 = (n39786 & n60372) | (n39786 & n60594) | (n60372 & n60594);
  assign n60596 = n39383 | n39786;
  assign n60597 = n60372 | n60596;
  assign n39789 = ~n60595 & n60597;
  assign n39790 = x151 & x214;
  assign n39791 = n39789 & n39790;
  assign n39792 = n39789 | n39790;
  assign n39793 = ~n39791 & n39792;
  assign n60598 = n39390 & n39793;
  assign n60599 = (n39793 & n60376) | (n39793 & n60598) | (n60376 & n60598);
  assign n60600 = n39390 | n39793;
  assign n60601 = n60376 | n60600;
  assign n39796 = ~n60599 & n60601;
  assign n39797 = x150 & x215;
  assign n39798 = n39796 & n39797;
  assign n39799 = n39796 | n39797;
  assign n39800 = ~n39798 & n39799;
  assign n60602 = n39397 & n39800;
  assign n60603 = (n39800 & n60380) | (n39800 & n60602) | (n60380 & n60602);
  assign n60604 = n39397 | n39800;
  assign n60605 = n60380 | n60604;
  assign n39803 = ~n60603 & n60605;
  assign n39804 = x149 & x216;
  assign n39805 = n39803 & n39804;
  assign n39806 = n39803 | n39804;
  assign n39807 = ~n39805 & n39806;
  assign n60606 = n39404 & n39807;
  assign n60607 = (n39807 & n60384) | (n39807 & n60606) | (n60384 & n60606);
  assign n60608 = n39404 | n39807;
  assign n60609 = n60384 | n60608;
  assign n39810 = ~n60607 & n60609;
  assign n39811 = x148 & x217;
  assign n39812 = n39810 & n39811;
  assign n39813 = n39810 | n39811;
  assign n39814 = ~n39812 & n39813;
  assign n60610 = n39411 & n39814;
  assign n60611 = (n39814 & n60388) | (n39814 & n60610) | (n60388 & n60610);
  assign n60612 = n39411 | n39814;
  assign n60613 = n60388 | n60612;
  assign n39817 = ~n60611 & n60613;
  assign n39818 = x147 & x218;
  assign n39819 = n39817 & n39818;
  assign n39820 = n39817 | n39818;
  assign n39821 = ~n39819 & n39820;
  assign n60614 = n39418 & n39821;
  assign n60615 = (n39821 & n60392) | (n39821 & n60614) | (n60392 & n60614);
  assign n60616 = n39418 | n39821;
  assign n60617 = n60392 | n60616;
  assign n39824 = ~n60615 & n60617;
  assign n39825 = x146 & x219;
  assign n39826 = n39824 & n39825;
  assign n39827 = n39824 | n39825;
  assign n39828 = ~n39826 & n39827;
  assign n60618 = n39425 & n39828;
  assign n60619 = (n39828 & n60396) | (n39828 & n60618) | (n60396 & n60618);
  assign n60620 = n39425 | n39828;
  assign n60621 = n60396 | n60620;
  assign n39831 = ~n60619 & n60621;
  assign n39832 = x145 & x220;
  assign n39833 = n39831 & n39832;
  assign n39834 = n39831 | n39832;
  assign n39835 = ~n39833 & n39834;
  assign n60622 = n39432 & n39835;
  assign n60623 = (n39835 & n60400) | (n39835 & n60622) | (n60400 & n60622);
  assign n60624 = n39432 | n39835;
  assign n60625 = n60400 | n60624;
  assign n39838 = ~n60623 & n60625;
  assign n39839 = x144 & x221;
  assign n39840 = n39838 & n39839;
  assign n39841 = n39838 | n39839;
  assign n39842 = ~n39840 & n39841;
  assign n60626 = n39439 & n39842;
  assign n60627 = (n39842 & n60404) | (n39842 & n60626) | (n60404 & n60626);
  assign n60628 = n39439 | n39842;
  assign n60629 = n60404 | n60628;
  assign n39845 = ~n60627 & n60629;
  assign n39846 = x143 & x222;
  assign n39847 = n39845 & n39846;
  assign n39848 = n39845 | n39846;
  assign n39849 = ~n39847 & n39848;
  assign n60630 = n39446 & n39849;
  assign n60631 = (n39849 & n60408) | (n39849 & n60630) | (n60408 & n60630);
  assign n60632 = n39446 | n39849;
  assign n60633 = n60408 | n60632;
  assign n39852 = ~n60631 & n60633;
  assign n39853 = x142 & x223;
  assign n39854 = n39852 & n39853;
  assign n39855 = n39852 | n39853;
  assign n39856 = ~n39854 & n39855;
  assign n60634 = n39453 & n39856;
  assign n60635 = (n39856 & n60412) | (n39856 & n60634) | (n60412 & n60634);
  assign n60636 = n39453 | n39856;
  assign n60637 = n60412 | n60636;
  assign n39859 = ~n60635 & n60637;
  assign n39860 = x141 & x224;
  assign n39861 = n39859 & n39860;
  assign n39862 = n39859 | n39860;
  assign n39863 = ~n39861 & n39862;
  assign n60638 = n39460 & n39863;
  assign n60639 = (n39863 & n60416) | (n39863 & n60638) | (n60416 & n60638);
  assign n60640 = n39460 | n39863;
  assign n60641 = n60416 | n60640;
  assign n39866 = ~n60639 & n60641;
  assign n39867 = x140 & x225;
  assign n39868 = n39866 & n39867;
  assign n39869 = n39866 | n39867;
  assign n39870 = ~n39868 & n39869;
  assign n60642 = n39467 & n39870;
  assign n60643 = (n39870 & n60420) | (n39870 & n60642) | (n60420 & n60642);
  assign n60644 = n39467 | n39870;
  assign n60645 = n60420 | n60644;
  assign n39873 = ~n60643 & n60645;
  assign n39874 = x139 & x226;
  assign n39875 = n39873 & n39874;
  assign n39876 = n39873 | n39874;
  assign n39877 = ~n39875 & n39876;
  assign n60646 = n39474 & n39877;
  assign n60647 = (n39877 & n60424) | (n39877 & n60646) | (n60424 & n60646);
  assign n60648 = n39474 | n39877;
  assign n60649 = n60424 | n60648;
  assign n39880 = ~n60647 & n60649;
  assign n39881 = x138 & x227;
  assign n39882 = n39880 & n39881;
  assign n39883 = n39880 | n39881;
  assign n39884 = ~n39882 & n39883;
  assign n60650 = n39481 & n39884;
  assign n60651 = (n39884 & n60428) | (n39884 & n60650) | (n60428 & n60650);
  assign n60652 = n39481 | n39884;
  assign n60653 = n60428 | n60652;
  assign n39887 = ~n60651 & n60653;
  assign n39888 = x137 & x228;
  assign n39889 = n39887 & n39888;
  assign n39890 = n39887 | n39888;
  assign n39891 = ~n39889 & n39890;
  assign n60654 = n39488 & n39891;
  assign n60655 = (n39891 & n60432) | (n39891 & n60654) | (n60432 & n60654);
  assign n60656 = n39488 | n39891;
  assign n60657 = n60432 | n60656;
  assign n39894 = ~n60655 & n60657;
  assign n39895 = x136 & x229;
  assign n39896 = n39894 & n39895;
  assign n39897 = n39894 | n39895;
  assign n39898 = ~n39896 & n39897;
  assign n60658 = n39495 & n39898;
  assign n60659 = (n39898 & n60436) | (n39898 & n60658) | (n60436 & n60658);
  assign n60660 = n39495 | n39898;
  assign n60661 = n60436 | n60660;
  assign n39901 = ~n60659 & n60661;
  assign n39902 = x135 & x230;
  assign n39903 = n39901 & n39902;
  assign n39904 = n39901 | n39902;
  assign n39905 = ~n39903 & n39904;
  assign n60662 = n39502 & n39905;
  assign n60663 = (n39905 & n60440) | (n39905 & n60662) | (n60440 & n60662);
  assign n60664 = n39502 | n39905;
  assign n60665 = n60440 | n60664;
  assign n39908 = ~n60663 & n60665;
  assign n39909 = x134 & x231;
  assign n39910 = n39908 & n39909;
  assign n39911 = n39908 | n39909;
  assign n39912 = ~n39910 & n39911;
  assign n60666 = n39509 & n39912;
  assign n60667 = (n39912 & n60444) | (n39912 & n60666) | (n60444 & n60666);
  assign n60668 = n39509 | n39912;
  assign n60669 = n60444 | n60668;
  assign n39915 = ~n60667 & n60669;
  assign n39916 = x133 & x232;
  assign n39917 = n39915 & n39916;
  assign n39918 = n39915 | n39916;
  assign n39919 = ~n39917 & n39918;
  assign n60670 = n39516 & n39919;
  assign n60671 = (n39919 & n60448) | (n39919 & n60670) | (n60448 & n60670);
  assign n60672 = n39516 | n39919;
  assign n60673 = n60448 | n60672;
  assign n39922 = ~n60671 & n60673;
  assign n39923 = x132 & x233;
  assign n39924 = n39922 & n39923;
  assign n39925 = n39922 | n39923;
  assign n39926 = ~n39924 & n39925;
  assign n60674 = n39523 & n39926;
  assign n60675 = (n39926 & n60452) | (n39926 & n60674) | (n60452 & n60674);
  assign n60676 = n39523 | n39926;
  assign n60677 = n60452 | n60676;
  assign n39929 = ~n60675 & n60677;
  assign n39930 = x131 & x234;
  assign n39931 = n39929 & n39930;
  assign n39932 = n39929 | n39930;
  assign n39933 = ~n39931 & n39932;
  assign n60678 = n39530 & n39933;
  assign n60679 = (n39933 & n60456) | (n39933 & n60678) | (n60456 & n60678);
  assign n60680 = n39530 | n39933;
  assign n60681 = n60456 | n60680;
  assign n39936 = ~n60679 & n60681;
  assign n39937 = x130 & x235;
  assign n39938 = n39936 & n39937;
  assign n39939 = n39936 | n39937;
  assign n39940 = ~n39938 & n39939;
  assign n60682 = n39537 & n39940;
  assign n60683 = (n39940 & n60461) | (n39940 & n60682) | (n60461 & n60682);
  assign n60684 = n39537 | n39940;
  assign n60685 = n60461 | n60684;
  assign n39943 = ~n60683 & n60685;
  assign n39944 = x129 & x236;
  assign n39945 = n39943 & n39944;
  assign n39946 = n39943 | n39944;
  assign n39947 = ~n39945 & n39946;
  assign n60471 = n39544 | n39546;
  assign n60686 = n39947 & n60471;
  assign n60687 = n39544 & n39947;
  assign n60688 = (n60244 & n60686) | (n60244 & n60687) | (n60686 & n60687);
  assign n60689 = n39947 | n60471;
  assign n60690 = n39544 | n39947;
  assign n60691 = (n60244 & n60689) | (n60244 & n60690) | (n60689 & n60690);
  assign n39950 = ~n60688 & n60691;
  assign n39951 = x128 & x237;
  assign n39952 = n39950 & n39951;
  assign n39953 = n39950 | n39951;
  assign n39954 = ~n39952 & n39953;
  assign n60469 = n39551 | n39553;
  assign n72649 = n39954 & n60469;
  assign n72650 = n39551 & n39954;
  assign n72651 = (n60242 & n72649) | (n60242 & n72650) | (n72649 & n72650);
  assign n72652 = n39954 | n60469;
  assign n72653 = n39551 | n39954;
  assign n72654 = (n60242 & n72652) | (n60242 & n72653) | (n72652 & n72653);
  assign n39957 = ~n72651 & n72654;
  assign n39958 = x127 & x238;
  assign n39959 = n39957 & n39958;
  assign n39960 = n39957 | n39958;
  assign n39961 = ~n39959 & n39960;
  assign n60467 = n39558 | n39560;
  assign n72655 = n39961 & n60467;
  assign n72656 = n39558 & n39961;
  assign n72657 = (n60240 & n72655) | (n60240 & n72656) | (n72655 & n72656);
  assign n72658 = n39961 | n60467;
  assign n72659 = n39558 | n39961;
  assign n72660 = (n60240 & n72658) | (n60240 & n72659) | (n72658 & n72659);
  assign n39964 = ~n72657 & n72660;
  assign n39965 = x126 & x239;
  assign n39966 = n39964 & n39965;
  assign n39967 = n39964 | n39965;
  assign n39968 = ~n39966 & n39967;
  assign n39969 = n60466 & n39968;
  assign n39970 = n60466 | n39968;
  assign n39971 = ~n39969 & n39970;
  assign n60468 = (n39558 & n60240) | (n39558 & n60467) | (n60240 & n60467);
  assign n60470 = (n39551 & n60242) | (n39551 & n60469) | (n60242 & n60469);
  assign n60704 = n39742 | n39744;
  assign n72663 = n39341 | n39742;
  assign n72664 = (n39742 & n39744) | (n39742 & n72663) | (n39744 & n72663);
  assign n72665 = (n60350 & n60704) | (n60350 & n72664) | (n60704 & n72664);
  assign n72666 = (n60349 & n60704) | (n60349 & n72664) | (n60704 & n72664);
  assign n72667 = (n72349 & n72665) | (n72349 & n72666) | (n72665 & n72666);
  assign n60709 = n39721 | n39723;
  assign n72668 = n39320 | n39721;
  assign n72669 = (n39721 & n39723) | (n39721 & n72668) | (n39723 & n72668);
  assign n72670 = (n60340 & n60709) | (n60340 & n72669) | (n60709 & n72669);
  assign n72671 = (n60339 & n60709) | (n60339 & n72669) | (n60709 & n72669);
  assign n72672 = (n72354 & n72670) | (n72354 & n72671) | (n72670 & n72671);
  assign n60487 = (n60109 & n72561) | (n60109 & n60486) | (n72561 & n60486);
  assign n60714 = n39700 | n39702;
  assign n72673 = n39299 | n39700;
  assign n72674 = (n39700 & n39702) | (n39700 & n72673) | (n39702 & n72673);
  assign n72675 = (n60330 & n60714) | (n60330 & n72674) | (n60714 & n72674);
  assign n72676 = (n60329 & n60714) | (n60329 & n72674) | (n60714 & n72674);
  assign n72677 = (n60035 & n72675) | (n60035 & n72676) | (n72675 & n72676);
  assign n60492 = (n60099 & n72563) | (n60099 & n60491) | (n72563 & n60491);
  assign n60719 = n39679 | n39681;
  assign n72678 = n39278 | n39679;
  assign n72679 = (n39679 & n39681) | (n39679 & n72678) | (n39681 & n72678);
  assign n72680 = (n60320 & n60719) | (n60320 & n72679) | (n60719 & n72679);
  assign n72681 = (n60319 & n60719) | (n60319 & n72679) | (n60719 & n72679);
  assign n72682 = (n60040 & n72680) | (n60040 & n72681) | (n72680 & n72681);
  assign n60497 = (n60089 & n72565) | (n60089 & n60496) | (n72565 & n60496);
  assign n60724 = n39658 | n39660;
  assign n72683 = n39257 | n39658;
  assign n72684 = (n39658 & n39660) | (n39658 & n72683) | (n39660 & n72683);
  assign n72685 = (n60310 & n60724) | (n60310 & n72684) | (n60724 & n72684);
  assign n72686 = (n60309 & n60724) | (n60309 & n72684) | (n60724 & n72684);
  assign n72687 = (n60045 & n72685) | (n60045 & n72686) | (n72685 & n72686);
  assign n60502 = (n60079 & n72567) | (n60079 & n60501) | (n72567 & n60501);
  assign n60729 = n39637 | n39639;
  assign n72688 = n39236 | n39637;
  assign n72689 = (n39637 & n39639) | (n39637 & n72688) | (n39639 & n72688);
  assign n72690 = (n60300 & n60729) | (n60300 & n72689) | (n60729 & n72689);
  assign n72691 = (n60299 & n60729) | (n60299 & n72689) | (n60729 & n72689);
  assign n72692 = (n60050 & n72690) | (n60050 & n72691) | (n72690 & n72691);
  assign n72693 = n39229 | n39630;
  assign n72694 = (n39630 & n39632) | (n39630 & n72693) | (n39632 & n72693);
  assign n60732 = n39630 | n60516;
  assign n60733 = (n72495 & n72694) | (n72495 & n60732) | (n72694 & n60732);
  assign n40022 = x175 & x191;
  assign n72695 = n40022 & n72581;
  assign n72696 = (n39625 & n40022) | (n39625 & n72695) | (n40022 & n72695);
  assign n60737 = n40022 & n72581;
  assign n60738 = (n72574 & n72696) | (n72574 & n60737) | (n72696 & n60737);
  assign n72697 = n40022 | n72581;
  assign n72698 = n39625 | n72697;
  assign n60740 = n40022 | n72581;
  assign n60741 = (n72574 & n72698) | (n72574 & n60740) | (n72698 & n60740);
  assign n40025 = ~n60738 & n60741;
  assign n40026 = n60733 & n40025;
  assign n40027 = n60733 | n40025;
  assign n40028 = ~n40026 & n40027;
  assign n40029 = x174 & x192;
  assign n40030 = n40028 & n40029;
  assign n40031 = n40028 | n40029;
  assign n40032 = ~n40030 & n40031;
  assign n40033 = n72692 & n40032;
  assign n40034 = n72692 | n40032;
  assign n40035 = ~n40033 & n40034;
  assign n40036 = x173 & x193;
  assign n40037 = n40035 & n40036;
  assign n40038 = n40035 | n40036;
  assign n40039 = ~n40037 & n40038;
  assign n60726 = n39644 | n39646;
  assign n60742 = n40039 & n60726;
  assign n60743 = n39644 & n40039;
  assign n60744 = (n60502 & n60742) | (n60502 & n60743) | (n60742 & n60743);
  assign n60745 = n40039 | n60726;
  assign n60746 = n39644 | n40039;
  assign n60747 = (n60502 & n60745) | (n60502 & n60746) | (n60745 & n60746);
  assign n40042 = ~n60744 & n60747;
  assign n40043 = x172 & x194;
  assign n40044 = n40042 & n40043;
  assign n40045 = n40042 | n40043;
  assign n40046 = ~n40044 & n40045;
  assign n60748 = n39651 & n40046;
  assign n60749 = (n40046 & n60528) | (n40046 & n60748) | (n60528 & n60748);
  assign n60750 = n39651 | n40046;
  assign n60751 = n60528 | n60750;
  assign n40049 = ~n60749 & n60751;
  assign n40050 = x171 & x195;
  assign n40051 = n40049 & n40050;
  assign n40052 = n40049 | n40050;
  assign n40053 = ~n40051 & n40052;
  assign n40054 = n72687 & n40053;
  assign n40055 = n72687 | n40053;
  assign n40056 = ~n40054 & n40055;
  assign n40057 = x170 & x196;
  assign n40058 = n40056 & n40057;
  assign n40059 = n40056 | n40057;
  assign n40060 = ~n40058 & n40059;
  assign n60721 = n39665 | n39667;
  assign n60752 = n40060 & n60721;
  assign n60753 = n39665 & n40060;
  assign n60754 = (n60497 & n60752) | (n60497 & n60753) | (n60752 & n60753);
  assign n60755 = n40060 | n60721;
  assign n60756 = n39665 | n40060;
  assign n60757 = (n60497 & n60755) | (n60497 & n60756) | (n60755 & n60756);
  assign n40063 = ~n60754 & n60757;
  assign n40064 = x169 & x197;
  assign n40065 = n40063 & n40064;
  assign n40066 = n40063 | n40064;
  assign n40067 = ~n40065 & n40066;
  assign n60758 = n39672 & n40067;
  assign n60759 = (n40067 & n60538) | (n40067 & n60758) | (n60538 & n60758);
  assign n60760 = n39672 | n40067;
  assign n60761 = n60538 | n60760;
  assign n40070 = ~n60759 & n60761;
  assign n40071 = x168 & x198;
  assign n40072 = n40070 & n40071;
  assign n40073 = n40070 | n40071;
  assign n40074 = ~n40072 & n40073;
  assign n40075 = n72682 & n40074;
  assign n40076 = n72682 | n40074;
  assign n40077 = ~n40075 & n40076;
  assign n40078 = x167 & x199;
  assign n40079 = n40077 & n40078;
  assign n40080 = n40077 | n40078;
  assign n40081 = ~n40079 & n40080;
  assign n60716 = n39686 | n39688;
  assign n60762 = n40081 & n60716;
  assign n60763 = n39686 & n40081;
  assign n60764 = (n60492 & n60762) | (n60492 & n60763) | (n60762 & n60763);
  assign n60765 = n40081 | n60716;
  assign n60766 = n39686 | n40081;
  assign n60767 = (n60492 & n60765) | (n60492 & n60766) | (n60765 & n60766);
  assign n40084 = ~n60764 & n60767;
  assign n40085 = x166 & x200;
  assign n40086 = n40084 & n40085;
  assign n40087 = n40084 | n40085;
  assign n40088 = ~n40086 & n40087;
  assign n60768 = n39693 & n40088;
  assign n60769 = (n40088 & n60548) | (n40088 & n60768) | (n60548 & n60768);
  assign n60770 = n39693 | n40088;
  assign n60771 = n60548 | n60770;
  assign n40091 = ~n60769 & n60771;
  assign n40092 = x165 & x201;
  assign n40093 = n40091 & n40092;
  assign n40094 = n40091 | n40092;
  assign n40095 = ~n40093 & n40094;
  assign n40096 = n72677 & n40095;
  assign n40097 = n72677 | n40095;
  assign n40098 = ~n40096 & n40097;
  assign n40099 = x164 & x202;
  assign n40100 = n40098 & n40099;
  assign n40101 = n40098 | n40099;
  assign n40102 = ~n40100 & n40101;
  assign n60711 = n39707 | n39709;
  assign n60772 = n40102 & n60711;
  assign n60773 = n39707 & n40102;
  assign n60774 = (n60487 & n60772) | (n60487 & n60773) | (n60772 & n60773);
  assign n60775 = n40102 | n60711;
  assign n60776 = n39707 | n40102;
  assign n60777 = (n60487 & n60775) | (n60487 & n60776) | (n60775 & n60776);
  assign n40105 = ~n60774 & n60777;
  assign n40106 = x163 & x203;
  assign n40107 = n40105 & n40106;
  assign n40108 = n40105 | n40106;
  assign n40109 = ~n40107 & n40108;
  assign n60778 = n39714 & n40109;
  assign n60779 = (n40109 & n60558) | (n40109 & n60778) | (n60558 & n60778);
  assign n60780 = n39714 | n40109;
  assign n60781 = n60558 | n60780;
  assign n40112 = ~n60779 & n60781;
  assign n40113 = x162 & x204;
  assign n40114 = n40112 & n40113;
  assign n40115 = n40112 | n40113;
  assign n40116 = ~n40114 & n40115;
  assign n40117 = n72672 & n40116;
  assign n40118 = n72672 | n40116;
  assign n40119 = ~n40117 & n40118;
  assign n40120 = x161 & x205;
  assign n40121 = n40119 & n40120;
  assign n40122 = n40119 | n40120;
  assign n40123 = ~n40121 & n40122;
  assign n60706 = n39728 | n39730;
  assign n60782 = n40123 & n60706;
  assign n60783 = n39728 & n40123;
  assign n60784 = (n72559 & n60782) | (n72559 & n60783) | (n60782 & n60783);
  assign n60785 = n40123 | n60706;
  assign n60786 = n39728 | n40123;
  assign n60787 = (n72559 & n60785) | (n72559 & n60786) | (n60785 & n60786);
  assign n40126 = ~n60784 & n60787;
  assign n40127 = x160 & x206;
  assign n40128 = n40126 & n40127;
  assign n40129 = n40126 | n40127;
  assign n40130 = ~n40128 & n40129;
  assign n60788 = n39735 & n40130;
  assign n72699 = (n40130 & n60567) | (n40130 & n60788) | (n60567 & n60788);
  assign n72700 = (n40130 & n60566) | (n40130 & n60788) | (n60566 & n60788);
  assign n72701 = (n72470 & n72699) | (n72470 & n72700) | (n72699 & n72700);
  assign n60790 = n39735 | n40130;
  assign n72702 = n60567 | n60790;
  assign n72703 = n60566 | n60790;
  assign n72704 = (n72470 & n72702) | (n72470 & n72703) | (n72702 & n72703);
  assign n40133 = ~n72701 & n72704;
  assign n40134 = x159 & x207;
  assign n40135 = n40133 & n40134;
  assign n40136 = n40133 | n40134;
  assign n40137 = ~n40135 & n40136;
  assign n40138 = n72667 & n40137;
  assign n40139 = n72667 | n40137;
  assign n40140 = ~n40138 & n40139;
  assign n40141 = x158 & x208;
  assign n40142 = n40140 & n40141;
  assign n40143 = n40140 | n40141;
  assign n40144 = ~n40142 & n40143;
  assign n60701 = n39749 | n39751;
  assign n60792 = n40144 & n60701;
  assign n60793 = n39749 & n40144;
  assign n60794 = (n72554 & n60792) | (n72554 & n60793) | (n60792 & n60793);
  assign n60795 = n40144 | n60701;
  assign n60796 = n39749 | n40144;
  assign n60797 = (n72554 & n60795) | (n72554 & n60796) | (n60795 & n60796);
  assign n40147 = ~n60794 & n60797;
  assign n40148 = x157 & x209;
  assign n40149 = n40147 & n40148;
  assign n40150 = n40147 | n40148;
  assign n40151 = ~n40149 & n40150;
  assign n60798 = n39756 & n40151;
  assign n72705 = (n40151 & n60577) | (n40151 & n60798) | (n60577 & n60798);
  assign n72706 = (n40151 & n60576) | (n40151 & n60798) | (n60576 & n60798);
  assign n72707 = (n60249 & n72705) | (n60249 & n72706) | (n72705 & n72706);
  assign n60800 = n39756 | n40151;
  assign n72708 = n60577 | n60800;
  assign n72709 = n60576 | n60800;
  assign n72710 = (n60249 & n72708) | (n60249 & n72709) | (n72708 & n72709);
  assign n40154 = ~n72707 & n72710;
  assign n40155 = x156 & x210;
  assign n40156 = n40154 & n40155;
  assign n40157 = n40154 | n40155;
  assign n40158 = ~n40156 & n40157;
  assign n60699 = n39763 | n39765;
  assign n72711 = n40158 & n60699;
  assign n72661 = n39362 | n39763;
  assign n72662 = (n39763 & n39765) | (n39763 & n72661) | (n39765 & n72661);
  assign n72712 = n40158 & n72662;
  assign n72713 = (n72534 & n72711) | (n72534 & n72712) | (n72711 & n72712);
  assign n72714 = n40158 | n60699;
  assign n72715 = n40158 | n72662;
  assign n72716 = (n72534 & n72714) | (n72534 & n72715) | (n72714 & n72715);
  assign n40161 = ~n72713 & n72716;
  assign n40162 = x155 & x211;
  assign n40163 = n40161 & n40162;
  assign n40164 = n40161 | n40162;
  assign n40165 = ~n40163 & n40164;
  assign n60802 = n39770 & n40165;
  assign n72717 = (n40165 & n60586) | (n40165 & n60802) | (n60586 & n60802);
  assign n72718 = (n39772 & n40165) | (n39772 & n60802) | (n40165 & n60802);
  assign n72719 = (n60364 & n72717) | (n60364 & n72718) | (n72717 & n72718);
  assign n60804 = n39770 | n40165;
  assign n72720 = n60586 | n60804;
  assign n72721 = n39772 | n60804;
  assign n72722 = (n60364 & n72720) | (n60364 & n72721) | (n72720 & n72721);
  assign n40168 = ~n72719 & n72722;
  assign n40169 = x154 & x212;
  assign n40170 = n40168 & n40169;
  assign n40171 = n40168 | n40169;
  assign n40172 = ~n40170 & n40171;
  assign n60806 = n39777 & n40172;
  assign n60807 = (n40172 & n60591) | (n40172 & n60806) | (n60591 & n60806);
  assign n60808 = n39777 | n40172;
  assign n60809 = n60591 | n60808;
  assign n40175 = ~n60807 & n60809;
  assign n40176 = x153 & x213;
  assign n40177 = n40175 & n40176;
  assign n40178 = n40175 | n40176;
  assign n40179 = ~n40177 & n40178;
  assign n60810 = n39784 & n40179;
  assign n60811 = (n40179 & n60595) | (n40179 & n60810) | (n60595 & n60810);
  assign n60812 = n39784 | n40179;
  assign n60813 = n60595 | n60812;
  assign n40182 = ~n60811 & n60813;
  assign n40183 = x152 & x214;
  assign n40184 = n40182 & n40183;
  assign n40185 = n40182 | n40183;
  assign n40186 = ~n40184 & n40185;
  assign n60814 = n39791 & n40186;
  assign n60815 = (n40186 & n60599) | (n40186 & n60814) | (n60599 & n60814);
  assign n60816 = n39791 | n40186;
  assign n60817 = n60599 | n60816;
  assign n40189 = ~n60815 & n60817;
  assign n40190 = x151 & x215;
  assign n40191 = n40189 & n40190;
  assign n40192 = n40189 | n40190;
  assign n40193 = ~n40191 & n40192;
  assign n60818 = n39798 & n40193;
  assign n60819 = (n40193 & n60603) | (n40193 & n60818) | (n60603 & n60818);
  assign n60820 = n39798 | n40193;
  assign n60821 = n60603 | n60820;
  assign n40196 = ~n60819 & n60821;
  assign n40197 = x150 & x216;
  assign n40198 = n40196 & n40197;
  assign n40199 = n40196 | n40197;
  assign n40200 = ~n40198 & n40199;
  assign n60822 = n39805 & n40200;
  assign n60823 = (n40200 & n60607) | (n40200 & n60822) | (n60607 & n60822);
  assign n60824 = n39805 | n40200;
  assign n60825 = n60607 | n60824;
  assign n40203 = ~n60823 & n60825;
  assign n40204 = x149 & x217;
  assign n40205 = n40203 & n40204;
  assign n40206 = n40203 | n40204;
  assign n40207 = ~n40205 & n40206;
  assign n60826 = n39812 & n40207;
  assign n60827 = (n40207 & n60611) | (n40207 & n60826) | (n60611 & n60826);
  assign n60828 = n39812 | n40207;
  assign n60829 = n60611 | n60828;
  assign n40210 = ~n60827 & n60829;
  assign n40211 = x148 & x218;
  assign n40212 = n40210 & n40211;
  assign n40213 = n40210 | n40211;
  assign n40214 = ~n40212 & n40213;
  assign n60830 = n39819 & n40214;
  assign n60831 = (n40214 & n60615) | (n40214 & n60830) | (n60615 & n60830);
  assign n60832 = n39819 | n40214;
  assign n60833 = n60615 | n60832;
  assign n40217 = ~n60831 & n60833;
  assign n40218 = x147 & x219;
  assign n40219 = n40217 & n40218;
  assign n40220 = n40217 | n40218;
  assign n40221 = ~n40219 & n40220;
  assign n60834 = n39826 & n40221;
  assign n60835 = (n40221 & n60619) | (n40221 & n60834) | (n60619 & n60834);
  assign n60836 = n39826 | n40221;
  assign n60837 = n60619 | n60836;
  assign n40224 = ~n60835 & n60837;
  assign n40225 = x146 & x220;
  assign n40226 = n40224 & n40225;
  assign n40227 = n40224 | n40225;
  assign n40228 = ~n40226 & n40227;
  assign n60838 = n39833 & n40228;
  assign n60839 = (n40228 & n60623) | (n40228 & n60838) | (n60623 & n60838);
  assign n60840 = n39833 | n40228;
  assign n60841 = n60623 | n60840;
  assign n40231 = ~n60839 & n60841;
  assign n40232 = x145 & x221;
  assign n40233 = n40231 & n40232;
  assign n40234 = n40231 | n40232;
  assign n40235 = ~n40233 & n40234;
  assign n60842 = n39840 & n40235;
  assign n60843 = (n40235 & n60627) | (n40235 & n60842) | (n60627 & n60842);
  assign n60844 = n39840 | n40235;
  assign n60845 = n60627 | n60844;
  assign n40238 = ~n60843 & n60845;
  assign n40239 = x144 & x222;
  assign n40240 = n40238 & n40239;
  assign n40241 = n40238 | n40239;
  assign n40242 = ~n40240 & n40241;
  assign n60846 = n39847 & n40242;
  assign n60847 = (n40242 & n60631) | (n40242 & n60846) | (n60631 & n60846);
  assign n60848 = n39847 | n40242;
  assign n60849 = n60631 | n60848;
  assign n40245 = ~n60847 & n60849;
  assign n40246 = x143 & x223;
  assign n40247 = n40245 & n40246;
  assign n40248 = n40245 | n40246;
  assign n40249 = ~n40247 & n40248;
  assign n60850 = n39854 & n40249;
  assign n60851 = (n40249 & n60635) | (n40249 & n60850) | (n60635 & n60850);
  assign n60852 = n39854 | n40249;
  assign n60853 = n60635 | n60852;
  assign n40252 = ~n60851 & n60853;
  assign n40253 = x142 & x224;
  assign n40254 = n40252 & n40253;
  assign n40255 = n40252 | n40253;
  assign n40256 = ~n40254 & n40255;
  assign n60854 = n39861 & n40256;
  assign n60855 = (n40256 & n60639) | (n40256 & n60854) | (n60639 & n60854);
  assign n60856 = n39861 | n40256;
  assign n60857 = n60639 | n60856;
  assign n40259 = ~n60855 & n60857;
  assign n40260 = x141 & x225;
  assign n40261 = n40259 & n40260;
  assign n40262 = n40259 | n40260;
  assign n40263 = ~n40261 & n40262;
  assign n60858 = n39868 & n40263;
  assign n60859 = (n40263 & n60643) | (n40263 & n60858) | (n60643 & n60858);
  assign n60860 = n39868 | n40263;
  assign n60861 = n60643 | n60860;
  assign n40266 = ~n60859 & n60861;
  assign n40267 = x140 & x226;
  assign n40268 = n40266 & n40267;
  assign n40269 = n40266 | n40267;
  assign n40270 = ~n40268 & n40269;
  assign n60862 = n39875 & n40270;
  assign n60863 = (n40270 & n60647) | (n40270 & n60862) | (n60647 & n60862);
  assign n60864 = n39875 | n40270;
  assign n60865 = n60647 | n60864;
  assign n40273 = ~n60863 & n60865;
  assign n40274 = x139 & x227;
  assign n40275 = n40273 & n40274;
  assign n40276 = n40273 | n40274;
  assign n40277 = ~n40275 & n40276;
  assign n60866 = n39882 & n40277;
  assign n60867 = (n40277 & n60651) | (n40277 & n60866) | (n60651 & n60866);
  assign n60868 = n39882 | n40277;
  assign n60869 = n60651 | n60868;
  assign n40280 = ~n60867 & n60869;
  assign n40281 = x138 & x228;
  assign n40282 = n40280 & n40281;
  assign n40283 = n40280 | n40281;
  assign n40284 = ~n40282 & n40283;
  assign n60870 = n39889 & n40284;
  assign n60871 = (n40284 & n60655) | (n40284 & n60870) | (n60655 & n60870);
  assign n60872 = n39889 | n40284;
  assign n60873 = n60655 | n60872;
  assign n40287 = ~n60871 & n60873;
  assign n40288 = x137 & x229;
  assign n40289 = n40287 & n40288;
  assign n40290 = n40287 | n40288;
  assign n40291 = ~n40289 & n40290;
  assign n60874 = n39896 & n40291;
  assign n60875 = (n40291 & n60659) | (n40291 & n60874) | (n60659 & n60874);
  assign n60876 = n39896 | n40291;
  assign n60877 = n60659 | n60876;
  assign n40294 = ~n60875 & n60877;
  assign n40295 = x136 & x230;
  assign n40296 = n40294 & n40295;
  assign n40297 = n40294 | n40295;
  assign n40298 = ~n40296 & n40297;
  assign n60878 = n39903 & n40298;
  assign n60879 = (n40298 & n60663) | (n40298 & n60878) | (n60663 & n60878);
  assign n60880 = n39903 | n40298;
  assign n60881 = n60663 | n60880;
  assign n40301 = ~n60879 & n60881;
  assign n40302 = x135 & x231;
  assign n40303 = n40301 & n40302;
  assign n40304 = n40301 | n40302;
  assign n40305 = ~n40303 & n40304;
  assign n60882 = n39910 & n40305;
  assign n60883 = (n40305 & n60667) | (n40305 & n60882) | (n60667 & n60882);
  assign n60884 = n39910 | n40305;
  assign n60885 = n60667 | n60884;
  assign n40308 = ~n60883 & n60885;
  assign n40309 = x134 & x232;
  assign n40310 = n40308 & n40309;
  assign n40311 = n40308 | n40309;
  assign n40312 = ~n40310 & n40311;
  assign n60886 = n39917 & n40312;
  assign n60887 = (n40312 & n60671) | (n40312 & n60886) | (n60671 & n60886);
  assign n60888 = n39917 | n40312;
  assign n60889 = n60671 | n60888;
  assign n40315 = ~n60887 & n60889;
  assign n40316 = x133 & x233;
  assign n40317 = n40315 & n40316;
  assign n40318 = n40315 | n40316;
  assign n40319 = ~n40317 & n40318;
  assign n60890 = n39924 & n40319;
  assign n60891 = (n40319 & n60675) | (n40319 & n60890) | (n60675 & n60890);
  assign n60892 = n39924 | n40319;
  assign n60893 = n60675 | n60892;
  assign n40322 = ~n60891 & n60893;
  assign n40323 = x132 & x234;
  assign n40324 = n40322 & n40323;
  assign n40325 = n40322 | n40323;
  assign n40326 = ~n40324 & n40325;
  assign n60894 = n39931 & n40326;
  assign n60895 = (n40326 & n60679) | (n40326 & n60894) | (n60679 & n60894);
  assign n60896 = n39931 | n40326;
  assign n60897 = n60679 | n60896;
  assign n40329 = ~n60895 & n60897;
  assign n40330 = x131 & x235;
  assign n40331 = n40329 & n40330;
  assign n40332 = n40329 | n40330;
  assign n40333 = ~n40331 & n40332;
  assign n60898 = n39938 & n40333;
  assign n60899 = (n40333 & n60683) | (n40333 & n60898) | (n60683 & n60898);
  assign n60900 = n39938 | n40333;
  assign n60901 = n60683 | n60900;
  assign n40336 = ~n60899 & n60901;
  assign n40337 = x130 & x236;
  assign n40338 = n40336 & n40337;
  assign n40339 = n40336 | n40337;
  assign n40340 = ~n40338 & n40339;
  assign n60902 = n39945 & n40340;
  assign n60903 = (n40340 & n60688) | (n40340 & n60902) | (n60688 & n60902);
  assign n60904 = n39945 | n40340;
  assign n60905 = n60688 | n60904;
  assign n40343 = ~n60903 & n60905;
  assign n40344 = x129 & x237;
  assign n40345 = n40343 & n40344;
  assign n40346 = n40343 | n40344;
  assign n40347 = ~n40345 & n40346;
  assign n60696 = n39952 | n39954;
  assign n60906 = n40347 & n60696;
  assign n60907 = n39952 & n40347;
  assign n60908 = (n60470 & n60906) | (n60470 & n60907) | (n60906 & n60907);
  assign n60909 = n40347 | n60696;
  assign n60910 = n39952 | n40347;
  assign n60911 = (n60470 & n60909) | (n60470 & n60910) | (n60909 & n60910);
  assign n40350 = ~n60908 & n60911;
  assign n40351 = x128 & x238;
  assign n40352 = n40350 & n40351;
  assign n40353 = n40350 | n40351;
  assign n40354 = ~n40352 & n40353;
  assign n60694 = n39959 | n39961;
  assign n72723 = n40354 & n60694;
  assign n72724 = n39959 & n40354;
  assign n72725 = (n60468 & n72723) | (n60468 & n72724) | (n72723 & n72724);
  assign n72726 = n40354 | n60694;
  assign n72727 = n39959 | n40354;
  assign n72728 = (n60468 & n72726) | (n60468 & n72727) | (n72726 & n72727);
  assign n40357 = ~n72725 & n72728;
  assign n40358 = x127 & x239;
  assign n40359 = n40357 & n40358;
  assign n40360 = n40357 | n40358;
  assign n40361 = ~n40359 & n40360;
  assign n60692 = n39966 | n39968;
  assign n72729 = n40361 & n60692;
  assign n72730 = n39966 & n40361;
  assign n72731 = (n60466 & n72729) | (n60466 & n72730) | (n72729 & n72730);
  assign n72732 = n40361 | n60692;
  assign n72733 = n39966 | n40361;
  assign n72734 = (n60466 & n72732) | (n60466 & n72733) | (n72732 & n72733);
  assign n40364 = ~n72731 & n72734;
  assign n60693 = (n39966 & n60466) | (n39966 & n60692) | (n60466 & n60692);
  assign n60695 = (n39959 & n60468) | (n39959 & n60694) | (n60468 & n60694);
  assign n60700 = (n72534 & n72662) | (n72534 & n60699) | (n72662 & n60699);
  assign n60919 = n40149 | n40151;
  assign n72735 = n39756 | n40149;
  assign n72736 = (n40149 & n40151) | (n40149 & n72735) | (n40151 & n72735);
  assign n72737 = (n60577 & n60919) | (n60577 & n72736) | (n60919 & n72736);
  assign n72738 = (n60576 & n60919) | (n60576 & n72736) | (n60919 & n72736);
  assign n72739 = (n60249 & n72737) | (n60249 & n72738) | (n72737 & n72738);
  assign n60924 = n40128 | n40130;
  assign n72740 = n39735 | n40128;
  assign n72741 = (n40128 & n40130) | (n40128 & n72740) | (n40130 & n72740);
  assign n72742 = (n60567 & n60924) | (n60567 & n72741) | (n60924 & n72741);
  assign n72743 = (n60566 & n60924) | (n60566 & n72741) | (n60924 & n72741);
  assign n72744 = (n72470 & n72742) | (n72470 & n72743) | (n72742 & n72743);
  assign n40414 = x175 & x192;
  assign n72754 = n40414 & n72696;
  assign n72755 = n40414 & n60737;
  assign n72756 = (n72574 & n72754) | (n72574 & n72755) | (n72754 & n72755);
  assign n72753 = (n40025 & n40414) | (n40025 & n72756) | (n40414 & n72756);
  assign n60952 = (n60733 & n72753) | (n60733 & n72756) | (n72753 & n72756);
  assign n72758 = n40414 | n72696;
  assign n72759 = n40414 | n60737;
  assign n72760 = (n72574 & n72758) | (n72574 & n72759) | (n72758 & n72759);
  assign n72757 = n40025 | n72760;
  assign n60955 = (n60733 & n72757) | (n60733 & n72760) | (n72757 & n72760);
  assign n40417 = ~n60952 & n60955;
  assign n60957 = n40030 & n40417;
  assign n72761 = (n40032 & n40417) | (n40032 & n60957) | (n40417 & n60957);
  assign n60958 = (n72692 & n72761) | (n72692 & n60957) | (n72761 & n60957);
  assign n60960 = n40030 | n40417;
  assign n72762 = n40032 | n60960;
  assign n60961 = (n72692 & n72762) | (n72692 & n60960) | (n72762 & n60960);
  assign n40420 = ~n60958 & n60961;
  assign n40421 = x174 & x193;
  assign n40422 = n40420 & n40421;
  assign n40423 = n40420 | n40421;
  assign n40424 = ~n40422 & n40423;
  assign n60962 = n40037 & n40424;
  assign n72763 = (n40424 & n60743) | (n40424 & n60962) | (n60743 & n60962);
  assign n72764 = (n40424 & n60742) | (n40424 & n60962) | (n60742 & n60962);
  assign n72765 = (n60502 & n72763) | (n60502 & n72764) | (n72763 & n72764);
  assign n60964 = n40037 | n40424;
  assign n72766 = n60743 | n60964;
  assign n72767 = n60742 | n60964;
  assign n72768 = (n60502 & n72766) | (n60502 & n72767) | (n72766 & n72767);
  assign n40427 = ~n72765 & n72768;
  assign n40428 = x173 & x194;
  assign n40429 = n40427 & n40428;
  assign n40430 = n40427 | n40428;
  assign n40431 = ~n40429 & n40430;
  assign n60944 = n40044 | n40046;
  assign n72769 = n40431 & n60944;
  assign n72751 = n39651 | n40044;
  assign n72752 = (n40044 & n40046) | (n40044 & n72751) | (n40046 & n72751);
  assign n72770 = n40431 & n72752;
  assign n72771 = (n60528 & n72769) | (n60528 & n72770) | (n72769 & n72770);
  assign n72772 = n40431 | n60944;
  assign n72773 = n40431 | n72752;
  assign n72774 = (n60528 & n72772) | (n60528 & n72773) | (n72772 & n72773);
  assign n40434 = ~n72771 & n72774;
  assign n40435 = x172 & x195;
  assign n40436 = n40434 & n40435;
  assign n40437 = n40434 | n40435;
  assign n40438 = ~n40436 & n40437;
  assign n60941 = n40051 | n40053;
  assign n60966 = n40438 & n60941;
  assign n60967 = n40051 & n40438;
  assign n60968 = (n72687 & n60966) | (n72687 & n60967) | (n60966 & n60967);
  assign n60969 = n40438 | n60941;
  assign n60970 = n40051 | n40438;
  assign n60971 = (n72687 & n60969) | (n72687 & n60970) | (n60969 & n60970);
  assign n40441 = ~n60968 & n60971;
  assign n40442 = x171 & x196;
  assign n40443 = n40441 & n40442;
  assign n40444 = n40441 | n40442;
  assign n40445 = ~n40443 & n40444;
  assign n60972 = n40058 & n40445;
  assign n72775 = (n40445 & n60753) | (n40445 & n60972) | (n60753 & n60972);
  assign n72776 = (n40445 & n60752) | (n40445 & n60972) | (n60752 & n60972);
  assign n72777 = (n60497 & n72775) | (n60497 & n72776) | (n72775 & n72776);
  assign n60974 = n40058 | n40445;
  assign n72778 = n60753 | n60974;
  assign n72779 = n60752 | n60974;
  assign n72780 = (n60497 & n72778) | (n60497 & n72779) | (n72778 & n72779);
  assign n40448 = ~n72777 & n72780;
  assign n40449 = x170 & x197;
  assign n40450 = n40448 & n40449;
  assign n40451 = n40448 | n40449;
  assign n40452 = ~n40450 & n40451;
  assign n60939 = n40065 | n40067;
  assign n72781 = n40452 & n60939;
  assign n72749 = n39672 | n40065;
  assign n72750 = (n40065 & n40067) | (n40065 & n72749) | (n40067 & n72749);
  assign n72782 = n40452 & n72750;
  assign n72783 = (n60538 & n72781) | (n60538 & n72782) | (n72781 & n72782);
  assign n72784 = n40452 | n60939;
  assign n72785 = n40452 | n72750;
  assign n72786 = (n60538 & n72784) | (n60538 & n72785) | (n72784 & n72785);
  assign n40455 = ~n72783 & n72786;
  assign n40456 = x169 & x198;
  assign n40457 = n40455 & n40456;
  assign n40458 = n40455 | n40456;
  assign n40459 = ~n40457 & n40458;
  assign n60936 = n40072 | n40074;
  assign n60976 = n40459 & n60936;
  assign n60977 = n40072 & n40459;
  assign n60978 = (n72682 & n60976) | (n72682 & n60977) | (n60976 & n60977);
  assign n60979 = n40459 | n60936;
  assign n60980 = n40072 | n40459;
  assign n60981 = (n72682 & n60979) | (n72682 & n60980) | (n60979 & n60980);
  assign n40462 = ~n60978 & n60981;
  assign n40463 = x168 & x199;
  assign n40464 = n40462 & n40463;
  assign n40465 = n40462 | n40463;
  assign n40466 = ~n40464 & n40465;
  assign n60982 = n40079 & n40466;
  assign n72787 = (n40466 & n60763) | (n40466 & n60982) | (n60763 & n60982);
  assign n72788 = (n40466 & n60762) | (n40466 & n60982) | (n60762 & n60982);
  assign n72789 = (n60492 & n72787) | (n60492 & n72788) | (n72787 & n72788);
  assign n60984 = n40079 | n40466;
  assign n72790 = n60763 | n60984;
  assign n72791 = n60762 | n60984;
  assign n72792 = (n60492 & n72790) | (n60492 & n72791) | (n72790 & n72791);
  assign n40469 = ~n72789 & n72792;
  assign n40470 = x167 & x200;
  assign n40471 = n40469 & n40470;
  assign n40472 = n40469 | n40470;
  assign n40473 = ~n40471 & n40472;
  assign n60934 = n40086 | n40088;
  assign n72793 = n40473 & n60934;
  assign n72747 = n39693 | n40086;
  assign n72748 = (n40086 & n40088) | (n40086 & n72747) | (n40088 & n72747);
  assign n72794 = n40473 & n72748;
  assign n72795 = (n60548 & n72793) | (n60548 & n72794) | (n72793 & n72794);
  assign n72796 = n40473 | n60934;
  assign n72797 = n40473 | n72748;
  assign n72798 = (n60548 & n72796) | (n60548 & n72797) | (n72796 & n72797);
  assign n40476 = ~n72795 & n72798;
  assign n40477 = x166 & x201;
  assign n40478 = n40476 & n40477;
  assign n40479 = n40476 | n40477;
  assign n40480 = ~n40478 & n40479;
  assign n60931 = n40093 | n40095;
  assign n60986 = n40480 & n60931;
  assign n60987 = n40093 & n40480;
  assign n60988 = (n72677 & n60986) | (n72677 & n60987) | (n60986 & n60987);
  assign n60989 = n40480 | n60931;
  assign n60990 = n40093 | n40480;
  assign n60991 = (n72677 & n60989) | (n72677 & n60990) | (n60989 & n60990);
  assign n40483 = ~n60988 & n60991;
  assign n40484 = x165 & x202;
  assign n40485 = n40483 & n40484;
  assign n40486 = n40483 | n40484;
  assign n40487 = ~n40485 & n40486;
  assign n60992 = n40100 & n40487;
  assign n72799 = (n40487 & n60773) | (n40487 & n60992) | (n60773 & n60992);
  assign n72800 = (n40487 & n60772) | (n40487 & n60992) | (n60772 & n60992);
  assign n72801 = (n60487 & n72799) | (n60487 & n72800) | (n72799 & n72800);
  assign n60994 = n40100 | n40487;
  assign n72802 = n60773 | n60994;
  assign n72803 = n60772 | n60994;
  assign n72804 = (n60487 & n72802) | (n60487 & n72803) | (n72802 & n72803);
  assign n40490 = ~n72801 & n72804;
  assign n40491 = x164 & x203;
  assign n40492 = n40490 & n40491;
  assign n40493 = n40490 | n40491;
  assign n40494 = ~n40492 & n40493;
  assign n60929 = n40107 | n40109;
  assign n72805 = n40494 & n60929;
  assign n72745 = n39714 | n40107;
  assign n72746 = (n40107 & n40109) | (n40107 & n72745) | (n40109 & n72745);
  assign n72806 = n40494 & n72746;
  assign n72807 = (n60558 & n72805) | (n60558 & n72806) | (n72805 & n72806);
  assign n72808 = n40494 | n60929;
  assign n72809 = n40494 | n72746;
  assign n72810 = (n60558 & n72808) | (n60558 & n72809) | (n72808 & n72809);
  assign n40497 = ~n72807 & n72810;
  assign n40498 = x163 & x204;
  assign n40499 = n40497 & n40498;
  assign n40500 = n40497 | n40498;
  assign n40501 = ~n40499 & n40500;
  assign n60926 = n40114 | n40116;
  assign n60996 = n40501 & n60926;
  assign n60997 = n40114 & n40501;
  assign n60998 = (n72672 & n60996) | (n72672 & n60997) | (n60996 & n60997);
  assign n60999 = n40501 | n60926;
  assign n61000 = n40114 | n40501;
  assign n61001 = (n72672 & n60999) | (n72672 & n61000) | (n60999 & n61000);
  assign n40504 = ~n60998 & n61001;
  assign n40505 = x162 & x205;
  assign n40506 = n40504 & n40505;
  assign n40507 = n40504 | n40505;
  assign n40508 = ~n40506 & n40507;
  assign n61002 = n40121 & n40508;
  assign n72811 = (n40508 & n60783) | (n40508 & n61002) | (n60783 & n61002);
  assign n72812 = (n40508 & n60782) | (n40508 & n61002) | (n60782 & n61002);
  assign n72813 = (n72559 & n72811) | (n72559 & n72812) | (n72811 & n72812);
  assign n61004 = n40121 | n40508;
  assign n72814 = n60783 | n61004;
  assign n72815 = n60782 | n61004;
  assign n72816 = (n72559 & n72814) | (n72559 & n72815) | (n72814 & n72815);
  assign n40511 = ~n72813 & n72816;
  assign n40512 = x161 & x206;
  assign n40513 = n40511 & n40512;
  assign n40514 = n40511 | n40512;
  assign n40515 = ~n40513 & n40514;
  assign n40516 = n72744 & n40515;
  assign n40517 = n72744 | n40515;
  assign n40518 = ~n40516 & n40517;
  assign n40519 = x160 & x207;
  assign n40520 = n40518 & n40519;
  assign n40521 = n40518 | n40519;
  assign n40522 = ~n40520 & n40521;
  assign n60921 = n40135 | n40137;
  assign n61006 = n40522 & n60921;
  assign n61007 = n40135 & n40522;
  assign n61008 = (n72667 & n61006) | (n72667 & n61007) | (n61006 & n61007);
  assign n61009 = n40522 | n60921;
  assign n61010 = n40135 | n40522;
  assign n61011 = (n72667 & n61009) | (n72667 & n61010) | (n61009 & n61010);
  assign n40525 = ~n61008 & n61011;
  assign n40526 = x159 & x208;
  assign n40527 = n40525 & n40526;
  assign n40528 = n40525 | n40526;
  assign n40529 = ~n40527 & n40528;
  assign n61012 = n40142 & n40529;
  assign n72817 = (n40529 & n60793) | (n40529 & n61012) | (n60793 & n61012);
  assign n72818 = (n40529 & n60792) | (n40529 & n61012) | (n60792 & n61012);
  assign n72819 = (n72554 & n72817) | (n72554 & n72818) | (n72817 & n72818);
  assign n61014 = n40142 | n40529;
  assign n72820 = n60793 | n61014;
  assign n72821 = n60792 | n61014;
  assign n72822 = (n72554 & n72820) | (n72554 & n72821) | (n72820 & n72821);
  assign n40532 = ~n72819 & n72822;
  assign n40533 = x158 & x209;
  assign n40534 = n40532 & n40533;
  assign n40535 = n40532 | n40533;
  assign n40536 = ~n40534 & n40535;
  assign n40537 = n72739 & n40536;
  assign n40538 = n72739 | n40536;
  assign n40539 = ~n40537 & n40538;
  assign n40540 = x157 & x210;
  assign n40541 = n40539 & n40540;
  assign n40542 = n40539 | n40540;
  assign n40543 = ~n40541 & n40542;
  assign n60916 = n40156 | n40158;
  assign n61016 = n40543 & n60916;
  assign n61017 = n40156 & n40543;
  assign n61018 = (n60700 & n61016) | (n60700 & n61017) | (n61016 & n61017);
  assign n61019 = n40543 | n60916;
  assign n61020 = n40156 | n40543;
  assign n61021 = (n60700 & n61019) | (n60700 & n61020) | (n61019 & n61020);
  assign n40546 = ~n61018 & n61021;
  assign n40547 = x156 & x211;
  assign n40548 = n40546 & n40547;
  assign n40549 = n40546 | n40547;
  assign n40550 = ~n40548 & n40549;
  assign n61022 = n40163 & n40550;
  assign n61023 = (n40550 & n72719) | (n40550 & n61022) | (n72719 & n61022);
  assign n61024 = n40163 | n40550;
  assign n61025 = n72719 | n61024;
  assign n40553 = ~n61023 & n61025;
  assign n40554 = x155 & x212;
  assign n40555 = n40553 & n40554;
  assign n40556 = n40553 | n40554;
  assign n40557 = ~n40555 & n40556;
  assign n61026 = n40170 & n40557;
  assign n61027 = (n40557 & n60807) | (n40557 & n61026) | (n60807 & n61026);
  assign n61028 = n40170 | n40557;
  assign n61029 = n60807 | n61028;
  assign n40560 = ~n61027 & n61029;
  assign n40561 = x154 & x213;
  assign n40562 = n40560 & n40561;
  assign n40563 = n40560 | n40561;
  assign n40564 = ~n40562 & n40563;
  assign n61030 = n40177 & n40564;
  assign n61031 = (n40564 & n60811) | (n40564 & n61030) | (n60811 & n61030);
  assign n61032 = n40177 | n40564;
  assign n61033 = n60811 | n61032;
  assign n40567 = ~n61031 & n61033;
  assign n40568 = x153 & x214;
  assign n40569 = n40567 & n40568;
  assign n40570 = n40567 | n40568;
  assign n40571 = ~n40569 & n40570;
  assign n61034 = n40184 & n40571;
  assign n61035 = (n40571 & n60815) | (n40571 & n61034) | (n60815 & n61034);
  assign n61036 = n40184 | n40571;
  assign n61037 = n60815 | n61036;
  assign n40574 = ~n61035 & n61037;
  assign n40575 = x152 & x215;
  assign n40576 = n40574 & n40575;
  assign n40577 = n40574 | n40575;
  assign n40578 = ~n40576 & n40577;
  assign n61038 = n40191 & n40578;
  assign n61039 = (n40578 & n60819) | (n40578 & n61038) | (n60819 & n61038);
  assign n61040 = n40191 | n40578;
  assign n61041 = n60819 | n61040;
  assign n40581 = ~n61039 & n61041;
  assign n40582 = x151 & x216;
  assign n40583 = n40581 & n40582;
  assign n40584 = n40581 | n40582;
  assign n40585 = ~n40583 & n40584;
  assign n61042 = n40198 & n40585;
  assign n61043 = (n40585 & n60823) | (n40585 & n61042) | (n60823 & n61042);
  assign n61044 = n40198 | n40585;
  assign n61045 = n60823 | n61044;
  assign n40588 = ~n61043 & n61045;
  assign n40589 = x150 & x217;
  assign n40590 = n40588 & n40589;
  assign n40591 = n40588 | n40589;
  assign n40592 = ~n40590 & n40591;
  assign n61046 = n40205 & n40592;
  assign n61047 = (n40592 & n60827) | (n40592 & n61046) | (n60827 & n61046);
  assign n61048 = n40205 | n40592;
  assign n61049 = n60827 | n61048;
  assign n40595 = ~n61047 & n61049;
  assign n40596 = x149 & x218;
  assign n40597 = n40595 & n40596;
  assign n40598 = n40595 | n40596;
  assign n40599 = ~n40597 & n40598;
  assign n61050 = n40212 & n40599;
  assign n61051 = (n40599 & n60831) | (n40599 & n61050) | (n60831 & n61050);
  assign n61052 = n40212 | n40599;
  assign n61053 = n60831 | n61052;
  assign n40602 = ~n61051 & n61053;
  assign n40603 = x148 & x219;
  assign n40604 = n40602 & n40603;
  assign n40605 = n40602 | n40603;
  assign n40606 = ~n40604 & n40605;
  assign n61054 = n40219 & n40606;
  assign n61055 = (n40606 & n60835) | (n40606 & n61054) | (n60835 & n61054);
  assign n61056 = n40219 | n40606;
  assign n61057 = n60835 | n61056;
  assign n40609 = ~n61055 & n61057;
  assign n40610 = x147 & x220;
  assign n40611 = n40609 & n40610;
  assign n40612 = n40609 | n40610;
  assign n40613 = ~n40611 & n40612;
  assign n61058 = n40226 & n40613;
  assign n61059 = (n40613 & n60839) | (n40613 & n61058) | (n60839 & n61058);
  assign n61060 = n40226 | n40613;
  assign n61061 = n60839 | n61060;
  assign n40616 = ~n61059 & n61061;
  assign n40617 = x146 & x221;
  assign n40618 = n40616 & n40617;
  assign n40619 = n40616 | n40617;
  assign n40620 = ~n40618 & n40619;
  assign n61062 = n40233 & n40620;
  assign n61063 = (n40620 & n60843) | (n40620 & n61062) | (n60843 & n61062);
  assign n61064 = n40233 | n40620;
  assign n61065 = n60843 | n61064;
  assign n40623 = ~n61063 & n61065;
  assign n40624 = x145 & x222;
  assign n40625 = n40623 & n40624;
  assign n40626 = n40623 | n40624;
  assign n40627 = ~n40625 & n40626;
  assign n61066 = n40240 & n40627;
  assign n61067 = (n40627 & n60847) | (n40627 & n61066) | (n60847 & n61066);
  assign n61068 = n40240 | n40627;
  assign n61069 = n60847 | n61068;
  assign n40630 = ~n61067 & n61069;
  assign n40631 = x144 & x223;
  assign n40632 = n40630 & n40631;
  assign n40633 = n40630 | n40631;
  assign n40634 = ~n40632 & n40633;
  assign n61070 = n40247 & n40634;
  assign n61071 = (n40634 & n60851) | (n40634 & n61070) | (n60851 & n61070);
  assign n61072 = n40247 | n40634;
  assign n61073 = n60851 | n61072;
  assign n40637 = ~n61071 & n61073;
  assign n40638 = x143 & x224;
  assign n40639 = n40637 & n40638;
  assign n40640 = n40637 | n40638;
  assign n40641 = ~n40639 & n40640;
  assign n61074 = n40254 & n40641;
  assign n61075 = (n40641 & n60855) | (n40641 & n61074) | (n60855 & n61074);
  assign n61076 = n40254 | n40641;
  assign n61077 = n60855 | n61076;
  assign n40644 = ~n61075 & n61077;
  assign n40645 = x142 & x225;
  assign n40646 = n40644 & n40645;
  assign n40647 = n40644 | n40645;
  assign n40648 = ~n40646 & n40647;
  assign n61078 = n40261 & n40648;
  assign n61079 = (n40648 & n60859) | (n40648 & n61078) | (n60859 & n61078);
  assign n61080 = n40261 | n40648;
  assign n61081 = n60859 | n61080;
  assign n40651 = ~n61079 & n61081;
  assign n40652 = x141 & x226;
  assign n40653 = n40651 & n40652;
  assign n40654 = n40651 | n40652;
  assign n40655 = ~n40653 & n40654;
  assign n61082 = n40268 & n40655;
  assign n61083 = (n40655 & n60863) | (n40655 & n61082) | (n60863 & n61082);
  assign n61084 = n40268 | n40655;
  assign n61085 = n60863 | n61084;
  assign n40658 = ~n61083 & n61085;
  assign n40659 = x140 & x227;
  assign n40660 = n40658 & n40659;
  assign n40661 = n40658 | n40659;
  assign n40662 = ~n40660 & n40661;
  assign n61086 = n40275 & n40662;
  assign n61087 = (n40662 & n60867) | (n40662 & n61086) | (n60867 & n61086);
  assign n61088 = n40275 | n40662;
  assign n61089 = n60867 | n61088;
  assign n40665 = ~n61087 & n61089;
  assign n40666 = x139 & x228;
  assign n40667 = n40665 & n40666;
  assign n40668 = n40665 | n40666;
  assign n40669 = ~n40667 & n40668;
  assign n61090 = n40282 & n40669;
  assign n61091 = (n40669 & n60871) | (n40669 & n61090) | (n60871 & n61090);
  assign n61092 = n40282 | n40669;
  assign n61093 = n60871 | n61092;
  assign n40672 = ~n61091 & n61093;
  assign n40673 = x138 & x229;
  assign n40674 = n40672 & n40673;
  assign n40675 = n40672 | n40673;
  assign n40676 = ~n40674 & n40675;
  assign n61094 = n40289 & n40676;
  assign n61095 = (n40676 & n60875) | (n40676 & n61094) | (n60875 & n61094);
  assign n61096 = n40289 | n40676;
  assign n61097 = n60875 | n61096;
  assign n40679 = ~n61095 & n61097;
  assign n40680 = x137 & x230;
  assign n40681 = n40679 & n40680;
  assign n40682 = n40679 | n40680;
  assign n40683 = ~n40681 & n40682;
  assign n61098 = n40296 & n40683;
  assign n61099 = (n40683 & n60879) | (n40683 & n61098) | (n60879 & n61098);
  assign n61100 = n40296 | n40683;
  assign n61101 = n60879 | n61100;
  assign n40686 = ~n61099 & n61101;
  assign n40687 = x136 & x231;
  assign n40688 = n40686 & n40687;
  assign n40689 = n40686 | n40687;
  assign n40690 = ~n40688 & n40689;
  assign n61102 = n40303 & n40690;
  assign n61103 = (n40690 & n60883) | (n40690 & n61102) | (n60883 & n61102);
  assign n61104 = n40303 | n40690;
  assign n61105 = n60883 | n61104;
  assign n40693 = ~n61103 & n61105;
  assign n40694 = x135 & x232;
  assign n40695 = n40693 & n40694;
  assign n40696 = n40693 | n40694;
  assign n40697 = ~n40695 & n40696;
  assign n61106 = n40310 & n40697;
  assign n61107 = (n40697 & n60887) | (n40697 & n61106) | (n60887 & n61106);
  assign n61108 = n40310 | n40697;
  assign n61109 = n60887 | n61108;
  assign n40700 = ~n61107 & n61109;
  assign n40701 = x134 & x233;
  assign n40702 = n40700 & n40701;
  assign n40703 = n40700 | n40701;
  assign n40704 = ~n40702 & n40703;
  assign n61110 = n40317 & n40704;
  assign n61111 = (n40704 & n60891) | (n40704 & n61110) | (n60891 & n61110);
  assign n61112 = n40317 | n40704;
  assign n61113 = n60891 | n61112;
  assign n40707 = ~n61111 & n61113;
  assign n40708 = x133 & x234;
  assign n40709 = n40707 & n40708;
  assign n40710 = n40707 | n40708;
  assign n40711 = ~n40709 & n40710;
  assign n61114 = n40324 & n40711;
  assign n61115 = (n40711 & n60895) | (n40711 & n61114) | (n60895 & n61114);
  assign n61116 = n40324 | n40711;
  assign n61117 = n60895 | n61116;
  assign n40714 = ~n61115 & n61117;
  assign n40715 = x132 & x235;
  assign n40716 = n40714 & n40715;
  assign n40717 = n40714 | n40715;
  assign n40718 = ~n40716 & n40717;
  assign n61118 = n40331 & n40718;
  assign n61119 = (n40718 & n60899) | (n40718 & n61118) | (n60899 & n61118);
  assign n61120 = n40331 | n40718;
  assign n61121 = n60899 | n61120;
  assign n40721 = ~n61119 & n61121;
  assign n40722 = x131 & x236;
  assign n40723 = n40721 & n40722;
  assign n40724 = n40721 | n40722;
  assign n40725 = ~n40723 & n40724;
  assign n61122 = n40338 & n40725;
  assign n61123 = (n40725 & n60903) | (n40725 & n61122) | (n60903 & n61122);
  assign n61124 = n40338 | n40725;
  assign n61125 = n60903 | n61124;
  assign n40728 = ~n61123 & n61125;
  assign n40729 = x130 & x237;
  assign n40730 = n40728 & n40729;
  assign n40731 = n40728 | n40729;
  assign n40732 = ~n40730 & n40731;
  assign n61126 = n40345 & n40732;
  assign n61127 = (n40732 & n60908) | (n40732 & n61126) | (n60908 & n61126);
  assign n61128 = n40345 | n40732;
  assign n61129 = n60908 | n61128;
  assign n40735 = ~n61127 & n61129;
  assign n40736 = x129 & x238;
  assign n40737 = n40735 & n40736;
  assign n40738 = n40735 | n40736;
  assign n40739 = ~n40737 & n40738;
  assign n60914 = n40352 | n40354;
  assign n61130 = n40739 & n60914;
  assign n61131 = n40352 & n40739;
  assign n61132 = (n60695 & n61130) | (n60695 & n61131) | (n61130 & n61131);
  assign n61133 = n40739 | n60914;
  assign n61134 = n40352 | n40739;
  assign n61135 = (n60695 & n61133) | (n60695 & n61134) | (n61133 & n61134);
  assign n40742 = ~n61132 & n61135;
  assign n40743 = x128 & x239;
  assign n40744 = n40742 & n40743;
  assign n40745 = n40742 | n40743;
  assign n40746 = ~n40744 & n40745;
  assign n60912 = n40359 | n40361;
  assign n72823 = n40746 & n60912;
  assign n72824 = n40359 & n40746;
  assign n72825 = (n60693 & n72823) | (n60693 & n72824) | (n72823 & n72824);
  assign n72826 = n40746 | n60912;
  assign n72827 = n40359 | n40746;
  assign n72828 = (n60693 & n72826) | (n60693 & n72827) | (n72826 & n72827);
  assign n40749 = ~n72825 & n72828;
  assign n60913 = (n40359 & n60693) | (n40359 & n60912) | (n60693 & n60912);
  assign n61144 = n40527 | n40529;
  assign n72831 = n40142 | n40527;
  assign n72832 = (n40527 & n40529) | (n40527 & n72831) | (n40529 & n72831);
  assign n72833 = (n60793 & n61144) | (n60793 & n72832) | (n61144 & n72832);
  assign n72834 = (n60792 & n61144) | (n60792 & n72832) | (n61144 & n72832);
  assign n72835 = (n72554 & n72833) | (n72554 & n72834) | (n72833 & n72834);
  assign n61149 = n40506 | n40508;
  assign n72836 = n40121 | n40506;
  assign n72837 = (n40506 & n40508) | (n40506 & n72836) | (n40508 & n72836);
  assign n72838 = (n60783 & n61149) | (n60783 & n72837) | (n61149 & n72837);
  assign n72839 = (n60782 & n61149) | (n60782 & n72837) | (n61149 & n72837);
  assign n72840 = (n72559 & n72838) | (n72559 & n72839) | (n72838 & n72839);
  assign n60930 = (n60558 & n72746) | (n60558 & n60929) | (n72746 & n60929);
  assign n61154 = n40485 | n40487;
  assign n72841 = n40100 | n40485;
  assign n72842 = (n40485 & n40487) | (n40485 & n72841) | (n40487 & n72841);
  assign n72843 = (n60773 & n61154) | (n60773 & n72842) | (n61154 & n72842);
  assign n72844 = (n60772 & n61154) | (n60772 & n72842) | (n61154 & n72842);
  assign n72845 = (n60487 & n72843) | (n60487 & n72844) | (n72843 & n72844);
  assign n60935 = (n60548 & n72748) | (n60548 & n60934) | (n72748 & n60934);
  assign n61159 = n40464 | n40466;
  assign n72846 = n40079 | n40464;
  assign n72847 = (n40464 & n40466) | (n40464 & n72846) | (n40466 & n72846);
  assign n72848 = (n60763 & n61159) | (n60763 & n72847) | (n61159 & n72847);
  assign n72849 = (n60762 & n61159) | (n60762 & n72847) | (n61159 & n72847);
  assign n72850 = (n60492 & n72848) | (n60492 & n72849) | (n72848 & n72849);
  assign n60940 = (n60538 & n72750) | (n60538 & n60939) | (n72750 & n60939);
  assign n61164 = n40443 | n40445;
  assign n72851 = n40058 | n40443;
  assign n72852 = (n40443 & n40445) | (n40443 & n72851) | (n40445 & n72851);
  assign n72853 = (n60753 & n61164) | (n60753 & n72852) | (n61164 & n72852);
  assign n72854 = (n60752 & n61164) | (n60752 & n72852) | (n61164 & n72852);
  assign n72855 = (n60497 & n72853) | (n60497 & n72854) | (n72853 & n72854);
  assign n60945 = (n60528 & n72752) | (n60528 & n60944) | (n72752 & n60944);
  assign n61169 = n40422 | n40424;
  assign n72856 = n40037 | n40422;
  assign n72857 = (n40422 & n40424) | (n40422 & n72856) | (n40424 & n72856);
  assign n72858 = (n60743 & n61169) | (n60743 & n72857) | (n61169 & n72857);
  assign n72859 = (n60742 & n61169) | (n60742 & n72857) | (n61169 & n72857);
  assign n72860 = (n60502 & n72858) | (n60502 & n72859) | (n72858 & n72859);
  assign n40798 = x175 & x193;
  assign n72861 = n40798 & n72753;
  assign n72862 = n40798 & n72756;
  assign n72863 = (n60733 & n72861) | (n60733 & n72862) | (n72861 & n72862);
  assign n72864 = (n40798 & n72761) | (n40798 & n72863) | (n72761 & n72863);
  assign n72865 = (n40798 & n60957) | (n40798 & n72863) | (n60957 & n72863);
  assign n72866 = (n72692 & n72864) | (n72692 & n72865) | (n72864 & n72865);
  assign n72867 = n40798 | n72753;
  assign n72868 = n40798 | n72756;
  assign n72869 = (n60733 & n72867) | (n60733 & n72868) | (n72867 & n72868);
  assign n72870 = n72761 | n72869;
  assign n72871 = n60957 | n72869;
  assign n72872 = (n72692 & n72870) | (n72692 & n72871) | (n72870 & n72871);
  assign n40801 = ~n72866 & n72872;
  assign n40802 = n72860 & n40801;
  assign n40803 = n72860 | n40801;
  assign n40804 = ~n40802 & n40803;
  assign n40805 = x174 & x194;
  assign n40806 = n40804 & n40805;
  assign n40807 = n40804 | n40805;
  assign n40808 = ~n40806 & n40807;
  assign n61166 = n40429 | n40431;
  assign n61175 = n40808 & n61166;
  assign n61176 = n40429 & n40808;
  assign n61177 = (n60945 & n61175) | (n60945 & n61176) | (n61175 & n61176);
  assign n61178 = n40808 | n61166;
  assign n61179 = n40429 | n40808;
  assign n61180 = (n60945 & n61178) | (n60945 & n61179) | (n61178 & n61179);
  assign n40811 = ~n61177 & n61180;
  assign n40812 = x173 & x195;
  assign n40813 = n40811 & n40812;
  assign n40814 = n40811 | n40812;
  assign n40815 = ~n40813 & n40814;
  assign n61181 = n40436 & n40815;
  assign n61182 = (n40815 & n60968) | (n40815 & n61181) | (n60968 & n61181);
  assign n61183 = n40436 | n40815;
  assign n61184 = n60968 | n61183;
  assign n40818 = ~n61182 & n61184;
  assign n40819 = x172 & x196;
  assign n40820 = n40818 & n40819;
  assign n40821 = n40818 | n40819;
  assign n40822 = ~n40820 & n40821;
  assign n40823 = n72855 & n40822;
  assign n40824 = n72855 | n40822;
  assign n40825 = ~n40823 & n40824;
  assign n40826 = x171 & x197;
  assign n40827 = n40825 & n40826;
  assign n40828 = n40825 | n40826;
  assign n40829 = ~n40827 & n40828;
  assign n61161 = n40450 | n40452;
  assign n61185 = n40829 & n61161;
  assign n61186 = n40450 & n40829;
  assign n61187 = (n60940 & n61185) | (n60940 & n61186) | (n61185 & n61186);
  assign n61188 = n40829 | n61161;
  assign n61189 = n40450 | n40829;
  assign n61190 = (n60940 & n61188) | (n60940 & n61189) | (n61188 & n61189);
  assign n40832 = ~n61187 & n61190;
  assign n40833 = x170 & x198;
  assign n40834 = n40832 & n40833;
  assign n40835 = n40832 | n40833;
  assign n40836 = ~n40834 & n40835;
  assign n61191 = n40457 & n40836;
  assign n61192 = (n40836 & n60978) | (n40836 & n61191) | (n60978 & n61191);
  assign n61193 = n40457 | n40836;
  assign n61194 = n60978 | n61193;
  assign n40839 = ~n61192 & n61194;
  assign n40840 = x169 & x199;
  assign n40841 = n40839 & n40840;
  assign n40842 = n40839 | n40840;
  assign n40843 = ~n40841 & n40842;
  assign n40844 = n72850 & n40843;
  assign n40845 = n72850 | n40843;
  assign n40846 = ~n40844 & n40845;
  assign n40847 = x168 & x200;
  assign n40848 = n40846 & n40847;
  assign n40849 = n40846 | n40847;
  assign n40850 = ~n40848 & n40849;
  assign n61156 = n40471 | n40473;
  assign n61195 = n40850 & n61156;
  assign n61196 = n40471 & n40850;
  assign n61197 = (n60935 & n61195) | (n60935 & n61196) | (n61195 & n61196);
  assign n61198 = n40850 | n61156;
  assign n61199 = n40471 | n40850;
  assign n61200 = (n60935 & n61198) | (n60935 & n61199) | (n61198 & n61199);
  assign n40853 = ~n61197 & n61200;
  assign n40854 = x167 & x201;
  assign n40855 = n40853 & n40854;
  assign n40856 = n40853 | n40854;
  assign n40857 = ~n40855 & n40856;
  assign n61201 = n40478 & n40857;
  assign n61202 = (n40857 & n60988) | (n40857 & n61201) | (n60988 & n61201);
  assign n61203 = n40478 | n40857;
  assign n61204 = n60988 | n61203;
  assign n40860 = ~n61202 & n61204;
  assign n40861 = x166 & x202;
  assign n40862 = n40860 & n40861;
  assign n40863 = n40860 | n40861;
  assign n40864 = ~n40862 & n40863;
  assign n40865 = n72845 & n40864;
  assign n40866 = n72845 | n40864;
  assign n40867 = ~n40865 & n40866;
  assign n40868 = x165 & x203;
  assign n40869 = n40867 & n40868;
  assign n40870 = n40867 | n40868;
  assign n40871 = ~n40869 & n40870;
  assign n61151 = n40492 | n40494;
  assign n61205 = n40871 & n61151;
  assign n61206 = n40492 & n40871;
  assign n61207 = (n60930 & n61205) | (n60930 & n61206) | (n61205 & n61206);
  assign n61208 = n40871 | n61151;
  assign n61209 = n40492 | n40871;
  assign n61210 = (n60930 & n61208) | (n60930 & n61209) | (n61208 & n61209);
  assign n40874 = ~n61207 & n61210;
  assign n40875 = x164 & x204;
  assign n40876 = n40874 & n40875;
  assign n40877 = n40874 | n40875;
  assign n40878 = ~n40876 & n40877;
  assign n61211 = n40499 & n40878;
  assign n61212 = (n40878 & n60998) | (n40878 & n61211) | (n60998 & n61211);
  assign n61213 = n40499 | n40878;
  assign n61214 = n60998 | n61213;
  assign n40881 = ~n61212 & n61214;
  assign n40882 = x163 & x205;
  assign n40883 = n40881 & n40882;
  assign n40884 = n40881 | n40882;
  assign n40885 = ~n40883 & n40884;
  assign n40886 = n72840 & n40885;
  assign n40887 = n72840 | n40885;
  assign n40888 = ~n40886 & n40887;
  assign n40889 = x162 & x206;
  assign n40890 = n40888 & n40889;
  assign n40891 = n40888 | n40889;
  assign n40892 = ~n40890 & n40891;
  assign n61146 = n40513 | n40515;
  assign n61215 = n40892 & n61146;
  assign n61216 = n40513 & n40892;
  assign n61217 = (n72744 & n61215) | (n72744 & n61216) | (n61215 & n61216);
  assign n61218 = n40892 | n61146;
  assign n61219 = n40513 | n40892;
  assign n61220 = (n72744 & n61218) | (n72744 & n61219) | (n61218 & n61219);
  assign n40895 = ~n61217 & n61220;
  assign n40896 = x161 & x207;
  assign n40897 = n40895 & n40896;
  assign n40898 = n40895 | n40896;
  assign n40899 = ~n40897 & n40898;
  assign n61221 = n40520 & n40899;
  assign n72873 = (n40899 & n61007) | (n40899 & n61221) | (n61007 & n61221);
  assign n72874 = (n40899 & n61006) | (n40899 & n61221) | (n61006 & n61221);
  assign n72875 = (n72667 & n72873) | (n72667 & n72874) | (n72873 & n72874);
  assign n61223 = n40520 | n40899;
  assign n72876 = n61007 | n61223;
  assign n72877 = n61006 | n61223;
  assign n72878 = (n72667 & n72876) | (n72667 & n72877) | (n72876 & n72877);
  assign n40902 = ~n72875 & n72878;
  assign n40903 = x160 & x208;
  assign n40904 = n40902 & n40903;
  assign n40905 = n40902 | n40903;
  assign n40906 = ~n40904 & n40905;
  assign n40907 = n72835 & n40906;
  assign n40908 = n72835 | n40906;
  assign n40909 = ~n40907 & n40908;
  assign n40910 = x159 & x209;
  assign n40911 = n40909 & n40910;
  assign n40912 = n40909 | n40910;
  assign n40913 = ~n40911 & n40912;
  assign n61141 = n40534 | n40536;
  assign n61225 = n40913 & n61141;
  assign n61226 = n40534 & n40913;
  assign n61227 = (n72739 & n61225) | (n72739 & n61226) | (n61225 & n61226);
  assign n61228 = n40913 | n61141;
  assign n61229 = n40534 | n40913;
  assign n61230 = (n72739 & n61228) | (n72739 & n61229) | (n61228 & n61229);
  assign n40916 = ~n61227 & n61230;
  assign n40917 = x158 & x210;
  assign n40918 = n40916 & n40917;
  assign n40919 = n40916 | n40917;
  assign n40920 = ~n40918 & n40919;
  assign n61231 = n40541 & n40920;
  assign n72879 = (n40920 & n61017) | (n40920 & n61231) | (n61017 & n61231);
  assign n72880 = (n40920 & n61016) | (n40920 & n61231) | (n61016 & n61231);
  assign n72881 = (n60700 & n72879) | (n60700 & n72880) | (n72879 & n72880);
  assign n61233 = n40541 | n40920;
  assign n72882 = n61017 | n61233;
  assign n72883 = n61016 | n61233;
  assign n72884 = (n60700 & n72882) | (n60700 & n72883) | (n72882 & n72883);
  assign n40923 = ~n72881 & n72884;
  assign n40924 = x157 & x211;
  assign n40925 = n40923 & n40924;
  assign n40926 = n40923 | n40924;
  assign n40927 = ~n40925 & n40926;
  assign n61139 = n40548 | n40550;
  assign n72885 = n40927 & n61139;
  assign n72829 = n40163 | n40548;
  assign n72830 = (n40548 & n40550) | (n40548 & n72829) | (n40550 & n72829);
  assign n72886 = n40927 & n72830;
  assign n72887 = (n72719 & n72885) | (n72719 & n72886) | (n72885 & n72886);
  assign n72888 = n40927 | n61139;
  assign n72889 = n40927 | n72830;
  assign n72890 = (n72719 & n72888) | (n72719 & n72889) | (n72888 & n72889);
  assign n40930 = ~n72887 & n72890;
  assign n40931 = x156 & x212;
  assign n40932 = n40930 & n40931;
  assign n40933 = n40930 | n40931;
  assign n40934 = ~n40932 & n40933;
  assign n61235 = n40555 & n40934;
  assign n72891 = (n40934 & n61026) | (n40934 & n61235) | (n61026 & n61235);
  assign n72892 = (n40557 & n40934) | (n40557 & n61235) | (n40934 & n61235);
  assign n72893 = (n60807 & n72891) | (n60807 & n72892) | (n72891 & n72892);
  assign n61237 = n40555 | n40934;
  assign n72894 = n61026 | n61237;
  assign n72895 = n40557 | n61237;
  assign n72896 = (n60807 & n72894) | (n60807 & n72895) | (n72894 & n72895);
  assign n40937 = ~n72893 & n72896;
  assign n40938 = x155 & x213;
  assign n40939 = n40937 & n40938;
  assign n40940 = n40937 | n40938;
  assign n40941 = ~n40939 & n40940;
  assign n61239 = n40562 & n40941;
  assign n61240 = (n40941 & n61031) | (n40941 & n61239) | (n61031 & n61239);
  assign n61241 = n40562 | n40941;
  assign n61242 = n61031 | n61241;
  assign n40944 = ~n61240 & n61242;
  assign n40945 = x154 & x214;
  assign n40946 = n40944 & n40945;
  assign n40947 = n40944 | n40945;
  assign n40948 = ~n40946 & n40947;
  assign n61243 = n40569 & n40948;
  assign n61244 = (n40948 & n61035) | (n40948 & n61243) | (n61035 & n61243);
  assign n61245 = n40569 | n40948;
  assign n61246 = n61035 | n61245;
  assign n40951 = ~n61244 & n61246;
  assign n40952 = x153 & x215;
  assign n40953 = n40951 & n40952;
  assign n40954 = n40951 | n40952;
  assign n40955 = ~n40953 & n40954;
  assign n61247 = n40576 & n40955;
  assign n61248 = (n40955 & n61039) | (n40955 & n61247) | (n61039 & n61247);
  assign n61249 = n40576 | n40955;
  assign n61250 = n61039 | n61249;
  assign n40958 = ~n61248 & n61250;
  assign n40959 = x152 & x216;
  assign n40960 = n40958 & n40959;
  assign n40961 = n40958 | n40959;
  assign n40962 = ~n40960 & n40961;
  assign n61251 = n40583 & n40962;
  assign n61252 = (n40962 & n61043) | (n40962 & n61251) | (n61043 & n61251);
  assign n61253 = n40583 | n40962;
  assign n61254 = n61043 | n61253;
  assign n40965 = ~n61252 & n61254;
  assign n40966 = x151 & x217;
  assign n40967 = n40965 & n40966;
  assign n40968 = n40965 | n40966;
  assign n40969 = ~n40967 & n40968;
  assign n61255 = n40590 & n40969;
  assign n61256 = (n40969 & n61047) | (n40969 & n61255) | (n61047 & n61255);
  assign n61257 = n40590 | n40969;
  assign n61258 = n61047 | n61257;
  assign n40972 = ~n61256 & n61258;
  assign n40973 = x150 & x218;
  assign n40974 = n40972 & n40973;
  assign n40975 = n40972 | n40973;
  assign n40976 = ~n40974 & n40975;
  assign n61259 = n40597 & n40976;
  assign n61260 = (n40976 & n61051) | (n40976 & n61259) | (n61051 & n61259);
  assign n61261 = n40597 | n40976;
  assign n61262 = n61051 | n61261;
  assign n40979 = ~n61260 & n61262;
  assign n40980 = x149 & x219;
  assign n40981 = n40979 & n40980;
  assign n40982 = n40979 | n40980;
  assign n40983 = ~n40981 & n40982;
  assign n61263 = n40604 & n40983;
  assign n61264 = (n40983 & n61055) | (n40983 & n61263) | (n61055 & n61263);
  assign n61265 = n40604 | n40983;
  assign n61266 = n61055 | n61265;
  assign n40986 = ~n61264 & n61266;
  assign n40987 = x148 & x220;
  assign n40988 = n40986 & n40987;
  assign n40989 = n40986 | n40987;
  assign n40990 = ~n40988 & n40989;
  assign n61267 = n40611 & n40990;
  assign n61268 = (n40990 & n61059) | (n40990 & n61267) | (n61059 & n61267);
  assign n61269 = n40611 | n40990;
  assign n61270 = n61059 | n61269;
  assign n40993 = ~n61268 & n61270;
  assign n40994 = x147 & x221;
  assign n40995 = n40993 & n40994;
  assign n40996 = n40993 | n40994;
  assign n40997 = ~n40995 & n40996;
  assign n61271 = n40618 & n40997;
  assign n61272 = (n40997 & n61063) | (n40997 & n61271) | (n61063 & n61271);
  assign n61273 = n40618 | n40997;
  assign n61274 = n61063 | n61273;
  assign n41000 = ~n61272 & n61274;
  assign n41001 = x146 & x222;
  assign n41002 = n41000 & n41001;
  assign n41003 = n41000 | n41001;
  assign n41004 = ~n41002 & n41003;
  assign n61275 = n40625 & n41004;
  assign n61276 = (n41004 & n61067) | (n41004 & n61275) | (n61067 & n61275);
  assign n61277 = n40625 | n41004;
  assign n61278 = n61067 | n61277;
  assign n41007 = ~n61276 & n61278;
  assign n41008 = x145 & x223;
  assign n41009 = n41007 & n41008;
  assign n41010 = n41007 | n41008;
  assign n41011 = ~n41009 & n41010;
  assign n61279 = n40632 & n41011;
  assign n61280 = (n41011 & n61071) | (n41011 & n61279) | (n61071 & n61279);
  assign n61281 = n40632 | n41011;
  assign n61282 = n61071 | n61281;
  assign n41014 = ~n61280 & n61282;
  assign n41015 = x144 & x224;
  assign n41016 = n41014 & n41015;
  assign n41017 = n41014 | n41015;
  assign n41018 = ~n41016 & n41017;
  assign n61283 = n40639 & n41018;
  assign n61284 = (n41018 & n61075) | (n41018 & n61283) | (n61075 & n61283);
  assign n61285 = n40639 | n41018;
  assign n61286 = n61075 | n61285;
  assign n41021 = ~n61284 & n61286;
  assign n41022 = x143 & x225;
  assign n41023 = n41021 & n41022;
  assign n41024 = n41021 | n41022;
  assign n41025 = ~n41023 & n41024;
  assign n61287 = n40646 & n41025;
  assign n61288 = (n41025 & n61079) | (n41025 & n61287) | (n61079 & n61287);
  assign n61289 = n40646 | n41025;
  assign n61290 = n61079 | n61289;
  assign n41028 = ~n61288 & n61290;
  assign n41029 = x142 & x226;
  assign n41030 = n41028 & n41029;
  assign n41031 = n41028 | n41029;
  assign n41032 = ~n41030 & n41031;
  assign n61291 = n40653 & n41032;
  assign n61292 = (n41032 & n61083) | (n41032 & n61291) | (n61083 & n61291);
  assign n61293 = n40653 | n41032;
  assign n61294 = n61083 | n61293;
  assign n41035 = ~n61292 & n61294;
  assign n41036 = x141 & x227;
  assign n41037 = n41035 & n41036;
  assign n41038 = n41035 | n41036;
  assign n41039 = ~n41037 & n41038;
  assign n61295 = n40660 & n41039;
  assign n61296 = (n41039 & n61087) | (n41039 & n61295) | (n61087 & n61295);
  assign n61297 = n40660 | n41039;
  assign n61298 = n61087 | n61297;
  assign n41042 = ~n61296 & n61298;
  assign n41043 = x140 & x228;
  assign n41044 = n41042 & n41043;
  assign n41045 = n41042 | n41043;
  assign n41046 = ~n41044 & n41045;
  assign n61299 = n40667 & n41046;
  assign n61300 = (n41046 & n61091) | (n41046 & n61299) | (n61091 & n61299);
  assign n61301 = n40667 | n41046;
  assign n61302 = n61091 | n61301;
  assign n41049 = ~n61300 & n61302;
  assign n41050 = x139 & x229;
  assign n41051 = n41049 & n41050;
  assign n41052 = n41049 | n41050;
  assign n41053 = ~n41051 & n41052;
  assign n61303 = n40674 & n41053;
  assign n61304 = (n41053 & n61095) | (n41053 & n61303) | (n61095 & n61303);
  assign n61305 = n40674 | n41053;
  assign n61306 = n61095 | n61305;
  assign n41056 = ~n61304 & n61306;
  assign n41057 = x138 & x230;
  assign n41058 = n41056 & n41057;
  assign n41059 = n41056 | n41057;
  assign n41060 = ~n41058 & n41059;
  assign n61307 = n40681 & n41060;
  assign n61308 = (n41060 & n61099) | (n41060 & n61307) | (n61099 & n61307);
  assign n61309 = n40681 | n41060;
  assign n61310 = n61099 | n61309;
  assign n41063 = ~n61308 & n61310;
  assign n41064 = x137 & x231;
  assign n41065 = n41063 & n41064;
  assign n41066 = n41063 | n41064;
  assign n41067 = ~n41065 & n41066;
  assign n61311 = n40688 & n41067;
  assign n61312 = (n41067 & n61103) | (n41067 & n61311) | (n61103 & n61311);
  assign n61313 = n40688 | n41067;
  assign n61314 = n61103 | n61313;
  assign n41070 = ~n61312 & n61314;
  assign n41071 = x136 & x232;
  assign n41072 = n41070 & n41071;
  assign n41073 = n41070 | n41071;
  assign n41074 = ~n41072 & n41073;
  assign n61315 = n40695 & n41074;
  assign n61316 = (n41074 & n61107) | (n41074 & n61315) | (n61107 & n61315);
  assign n61317 = n40695 | n41074;
  assign n61318 = n61107 | n61317;
  assign n41077 = ~n61316 & n61318;
  assign n41078 = x135 & x233;
  assign n41079 = n41077 & n41078;
  assign n41080 = n41077 | n41078;
  assign n41081 = ~n41079 & n41080;
  assign n61319 = n40702 & n41081;
  assign n61320 = (n41081 & n61111) | (n41081 & n61319) | (n61111 & n61319);
  assign n61321 = n40702 | n41081;
  assign n61322 = n61111 | n61321;
  assign n41084 = ~n61320 & n61322;
  assign n41085 = x134 & x234;
  assign n41086 = n41084 & n41085;
  assign n41087 = n41084 | n41085;
  assign n41088 = ~n41086 & n41087;
  assign n61323 = n40709 & n41088;
  assign n61324 = (n41088 & n61115) | (n41088 & n61323) | (n61115 & n61323);
  assign n61325 = n40709 | n41088;
  assign n61326 = n61115 | n61325;
  assign n41091 = ~n61324 & n61326;
  assign n41092 = x133 & x235;
  assign n41093 = n41091 & n41092;
  assign n41094 = n41091 | n41092;
  assign n41095 = ~n41093 & n41094;
  assign n61327 = n40716 & n41095;
  assign n61328 = (n41095 & n61119) | (n41095 & n61327) | (n61119 & n61327);
  assign n61329 = n40716 | n41095;
  assign n61330 = n61119 | n61329;
  assign n41098 = ~n61328 & n61330;
  assign n41099 = x132 & x236;
  assign n41100 = n41098 & n41099;
  assign n41101 = n41098 | n41099;
  assign n41102 = ~n41100 & n41101;
  assign n61331 = n40723 & n41102;
  assign n61332 = (n41102 & n61123) | (n41102 & n61331) | (n61123 & n61331);
  assign n61333 = n40723 | n41102;
  assign n61334 = n61123 | n61333;
  assign n41105 = ~n61332 & n61334;
  assign n41106 = x131 & x237;
  assign n41107 = n41105 & n41106;
  assign n41108 = n41105 | n41106;
  assign n41109 = ~n41107 & n41108;
  assign n61335 = n40730 & n41109;
  assign n61336 = (n41109 & n61127) | (n41109 & n61335) | (n61127 & n61335);
  assign n61337 = n40730 | n41109;
  assign n61338 = n61127 | n61337;
  assign n41112 = ~n61336 & n61338;
  assign n41113 = x130 & x238;
  assign n41114 = n41112 & n41113;
  assign n41115 = n41112 | n41113;
  assign n41116 = ~n41114 & n41115;
  assign n61339 = n40737 & n41116;
  assign n61340 = (n41116 & n61132) | (n41116 & n61339) | (n61132 & n61339);
  assign n61341 = n40737 | n41116;
  assign n61342 = n61132 | n61341;
  assign n41119 = ~n61340 & n61342;
  assign n41120 = x129 & x239;
  assign n41121 = n41119 & n41120;
  assign n41122 = n41119 | n41120;
  assign n41123 = ~n41121 & n41122;
  assign n61136 = n40744 | n40746;
  assign n61343 = n41123 & n61136;
  assign n61344 = n40744 & n41123;
  assign n61345 = (n60913 & n61343) | (n60913 & n61344) | (n61343 & n61344);
  assign n61346 = n41123 | n61136;
  assign n61347 = n40744 | n41123;
  assign n61348 = (n60913 & n61346) | (n60913 & n61347) | (n61346 & n61347);
  assign n41126 = ~n61345 & n61348;
  assign n61140 = (n72719 & n72830) | (n72719 & n61139) | (n72830 & n61139);
  assign n61352 = n40918 | n40920;
  assign n72897 = n40541 | n40918;
  assign n72898 = (n40918 & n40920) | (n40918 & n72897) | (n40920 & n72897);
  assign n72899 = (n61017 & n61352) | (n61017 & n72898) | (n61352 & n72898);
  assign n72900 = (n61016 & n61352) | (n61016 & n72898) | (n61352 & n72898);
  assign n72901 = (n60700 & n72899) | (n60700 & n72900) | (n72899 & n72900);
  assign n61357 = n40897 | n40899;
  assign n72902 = n40520 | n40897;
  assign n72903 = (n40897 & n40899) | (n40897 & n72902) | (n40899 & n72902);
  assign n72904 = (n61007 & n61357) | (n61007 & n72903) | (n61357 & n72903);
  assign n72905 = (n61006 & n61357) | (n61006 & n72903) | (n61357 & n72903);
  assign n72906 = (n72667 & n72904) | (n72667 & n72905) | (n72904 & n72905);
  assign n41174 = x175 & x194;
  assign n72915 = n41174 & n72866;
  assign n72916 = (n40801 & n41174) | (n40801 & n72915) | (n41174 & n72915);
  assign n61382 = n41174 & n72866;
  assign n61383 = (n72860 & n72916) | (n72860 & n61382) | (n72916 & n61382);
  assign n72917 = n41174 | n72866;
  assign n72918 = n40801 | n72917;
  assign n61385 = n41174 | n72866;
  assign n61386 = (n72860 & n72918) | (n72860 & n61385) | (n72918 & n61385);
  assign n41177 = ~n61383 & n61386;
  assign n61387 = n40806 & n41177;
  assign n72919 = (n41177 & n61176) | (n41177 & n61387) | (n61176 & n61387);
  assign n72920 = (n41177 & n61175) | (n41177 & n61387) | (n61175 & n61387);
  assign n72921 = (n60945 & n72919) | (n60945 & n72920) | (n72919 & n72920);
  assign n61389 = n40806 | n41177;
  assign n72922 = n61176 | n61389;
  assign n72923 = n61175 | n61389;
  assign n72924 = (n60945 & n72922) | (n60945 & n72923) | (n72922 & n72923);
  assign n41180 = ~n72921 & n72924;
  assign n41181 = x174 & x195;
  assign n41182 = n41180 & n41181;
  assign n41183 = n41180 | n41181;
  assign n41184 = ~n41182 & n41183;
  assign n61377 = n40813 | n40815;
  assign n72925 = n41184 & n61377;
  assign n72913 = n40436 | n40813;
  assign n72914 = (n40813 & n40815) | (n40813 & n72913) | (n40815 & n72913);
  assign n72926 = n41184 & n72914;
  assign n72927 = (n60968 & n72925) | (n60968 & n72926) | (n72925 & n72926);
  assign n72928 = n41184 | n61377;
  assign n72929 = n41184 | n72914;
  assign n72930 = (n60968 & n72928) | (n60968 & n72929) | (n72928 & n72929);
  assign n41187 = ~n72927 & n72930;
  assign n41188 = x173 & x196;
  assign n41189 = n41187 & n41188;
  assign n41190 = n41187 | n41188;
  assign n41191 = ~n41189 & n41190;
  assign n61374 = n40820 | n40822;
  assign n61391 = n41191 & n61374;
  assign n61392 = n40820 & n41191;
  assign n61393 = (n72855 & n61391) | (n72855 & n61392) | (n61391 & n61392);
  assign n61394 = n41191 | n61374;
  assign n61395 = n40820 | n41191;
  assign n61396 = (n72855 & n61394) | (n72855 & n61395) | (n61394 & n61395);
  assign n41194 = ~n61393 & n61396;
  assign n41195 = x172 & x197;
  assign n41196 = n41194 & n41195;
  assign n41197 = n41194 | n41195;
  assign n41198 = ~n41196 & n41197;
  assign n61397 = n40827 & n41198;
  assign n72931 = (n41198 & n61186) | (n41198 & n61397) | (n61186 & n61397);
  assign n72932 = (n41198 & n61185) | (n41198 & n61397) | (n61185 & n61397);
  assign n72933 = (n60940 & n72931) | (n60940 & n72932) | (n72931 & n72932);
  assign n61399 = n40827 | n41198;
  assign n72934 = n61186 | n61399;
  assign n72935 = n61185 | n61399;
  assign n72936 = (n60940 & n72934) | (n60940 & n72935) | (n72934 & n72935);
  assign n41201 = ~n72933 & n72936;
  assign n41202 = x171 & x198;
  assign n41203 = n41201 & n41202;
  assign n41204 = n41201 | n41202;
  assign n41205 = ~n41203 & n41204;
  assign n61372 = n40834 | n40836;
  assign n72937 = n41205 & n61372;
  assign n72911 = n40457 | n40834;
  assign n72912 = (n40834 & n40836) | (n40834 & n72911) | (n40836 & n72911);
  assign n72938 = n41205 & n72912;
  assign n72939 = (n60978 & n72937) | (n60978 & n72938) | (n72937 & n72938);
  assign n72940 = n41205 | n61372;
  assign n72941 = n41205 | n72912;
  assign n72942 = (n60978 & n72940) | (n60978 & n72941) | (n72940 & n72941);
  assign n41208 = ~n72939 & n72942;
  assign n41209 = x170 & x199;
  assign n41210 = n41208 & n41209;
  assign n41211 = n41208 | n41209;
  assign n41212 = ~n41210 & n41211;
  assign n61369 = n40841 | n40843;
  assign n61401 = n41212 & n61369;
  assign n61402 = n40841 & n41212;
  assign n61403 = (n72850 & n61401) | (n72850 & n61402) | (n61401 & n61402);
  assign n61404 = n41212 | n61369;
  assign n61405 = n40841 | n41212;
  assign n61406 = (n72850 & n61404) | (n72850 & n61405) | (n61404 & n61405);
  assign n41215 = ~n61403 & n61406;
  assign n41216 = x169 & x200;
  assign n41217 = n41215 & n41216;
  assign n41218 = n41215 | n41216;
  assign n41219 = ~n41217 & n41218;
  assign n61407 = n40848 & n41219;
  assign n72943 = (n41219 & n61196) | (n41219 & n61407) | (n61196 & n61407);
  assign n72944 = (n41219 & n61195) | (n41219 & n61407) | (n61195 & n61407);
  assign n72945 = (n60935 & n72943) | (n60935 & n72944) | (n72943 & n72944);
  assign n61409 = n40848 | n41219;
  assign n72946 = n61196 | n61409;
  assign n72947 = n61195 | n61409;
  assign n72948 = (n60935 & n72946) | (n60935 & n72947) | (n72946 & n72947);
  assign n41222 = ~n72945 & n72948;
  assign n41223 = x168 & x201;
  assign n41224 = n41222 & n41223;
  assign n41225 = n41222 | n41223;
  assign n41226 = ~n41224 & n41225;
  assign n61367 = n40855 | n40857;
  assign n72949 = n41226 & n61367;
  assign n72909 = n40478 | n40855;
  assign n72910 = (n40855 & n40857) | (n40855 & n72909) | (n40857 & n72909);
  assign n72950 = n41226 & n72910;
  assign n72951 = (n60988 & n72949) | (n60988 & n72950) | (n72949 & n72950);
  assign n72952 = n41226 | n61367;
  assign n72953 = n41226 | n72910;
  assign n72954 = (n60988 & n72952) | (n60988 & n72953) | (n72952 & n72953);
  assign n41229 = ~n72951 & n72954;
  assign n41230 = x167 & x202;
  assign n41231 = n41229 & n41230;
  assign n41232 = n41229 | n41230;
  assign n41233 = ~n41231 & n41232;
  assign n61364 = n40862 | n40864;
  assign n61411 = n41233 & n61364;
  assign n61412 = n40862 & n41233;
  assign n61413 = (n72845 & n61411) | (n72845 & n61412) | (n61411 & n61412);
  assign n61414 = n41233 | n61364;
  assign n61415 = n40862 | n41233;
  assign n61416 = (n72845 & n61414) | (n72845 & n61415) | (n61414 & n61415);
  assign n41236 = ~n61413 & n61416;
  assign n41237 = x166 & x203;
  assign n41238 = n41236 & n41237;
  assign n41239 = n41236 | n41237;
  assign n41240 = ~n41238 & n41239;
  assign n61417 = n40869 & n41240;
  assign n72955 = (n41240 & n61206) | (n41240 & n61417) | (n61206 & n61417);
  assign n72956 = (n41240 & n61205) | (n41240 & n61417) | (n61205 & n61417);
  assign n72957 = (n60930 & n72955) | (n60930 & n72956) | (n72955 & n72956);
  assign n61419 = n40869 | n41240;
  assign n72958 = n61206 | n61419;
  assign n72959 = n61205 | n61419;
  assign n72960 = (n60930 & n72958) | (n60930 & n72959) | (n72958 & n72959);
  assign n41243 = ~n72957 & n72960;
  assign n41244 = x165 & x204;
  assign n41245 = n41243 & n41244;
  assign n41246 = n41243 | n41244;
  assign n41247 = ~n41245 & n41246;
  assign n61362 = n40876 | n40878;
  assign n72961 = n41247 & n61362;
  assign n72907 = n40499 | n40876;
  assign n72908 = (n40876 & n40878) | (n40876 & n72907) | (n40878 & n72907);
  assign n72962 = n41247 & n72908;
  assign n72963 = (n60998 & n72961) | (n60998 & n72962) | (n72961 & n72962);
  assign n72964 = n41247 | n61362;
  assign n72965 = n41247 | n72908;
  assign n72966 = (n60998 & n72964) | (n60998 & n72965) | (n72964 & n72965);
  assign n41250 = ~n72963 & n72966;
  assign n41251 = x164 & x205;
  assign n41252 = n41250 & n41251;
  assign n41253 = n41250 | n41251;
  assign n41254 = ~n41252 & n41253;
  assign n61359 = n40883 | n40885;
  assign n61421 = n41254 & n61359;
  assign n61422 = n40883 & n41254;
  assign n61423 = (n72840 & n61421) | (n72840 & n61422) | (n61421 & n61422);
  assign n61424 = n41254 | n61359;
  assign n61425 = n40883 | n41254;
  assign n61426 = (n72840 & n61424) | (n72840 & n61425) | (n61424 & n61425);
  assign n41257 = ~n61423 & n61426;
  assign n41258 = x163 & x206;
  assign n41259 = n41257 & n41258;
  assign n41260 = n41257 | n41258;
  assign n41261 = ~n41259 & n41260;
  assign n61427 = n40890 & n41261;
  assign n72967 = (n41261 & n61216) | (n41261 & n61427) | (n61216 & n61427);
  assign n72968 = (n41261 & n61215) | (n41261 & n61427) | (n61215 & n61427);
  assign n72969 = (n72744 & n72967) | (n72744 & n72968) | (n72967 & n72968);
  assign n61429 = n40890 | n41261;
  assign n72970 = n61216 | n61429;
  assign n72971 = n61215 | n61429;
  assign n72972 = (n72744 & n72970) | (n72744 & n72971) | (n72970 & n72971);
  assign n41264 = ~n72969 & n72972;
  assign n41265 = x162 & x207;
  assign n41266 = n41264 & n41265;
  assign n41267 = n41264 | n41265;
  assign n41268 = ~n41266 & n41267;
  assign n41269 = n72906 & n41268;
  assign n41270 = n72906 | n41268;
  assign n41271 = ~n41269 & n41270;
  assign n41272 = x161 & x208;
  assign n41273 = n41271 & n41272;
  assign n41274 = n41271 | n41272;
  assign n41275 = ~n41273 & n41274;
  assign n61354 = n40904 | n40906;
  assign n61431 = n41275 & n61354;
  assign n61432 = n40904 & n41275;
  assign n61433 = (n72835 & n61431) | (n72835 & n61432) | (n61431 & n61432);
  assign n61434 = n41275 | n61354;
  assign n61435 = n40904 | n41275;
  assign n61436 = (n72835 & n61434) | (n72835 & n61435) | (n61434 & n61435);
  assign n41278 = ~n61433 & n61436;
  assign n41279 = x160 & x209;
  assign n41280 = n41278 & n41279;
  assign n41281 = n41278 | n41279;
  assign n41282 = ~n41280 & n41281;
  assign n61437 = n40911 & n41282;
  assign n72973 = (n41282 & n61226) | (n41282 & n61437) | (n61226 & n61437);
  assign n72974 = (n41282 & n61225) | (n41282 & n61437) | (n61225 & n61437);
  assign n72975 = (n72739 & n72973) | (n72739 & n72974) | (n72973 & n72974);
  assign n61439 = n40911 | n41282;
  assign n72976 = n61226 | n61439;
  assign n72977 = n61225 | n61439;
  assign n72978 = (n72739 & n72976) | (n72739 & n72977) | (n72976 & n72977);
  assign n41285 = ~n72975 & n72978;
  assign n41286 = x159 & x210;
  assign n41287 = n41285 & n41286;
  assign n41288 = n41285 | n41286;
  assign n41289 = ~n41287 & n41288;
  assign n41290 = n72901 & n41289;
  assign n41291 = n72901 | n41289;
  assign n41292 = ~n41290 & n41291;
  assign n41293 = x158 & x211;
  assign n41294 = n41292 & n41293;
  assign n41295 = n41292 | n41293;
  assign n41296 = ~n41294 & n41295;
  assign n61349 = n40925 | n40927;
  assign n61441 = n41296 & n61349;
  assign n61442 = n40925 & n41296;
  assign n61443 = (n61140 & n61441) | (n61140 & n61442) | (n61441 & n61442);
  assign n61444 = n41296 | n61349;
  assign n61445 = n40925 | n41296;
  assign n61446 = (n61140 & n61444) | (n61140 & n61445) | (n61444 & n61445);
  assign n41299 = ~n61443 & n61446;
  assign n41300 = x157 & x212;
  assign n41301 = n41299 & n41300;
  assign n41302 = n41299 | n41300;
  assign n41303 = ~n41301 & n41302;
  assign n61447 = n40932 & n41303;
  assign n61448 = (n41303 & n72893) | (n41303 & n61447) | (n72893 & n61447);
  assign n61449 = n40932 | n41303;
  assign n61450 = n72893 | n61449;
  assign n41306 = ~n61448 & n61450;
  assign n41307 = x156 & x213;
  assign n41308 = n41306 & n41307;
  assign n41309 = n41306 | n41307;
  assign n41310 = ~n41308 & n41309;
  assign n61451 = n40939 & n41310;
  assign n61452 = (n41310 & n61240) | (n41310 & n61451) | (n61240 & n61451);
  assign n61453 = n40939 | n41310;
  assign n61454 = n61240 | n61453;
  assign n41313 = ~n61452 & n61454;
  assign n41314 = x155 & x214;
  assign n41315 = n41313 & n41314;
  assign n41316 = n41313 | n41314;
  assign n41317 = ~n41315 & n41316;
  assign n61455 = n40946 & n41317;
  assign n61456 = (n41317 & n61244) | (n41317 & n61455) | (n61244 & n61455);
  assign n61457 = n40946 | n41317;
  assign n61458 = n61244 | n61457;
  assign n41320 = ~n61456 & n61458;
  assign n41321 = x154 & x215;
  assign n41322 = n41320 & n41321;
  assign n41323 = n41320 | n41321;
  assign n41324 = ~n41322 & n41323;
  assign n61459 = n40953 & n41324;
  assign n61460 = (n41324 & n61248) | (n41324 & n61459) | (n61248 & n61459);
  assign n61461 = n40953 | n41324;
  assign n61462 = n61248 | n61461;
  assign n41327 = ~n61460 & n61462;
  assign n41328 = x153 & x216;
  assign n41329 = n41327 & n41328;
  assign n41330 = n41327 | n41328;
  assign n41331 = ~n41329 & n41330;
  assign n61463 = n40960 & n41331;
  assign n61464 = (n41331 & n61252) | (n41331 & n61463) | (n61252 & n61463);
  assign n61465 = n40960 | n41331;
  assign n61466 = n61252 | n61465;
  assign n41334 = ~n61464 & n61466;
  assign n41335 = x152 & x217;
  assign n41336 = n41334 & n41335;
  assign n41337 = n41334 | n41335;
  assign n41338 = ~n41336 & n41337;
  assign n61467 = n40967 & n41338;
  assign n61468 = (n41338 & n61256) | (n41338 & n61467) | (n61256 & n61467);
  assign n61469 = n40967 | n41338;
  assign n61470 = n61256 | n61469;
  assign n41341 = ~n61468 & n61470;
  assign n41342 = x151 & x218;
  assign n41343 = n41341 & n41342;
  assign n41344 = n41341 | n41342;
  assign n41345 = ~n41343 & n41344;
  assign n61471 = n40974 & n41345;
  assign n61472 = (n41345 & n61260) | (n41345 & n61471) | (n61260 & n61471);
  assign n61473 = n40974 | n41345;
  assign n61474 = n61260 | n61473;
  assign n41348 = ~n61472 & n61474;
  assign n41349 = x150 & x219;
  assign n41350 = n41348 & n41349;
  assign n41351 = n41348 | n41349;
  assign n41352 = ~n41350 & n41351;
  assign n61475 = n40981 & n41352;
  assign n61476 = (n41352 & n61264) | (n41352 & n61475) | (n61264 & n61475);
  assign n61477 = n40981 | n41352;
  assign n61478 = n61264 | n61477;
  assign n41355 = ~n61476 & n61478;
  assign n41356 = x149 & x220;
  assign n41357 = n41355 & n41356;
  assign n41358 = n41355 | n41356;
  assign n41359 = ~n41357 & n41358;
  assign n61479 = n40988 & n41359;
  assign n61480 = (n41359 & n61268) | (n41359 & n61479) | (n61268 & n61479);
  assign n61481 = n40988 | n41359;
  assign n61482 = n61268 | n61481;
  assign n41362 = ~n61480 & n61482;
  assign n41363 = x148 & x221;
  assign n41364 = n41362 & n41363;
  assign n41365 = n41362 | n41363;
  assign n41366 = ~n41364 & n41365;
  assign n61483 = n40995 & n41366;
  assign n61484 = (n41366 & n61272) | (n41366 & n61483) | (n61272 & n61483);
  assign n61485 = n40995 | n41366;
  assign n61486 = n61272 | n61485;
  assign n41369 = ~n61484 & n61486;
  assign n41370 = x147 & x222;
  assign n41371 = n41369 & n41370;
  assign n41372 = n41369 | n41370;
  assign n41373 = ~n41371 & n41372;
  assign n61487 = n41002 & n41373;
  assign n61488 = (n41373 & n61276) | (n41373 & n61487) | (n61276 & n61487);
  assign n61489 = n41002 | n41373;
  assign n61490 = n61276 | n61489;
  assign n41376 = ~n61488 & n61490;
  assign n41377 = x146 & x223;
  assign n41378 = n41376 & n41377;
  assign n41379 = n41376 | n41377;
  assign n41380 = ~n41378 & n41379;
  assign n61491 = n41009 & n41380;
  assign n61492 = (n41380 & n61280) | (n41380 & n61491) | (n61280 & n61491);
  assign n61493 = n41009 | n41380;
  assign n61494 = n61280 | n61493;
  assign n41383 = ~n61492 & n61494;
  assign n41384 = x145 & x224;
  assign n41385 = n41383 & n41384;
  assign n41386 = n41383 | n41384;
  assign n41387 = ~n41385 & n41386;
  assign n61495 = n41016 & n41387;
  assign n61496 = (n41387 & n61284) | (n41387 & n61495) | (n61284 & n61495);
  assign n61497 = n41016 | n41387;
  assign n61498 = n61284 | n61497;
  assign n41390 = ~n61496 & n61498;
  assign n41391 = x144 & x225;
  assign n41392 = n41390 & n41391;
  assign n41393 = n41390 | n41391;
  assign n41394 = ~n41392 & n41393;
  assign n61499 = n41023 & n41394;
  assign n61500 = (n41394 & n61288) | (n41394 & n61499) | (n61288 & n61499);
  assign n61501 = n41023 | n41394;
  assign n61502 = n61288 | n61501;
  assign n41397 = ~n61500 & n61502;
  assign n41398 = x143 & x226;
  assign n41399 = n41397 & n41398;
  assign n41400 = n41397 | n41398;
  assign n41401 = ~n41399 & n41400;
  assign n61503 = n41030 & n41401;
  assign n61504 = (n41401 & n61292) | (n41401 & n61503) | (n61292 & n61503);
  assign n61505 = n41030 | n41401;
  assign n61506 = n61292 | n61505;
  assign n41404 = ~n61504 & n61506;
  assign n41405 = x142 & x227;
  assign n41406 = n41404 & n41405;
  assign n41407 = n41404 | n41405;
  assign n41408 = ~n41406 & n41407;
  assign n61507 = n41037 & n41408;
  assign n61508 = (n41408 & n61296) | (n41408 & n61507) | (n61296 & n61507);
  assign n61509 = n41037 | n41408;
  assign n61510 = n61296 | n61509;
  assign n41411 = ~n61508 & n61510;
  assign n41412 = x141 & x228;
  assign n41413 = n41411 & n41412;
  assign n41414 = n41411 | n41412;
  assign n41415 = ~n41413 & n41414;
  assign n61511 = n41044 & n41415;
  assign n61512 = (n41415 & n61300) | (n41415 & n61511) | (n61300 & n61511);
  assign n61513 = n41044 | n41415;
  assign n61514 = n61300 | n61513;
  assign n41418 = ~n61512 & n61514;
  assign n41419 = x140 & x229;
  assign n41420 = n41418 & n41419;
  assign n41421 = n41418 | n41419;
  assign n41422 = ~n41420 & n41421;
  assign n61515 = n41051 & n41422;
  assign n61516 = (n41422 & n61304) | (n41422 & n61515) | (n61304 & n61515);
  assign n61517 = n41051 | n41422;
  assign n61518 = n61304 | n61517;
  assign n41425 = ~n61516 & n61518;
  assign n41426 = x139 & x230;
  assign n41427 = n41425 & n41426;
  assign n41428 = n41425 | n41426;
  assign n41429 = ~n41427 & n41428;
  assign n61519 = n41058 & n41429;
  assign n61520 = (n41429 & n61308) | (n41429 & n61519) | (n61308 & n61519);
  assign n61521 = n41058 | n41429;
  assign n61522 = n61308 | n61521;
  assign n41432 = ~n61520 & n61522;
  assign n41433 = x138 & x231;
  assign n41434 = n41432 & n41433;
  assign n41435 = n41432 | n41433;
  assign n41436 = ~n41434 & n41435;
  assign n61523 = n41065 & n41436;
  assign n61524 = (n41436 & n61312) | (n41436 & n61523) | (n61312 & n61523);
  assign n61525 = n41065 | n41436;
  assign n61526 = n61312 | n61525;
  assign n41439 = ~n61524 & n61526;
  assign n41440 = x137 & x232;
  assign n41441 = n41439 & n41440;
  assign n41442 = n41439 | n41440;
  assign n41443 = ~n41441 & n41442;
  assign n61527 = n41072 & n41443;
  assign n61528 = (n41443 & n61316) | (n41443 & n61527) | (n61316 & n61527);
  assign n61529 = n41072 | n41443;
  assign n61530 = n61316 | n61529;
  assign n41446 = ~n61528 & n61530;
  assign n41447 = x136 & x233;
  assign n41448 = n41446 & n41447;
  assign n41449 = n41446 | n41447;
  assign n41450 = ~n41448 & n41449;
  assign n61531 = n41079 & n41450;
  assign n61532 = (n41450 & n61320) | (n41450 & n61531) | (n61320 & n61531);
  assign n61533 = n41079 | n41450;
  assign n61534 = n61320 | n61533;
  assign n41453 = ~n61532 & n61534;
  assign n41454 = x135 & x234;
  assign n41455 = n41453 & n41454;
  assign n41456 = n41453 | n41454;
  assign n41457 = ~n41455 & n41456;
  assign n61535 = n41086 & n41457;
  assign n61536 = (n41457 & n61324) | (n41457 & n61535) | (n61324 & n61535);
  assign n61537 = n41086 | n41457;
  assign n61538 = n61324 | n61537;
  assign n41460 = ~n61536 & n61538;
  assign n41461 = x134 & x235;
  assign n41462 = n41460 & n41461;
  assign n41463 = n41460 | n41461;
  assign n41464 = ~n41462 & n41463;
  assign n61539 = n41093 & n41464;
  assign n61540 = (n41464 & n61328) | (n41464 & n61539) | (n61328 & n61539);
  assign n61541 = n41093 | n41464;
  assign n61542 = n61328 | n61541;
  assign n41467 = ~n61540 & n61542;
  assign n41468 = x133 & x236;
  assign n41469 = n41467 & n41468;
  assign n41470 = n41467 | n41468;
  assign n41471 = ~n41469 & n41470;
  assign n61543 = n41100 & n41471;
  assign n61544 = (n41471 & n61332) | (n41471 & n61543) | (n61332 & n61543);
  assign n61545 = n41100 | n41471;
  assign n61546 = n61332 | n61545;
  assign n41474 = ~n61544 & n61546;
  assign n41475 = x132 & x237;
  assign n41476 = n41474 & n41475;
  assign n41477 = n41474 | n41475;
  assign n41478 = ~n41476 & n41477;
  assign n61547 = n41107 & n41478;
  assign n61548 = (n41478 & n61336) | (n41478 & n61547) | (n61336 & n61547);
  assign n61549 = n41107 | n41478;
  assign n61550 = n61336 | n61549;
  assign n41481 = ~n61548 & n61550;
  assign n41482 = x131 & x238;
  assign n41483 = n41481 & n41482;
  assign n41484 = n41481 | n41482;
  assign n41485 = ~n41483 & n41484;
  assign n61551 = n41114 & n41485;
  assign n61552 = (n41485 & n61340) | (n41485 & n61551) | (n61340 & n61551);
  assign n61553 = n41114 | n41485;
  assign n61554 = n61340 | n61553;
  assign n41488 = ~n61552 & n61554;
  assign n41489 = x130 & x239;
  assign n41490 = n41488 & n41489;
  assign n41491 = n41488 | n41489;
  assign n41492 = ~n41490 & n41491;
  assign n61555 = n41121 & n41492;
  assign n61556 = (n41492 & n61345) | (n41492 & n61555) | (n61345 & n61555);
  assign n61557 = n41121 | n41492;
  assign n61558 = n61345 | n61557;
  assign n41495 = ~n61556 & n61558;
  assign n61565 = n41280 | n41282;
  assign n72981 = n40911 | n41280;
  assign n72982 = (n41280 & n41282) | (n41280 & n72981) | (n41282 & n72981);
  assign n72983 = (n61226 & n61565) | (n61226 & n72982) | (n61565 & n72982);
  assign n72984 = (n61225 & n61565) | (n61225 & n72982) | (n61565 & n72982);
  assign n72985 = (n72739 & n72983) | (n72739 & n72984) | (n72983 & n72984);
  assign n61570 = n41259 | n41261;
  assign n72986 = n40890 | n41259;
  assign n72987 = (n41259 & n41261) | (n41259 & n72986) | (n41261 & n72986);
  assign n72988 = (n61216 & n61570) | (n61216 & n72987) | (n61570 & n72987);
  assign n72989 = (n61215 & n61570) | (n61215 & n72987) | (n61570 & n72987);
  assign n72990 = (n72744 & n72988) | (n72744 & n72989) | (n72988 & n72989);
  assign n61363 = (n60998 & n72908) | (n60998 & n61362) | (n72908 & n61362);
  assign n61575 = n41238 | n41240;
  assign n72991 = n40869 | n41238;
  assign n72992 = (n41238 & n41240) | (n41238 & n72991) | (n41240 & n72991);
  assign n72993 = (n61206 & n61575) | (n61206 & n72992) | (n61575 & n72992);
  assign n72994 = (n61205 & n61575) | (n61205 & n72992) | (n61575 & n72992);
  assign n72995 = (n60930 & n72993) | (n60930 & n72994) | (n72993 & n72994);
  assign n61368 = (n60988 & n72910) | (n60988 & n61367) | (n72910 & n61367);
  assign n61580 = n41217 | n41219;
  assign n72996 = n40848 | n41217;
  assign n72997 = (n41217 & n41219) | (n41217 & n72996) | (n41219 & n72996);
  assign n72998 = (n61196 & n61580) | (n61196 & n72997) | (n61580 & n72997);
  assign n72999 = (n61195 & n61580) | (n61195 & n72997) | (n61580 & n72997);
  assign n73000 = (n60935 & n72998) | (n60935 & n72999) | (n72998 & n72999);
  assign n61373 = (n60978 & n72912) | (n60978 & n61372) | (n72912 & n61372);
  assign n61585 = n41196 | n41198;
  assign n73001 = n40827 | n41196;
  assign n73002 = (n41196 & n41198) | (n41196 & n73001) | (n41198 & n73001);
  assign n73003 = (n61186 & n61585) | (n61186 & n73002) | (n61585 & n73002);
  assign n73004 = (n61185 & n61585) | (n61185 & n73002) | (n61585 & n73002);
  assign n73005 = (n60940 & n73003) | (n60940 & n73004) | (n73003 & n73004);
  assign n41542 = x175 & x195;
  assign n61590 = n41177 | n61383;
  assign n73006 = (n40806 & n61383) | (n40806 & n61590) | (n61383 & n61590);
  assign n61592 = n41542 & n73006;
  assign n73007 = n41542 & n61383;
  assign n73008 = (n41177 & n41542) | (n41177 & n73007) | (n41542 & n73007);
  assign n73009 = (n61176 & n61592) | (n61176 & n73008) | (n61592 & n73008);
  assign n73010 = (n61175 & n61592) | (n61175 & n73008) | (n61592 & n73008);
  assign n73011 = (n60945 & n73009) | (n60945 & n73010) | (n73009 & n73010);
  assign n61595 = n41542 | n73006;
  assign n73012 = n41542 | n61383;
  assign n73013 = n41177 | n73012;
  assign n73014 = (n61176 & n61595) | (n61176 & n73013) | (n61595 & n73013);
  assign n73015 = (n61175 & n61595) | (n61175 & n73013) | (n61595 & n73013);
  assign n73016 = (n60945 & n73014) | (n60945 & n73015) | (n73014 & n73015);
  assign n41545 = ~n73011 & n73016;
  assign n61599 = n41182 & n41545;
  assign n73017 = (n41184 & n41545) | (n41184 & n61599) | (n41545 & n61599);
  assign n73018 = (n61377 & n61599) | (n61377 & n73017) | (n61599 & n73017);
  assign n73019 = (n61599 & n72914) | (n61599 & n73017) | (n72914 & n73017);
  assign n73020 = (n60968 & n73018) | (n60968 & n73019) | (n73018 & n73019);
  assign n61602 = n41182 | n41545;
  assign n73021 = n41184 | n61602;
  assign n73022 = (n61377 & n61602) | (n61377 & n73021) | (n61602 & n73021);
  assign n73023 = (n61602 & n72914) | (n61602 & n73021) | (n72914 & n73021);
  assign n73024 = (n60968 & n73022) | (n60968 & n73023) | (n73022 & n73023);
  assign n41548 = ~n73020 & n73024;
  assign n41549 = x174 & x196;
  assign n41550 = n41548 & n41549;
  assign n41551 = n41548 | n41549;
  assign n41552 = ~n41550 & n41551;
  assign n61604 = n41189 & n41552;
  assign n61605 = (n41552 & n61393) | (n41552 & n61604) | (n61393 & n61604);
  assign n61606 = n41189 | n41552;
  assign n61607 = n61393 | n61606;
  assign n41555 = ~n61605 & n61607;
  assign n41556 = x173 & x197;
  assign n41557 = n41555 & n41556;
  assign n41558 = n41555 | n41556;
  assign n41559 = ~n41557 & n41558;
  assign n41560 = n73005 & n41559;
  assign n41561 = n73005 | n41559;
  assign n41562 = ~n41560 & n41561;
  assign n41563 = x172 & x198;
  assign n41564 = n41562 & n41563;
  assign n41565 = n41562 | n41563;
  assign n41566 = ~n41564 & n41565;
  assign n61582 = n41203 | n41205;
  assign n61608 = n41566 & n61582;
  assign n61609 = n41203 & n41566;
  assign n61610 = (n61373 & n61608) | (n61373 & n61609) | (n61608 & n61609);
  assign n61611 = n41566 | n61582;
  assign n61612 = n41203 | n41566;
  assign n61613 = (n61373 & n61611) | (n61373 & n61612) | (n61611 & n61612);
  assign n41569 = ~n61610 & n61613;
  assign n41570 = x171 & x199;
  assign n41571 = n41569 & n41570;
  assign n41572 = n41569 | n41570;
  assign n41573 = ~n41571 & n41572;
  assign n61614 = n41210 & n41573;
  assign n61615 = (n41573 & n61403) | (n41573 & n61614) | (n61403 & n61614);
  assign n61616 = n41210 | n41573;
  assign n61617 = n61403 | n61616;
  assign n41576 = ~n61615 & n61617;
  assign n41577 = x170 & x200;
  assign n41578 = n41576 & n41577;
  assign n41579 = n41576 | n41577;
  assign n41580 = ~n41578 & n41579;
  assign n41581 = n73000 & n41580;
  assign n41582 = n73000 | n41580;
  assign n41583 = ~n41581 & n41582;
  assign n41584 = x169 & x201;
  assign n41585 = n41583 & n41584;
  assign n41586 = n41583 | n41584;
  assign n41587 = ~n41585 & n41586;
  assign n61577 = n41224 | n41226;
  assign n61618 = n41587 & n61577;
  assign n61619 = n41224 & n41587;
  assign n61620 = (n61368 & n61618) | (n61368 & n61619) | (n61618 & n61619);
  assign n61621 = n41587 | n61577;
  assign n61622 = n41224 | n41587;
  assign n61623 = (n61368 & n61621) | (n61368 & n61622) | (n61621 & n61622);
  assign n41590 = ~n61620 & n61623;
  assign n41591 = x168 & x202;
  assign n41592 = n41590 & n41591;
  assign n41593 = n41590 | n41591;
  assign n41594 = ~n41592 & n41593;
  assign n61624 = n41231 & n41594;
  assign n61625 = (n41594 & n61413) | (n41594 & n61624) | (n61413 & n61624);
  assign n61626 = n41231 | n41594;
  assign n61627 = n61413 | n61626;
  assign n41597 = ~n61625 & n61627;
  assign n41598 = x167 & x203;
  assign n41599 = n41597 & n41598;
  assign n41600 = n41597 | n41598;
  assign n41601 = ~n41599 & n41600;
  assign n41602 = n72995 & n41601;
  assign n41603 = n72995 | n41601;
  assign n41604 = ~n41602 & n41603;
  assign n41605 = x166 & x204;
  assign n41606 = n41604 & n41605;
  assign n41607 = n41604 | n41605;
  assign n41608 = ~n41606 & n41607;
  assign n61572 = n41245 | n41247;
  assign n61628 = n41608 & n61572;
  assign n61629 = n41245 & n41608;
  assign n61630 = (n61363 & n61628) | (n61363 & n61629) | (n61628 & n61629);
  assign n61631 = n41608 | n61572;
  assign n61632 = n41245 | n41608;
  assign n61633 = (n61363 & n61631) | (n61363 & n61632) | (n61631 & n61632);
  assign n41611 = ~n61630 & n61633;
  assign n41612 = x165 & x205;
  assign n41613 = n41611 & n41612;
  assign n41614 = n41611 | n41612;
  assign n41615 = ~n41613 & n41614;
  assign n61634 = n41252 & n41615;
  assign n61635 = (n41615 & n61423) | (n41615 & n61634) | (n61423 & n61634);
  assign n61636 = n41252 | n41615;
  assign n61637 = n61423 | n61636;
  assign n41618 = ~n61635 & n61637;
  assign n41619 = x164 & x206;
  assign n41620 = n41618 & n41619;
  assign n41621 = n41618 | n41619;
  assign n41622 = ~n41620 & n41621;
  assign n41623 = n72990 & n41622;
  assign n41624 = n72990 | n41622;
  assign n41625 = ~n41623 & n41624;
  assign n41626 = x163 & x207;
  assign n41627 = n41625 & n41626;
  assign n41628 = n41625 | n41626;
  assign n41629 = ~n41627 & n41628;
  assign n61567 = n41266 | n41268;
  assign n61638 = n41629 & n61567;
  assign n61639 = n41266 & n41629;
  assign n61640 = (n72906 & n61638) | (n72906 & n61639) | (n61638 & n61639);
  assign n61641 = n41629 | n61567;
  assign n61642 = n41266 | n41629;
  assign n61643 = (n72906 & n61641) | (n72906 & n61642) | (n61641 & n61642);
  assign n41632 = ~n61640 & n61643;
  assign n41633 = x162 & x208;
  assign n41634 = n41632 & n41633;
  assign n41635 = n41632 | n41633;
  assign n41636 = ~n41634 & n41635;
  assign n61644 = n41273 & n41636;
  assign n73025 = (n41636 & n61432) | (n41636 & n61644) | (n61432 & n61644);
  assign n73026 = (n41636 & n61431) | (n41636 & n61644) | (n61431 & n61644);
  assign n73027 = (n72835 & n73025) | (n72835 & n73026) | (n73025 & n73026);
  assign n61646 = n41273 | n41636;
  assign n73028 = n61432 | n61646;
  assign n73029 = n61431 | n61646;
  assign n73030 = (n72835 & n73028) | (n72835 & n73029) | (n73028 & n73029);
  assign n41639 = ~n73027 & n73030;
  assign n41640 = x161 & x209;
  assign n41641 = n41639 & n41640;
  assign n41642 = n41639 | n41640;
  assign n41643 = ~n41641 & n41642;
  assign n41644 = n72985 & n41643;
  assign n41645 = n72985 | n41643;
  assign n41646 = ~n41644 & n41645;
  assign n41647 = x160 & x210;
  assign n41648 = n41646 & n41647;
  assign n41649 = n41646 | n41647;
  assign n41650 = ~n41648 & n41649;
  assign n61562 = n41287 | n41289;
  assign n61648 = n41650 & n61562;
  assign n61649 = n41287 & n41650;
  assign n61650 = (n72901 & n61648) | (n72901 & n61649) | (n61648 & n61649);
  assign n61651 = n41650 | n61562;
  assign n61652 = n41287 | n41650;
  assign n61653 = (n72901 & n61651) | (n72901 & n61652) | (n61651 & n61652);
  assign n41653 = ~n61650 & n61653;
  assign n41654 = x159 & x211;
  assign n41655 = n41653 & n41654;
  assign n41656 = n41653 | n41654;
  assign n41657 = ~n41655 & n41656;
  assign n61654 = n41294 & n41657;
  assign n73031 = (n41657 & n61442) | (n41657 & n61654) | (n61442 & n61654);
  assign n73032 = (n41657 & n61441) | (n41657 & n61654) | (n61441 & n61654);
  assign n73033 = (n61140 & n73031) | (n61140 & n73032) | (n73031 & n73032);
  assign n61656 = n41294 | n41657;
  assign n73034 = n61442 | n61656;
  assign n73035 = n61441 | n61656;
  assign n73036 = (n61140 & n73034) | (n61140 & n73035) | (n73034 & n73035);
  assign n41660 = ~n73033 & n73036;
  assign n41661 = x158 & x212;
  assign n41662 = n41660 & n41661;
  assign n41663 = n41660 | n41661;
  assign n41664 = ~n41662 & n41663;
  assign n61560 = n41301 | n41303;
  assign n73037 = n41664 & n61560;
  assign n72979 = n40932 | n41301;
  assign n72980 = (n41301 & n41303) | (n41301 & n72979) | (n41303 & n72979);
  assign n73038 = n41664 & n72980;
  assign n73039 = (n72893 & n73037) | (n72893 & n73038) | (n73037 & n73038);
  assign n73040 = n41664 | n61560;
  assign n73041 = n41664 | n72980;
  assign n73042 = (n72893 & n73040) | (n72893 & n73041) | (n73040 & n73041);
  assign n41667 = ~n73039 & n73042;
  assign n41668 = x157 & x213;
  assign n41669 = n41667 & n41668;
  assign n41670 = n41667 | n41668;
  assign n41671 = ~n41669 & n41670;
  assign n61658 = n41308 & n41671;
  assign n73043 = (n41671 & n61451) | (n41671 & n61658) | (n61451 & n61658);
  assign n73044 = (n41310 & n41671) | (n41310 & n61658) | (n41671 & n61658);
  assign n73045 = (n61240 & n73043) | (n61240 & n73044) | (n73043 & n73044);
  assign n61660 = n41308 | n41671;
  assign n73046 = n61451 | n61660;
  assign n73047 = n41310 | n61660;
  assign n73048 = (n61240 & n73046) | (n61240 & n73047) | (n73046 & n73047);
  assign n41674 = ~n73045 & n73048;
  assign n41675 = x156 & x214;
  assign n41676 = n41674 & n41675;
  assign n41677 = n41674 | n41675;
  assign n41678 = ~n41676 & n41677;
  assign n61662 = n41315 & n41678;
  assign n61663 = (n41678 & n61456) | (n41678 & n61662) | (n61456 & n61662);
  assign n61664 = n41315 | n41678;
  assign n61665 = n61456 | n61664;
  assign n41681 = ~n61663 & n61665;
  assign n41682 = x155 & x215;
  assign n41683 = n41681 & n41682;
  assign n41684 = n41681 | n41682;
  assign n41685 = ~n41683 & n41684;
  assign n61666 = n41322 & n41685;
  assign n61667 = (n41685 & n61460) | (n41685 & n61666) | (n61460 & n61666);
  assign n61668 = n41322 | n41685;
  assign n61669 = n61460 | n61668;
  assign n41688 = ~n61667 & n61669;
  assign n41689 = x154 & x216;
  assign n41690 = n41688 & n41689;
  assign n41691 = n41688 | n41689;
  assign n41692 = ~n41690 & n41691;
  assign n61670 = n41329 & n41692;
  assign n61671 = (n41692 & n61464) | (n41692 & n61670) | (n61464 & n61670);
  assign n61672 = n41329 | n41692;
  assign n61673 = n61464 | n61672;
  assign n41695 = ~n61671 & n61673;
  assign n41696 = x153 & x217;
  assign n41697 = n41695 & n41696;
  assign n41698 = n41695 | n41696;
  assign n41699 = ~n41697 & n41698;
  assign n61674 = n41336 & n41699;
  assign n61675 = (n41699 & n61468) | (n41699 & n61674) | (n61468 & n61674);
  assign n61676 = n41336 | n41699;
  assign n61677 = n61468 | n61676;
  assign n41702 = ~n61675 & n61677;
  assign n41703 = x152 & x218;
  assign n41704 = n41702 & n41703;
  assign n41705 = n41702 | n41703;
  assign n41706 = ~n41704 & n41705;
  assign n61678 = n41343 & n41706;
  assign n61679 = (n41706 & n61472) | (n41706 & n61678) | (n61472 & n61678);
  assign n61680 = n41343 | n41706;
  assign n61681 = n61472 | n61680;
  assign n41709 = ~n61679 & n61681;
  assign n41710 = x151 & x219;
  assign n41711 = n41709 & n41710;
  assign n41712 = n41709 | n41710;
  assign n41713 = ~n41711 & n41712;
  assign n61682 = n41350 & n41713;
  assign n61683 = (n41713 & n61476) | (n41713 & n61682) | (n61476 & n61682);
  assign n61684 = n41350 | n41713;
  assign n61685 = n61476 | n61684;
  assign n41716 = ~n61683 & n61685;
  assign n41717 = x150 & x220;
  assign n41718 = n41716 & n41717;
  assign n41719 = n41716 | n41717;
  assign n41720 = ~n41718 & n41719;
  assign n61686 = n41357 & n41720;
  assign n61687 = (n41720 & n61480) | (n41720 & n61686) | (n61480 & n61686);
  assign n61688 = n41357 | n41720;
  assign n61689 = n61480 | n61688;
  assign n41723 = ~n61687 & n61689;
  assign n41724 = x149 & x221;
  assign n41725 = n41723 & n41724;
  assign n41726 = n41723 | n41724;
  assign n41727 = ~n41725 & n41726;
  assign n61690 = n41364 & n41727;
  assign n61691 = (n41727 & n61484) | (n41727 & n61690) | (n61484 & n61690);
  assign n61692 = n41364 | n41727;
  assign n61693 = n61484 | n61692;
  assign n41730 = ~n61691 & n61693;
  assign n41731 = x148 & x222;
  assign n41732 = n41730 & n41731;
  assign n41733 = n41730 | n41731;
  assign n41734 = ~n41732 & n41733;
  assign n61694 = n41371 & n41734;
  assign n61695 = (n41734 & n61488) | (n41734 & n61694) | (n61488 & n61694);
  assign n61696 = n41371 | n41734;
  assign n61697 = n61488 | n61696;
  assign n41737 = ~n61695 & n61697;
  assign n41738 = x147 & x223;
  assign n41739 = n41737 & n41738;
  assign n41740 = n41737 | n41738;
  assign n41741 = ~n41739 & n41740;
  assign n61698 = n41378 & n41741;
  assign n61699 = (n41741 & n61492) | (n41741 & n61698) | (n61492 & n61698);
  assign n61700 = n41378 | n41741;
  assign n61701 = n61492 | n61700;
  assign n41744 = ~n61699 & n61701;
  assign n41745 = x146 & x224;
  assign n41746 = n41744 & n41745;
  assign n41747 = n41744 | n41745;
  assign n41748 = ~n41746 & n41747;
  assign n61702 = n41385 & n41748;
  assign n61703 = (n41748 & n61496) | (n41748 & n61702) | (n61496 & n61702);
  assign n61704 = n41385 | n41748;
  assign n61705 = n61496 | n61704;
  assign n41751 = ~n61703 & n61705;
  assign n41752 = x145 & x225;
  assign n41753 = n41751 & n41752;
  assign n41754 = n41751 | n41752;
  assign n41755 = ~n41753 & n41754;
  assign n61706 = n41392 & n41755;
  assign n61707 = (n41755 & n61500) | (n41755 & n61706) | (n61500 & n61706);
  assign n61708 = n41392 | n41755;
  assign n61709 = n61500 | n61708;
  assign n41758 = ~n61707 & n61709;
  assign n41759 = x144 & x226;
  assign n41760 = n41758 & n41759;
  assign n41761 = n41758 | n41759;
  assign n41762 = ~n41760 & n41761;
  assign n61710 = n41399 & n41762;
  assign n61711 = (n41762 & n61504) | (n41762 & n61710) | (n61504 & n61710);
  assign n61712 = n41399 | n41762;
  assign n61713 = n61504 | n61712;
  assign n41765 = ~n61711 & n61713;
  assign n41766 = x143 & x227;
  assign n41767 = n41765 & n41766;
  assign n41768 = n41765 | n41766;
  assign n41769 = ~n41767 & n41768;
  assign n61714 = n41406 & n41769;
  assign n61715 = (n41769 & n61508) | (n41769 & n61714) | (n61508 & n61714);
  assign n61716 = n41406 | n41769;
  assign n61717 = n61508 | n61716;
  assign n41772 = ~n61715 & n61717;
  assign n41773 = x142 & x228;
  assign n41774 = n41772 & n41773;
  assign n41775 = n41772 | n41773;
  assign n41776 = ~n41774 & n41775;
  assign n61718 = n41413 & n41776;
  assign n61719 = (n41776 & n61512) | (n41776 & n61718) | (n61512 & n61718);
  assign n61720 = n41413 | n41776;
  assign n61721 = n61512 | n61720;
  assign n41779 = ~n61719 & n61721;
  assign n41780 = x141 & x229;
  assign n41781 = n41779 & n41780;
  assign n41782 = n41779 | n41780;
  assign n41783 = ~n41781 & n41782;
  assign n61722 = n41420 & n41783;
  assign n61723 = (n41783 & n61516) | (n41783 & n61722) | (n61516 & n61722);
  assign n61724 = n41420 | n41783;
  assign n61725 = n61516 | n61724;
  assign n41786 = ~n61723 & n61725;
  assign n41787 = x140 & x230;
  assign n41788 = n41786 & n41787;
  assign n41789 = n41786 | n41787;
  assign n41790 = ~n41788 & n41789;
  assign n61726 = n41427 & n41790;
  assign n61727 = (n41790 & n61520) | (n41790 & n61726) | (n61520 & n61726);
  assign n61728 = n41427 | n41790;
  assign n61729 = n61520 | n61728;
  assign n41793 = ~n61727 & n61729;
  assign n41794 = x139 & x231;
  assign n41795 = n41793 & n41794;
  assign n41796 = n41793 | n41794;
  assign n41797 = ~n41795 & n41796;
  assign n61730 = n41434 & n41797;
  assign n61731 = (n41797 & n61524) | (n41797 & n61730) | (n61524 & n61730);
  assign n61732 = n41434 | n41797;
  assign n61733 = n61524 | n61732;
  assign n41800 = ~n61731 & n61733;
  assign n41801 = x138 & x232;
  assign n41802 = n41800 & n41801;
  assign n41803 = n41800 | n41801;
  assign n41804 = ~n41802 & n41803;
  assign n61734 = n41441 & n41804;
  assign n61735 = (n41804 & n61528) | (n41804 & n61734) | (n61528 & n61734);
  assign n61736 = n41441 | n41804;
  assign n61737 = n61528 | n61736;
  assign n41807 = ~n61735 & n61737;
  assign n41808 = x137 & x233;
  assign n41809 = n41807 & n41808;
  assign n41810 = n41807 | n41808;
  assign n41811 = ~n41809 & n41810;
  assign n61738 = n41448 & n41811;
  assign n61739 = (n41811 & n61532) | (n41811 & n61738) | (n61532 & n61738);
  assign n61740 = n41448 | n41811;
  assign n61741 = n61532 | n61740;
  assign n41814 = ~n61739 & n61741;
  assign n41815 = x136 & x234;
  assign n41816 = n41814 & n41815;
  assign n41817 = n41814 | n41815;
  assign n41818 = ~n41816 & n41817;
  assign n61742 = n41455 & n41818;
  assign n61743 = (n41818 & n61536) | (n41818 & n61742) | (n61536 & n61742);
  assign n61744 = n41455 | n41818;
  assign n61745 = n61536 | n61744;
  assign n41821 = ~n61743 & n61745;
  assign n41822 = x135 & x235;
  assign n41823 = n41821 & n41822;
  assign n41824 = n41821 | n41822;
  assign n41825 = ~n41823 & n41824;
  assign n61746 = n41462 & n41825;
  assign n61747 = (n41825 & n61540) | (n41825 & n61746) | (n61540 & n61746);
  assign n61748 = n41462 | n41825;
  assign n61749 = n61540 | n61748;
  assign n41828 = ~n61747 & n61749;
  assign n41829 = x134 & x236;
  assign n41830 = n41828 & n41829;
  assign n41831 = n41828 | n41829;
  assign n41832 = ~n41830 & n41831;
  assign n61750 = n41469 & n41832;
  assign n61751 = (n41832 & n61544) | (n41832 & n61750) | (n61544 & n61750);
  assign n61752 = n41469 | n41832;
  assign n61753 = n61544 | n61752;
  assign n41835 = ~n61751 & n61753;
  assign n41836 = x133 & x237;
  assign n41837 = n41835 & n41836;
  assign n41838 = n41835 | n41836;
  assign n41839 = ~n41837 & n41838;
  assign n61754 = n41476 & n41839;
  assign n61755 = (n41839 & n61548) | (n41839 & n61754) | (n61548 & n61754);
  assign n61756 = n41476 | n41839;
  assign n61757 = n61548 | n61756;
  assign n41842 = ~n61755 & n61757;
  assign n41843 = x132 & x238;
  assign n41844 = n41842 & n41843;
  assign n41845 = n41842 | n41843;
  assign n41846 = ~n41844 & n41845;
  assign n61758 = n41483 & n41846;
  assign n61759 = (n41846 & n61552) | (n41846 & n61758) | (n61552 & n61758);
  assign n61760 = n41483 | n41846;
  assign n61761 = n61552 | n61760;
  assign n41849 = ~n61759 & n61761;
  assign n41850 = x131 & x239;
  assign n41851 = n41849 & n41850;
  assign n41852 = n41849 | n41850;
  assign n41853 = ~n41851 & n41852;
  assign n61762 = n41490 & n41853;
  assign n61763 = (n41853 & n61556) | (n41853 & n61762) | (n61556 & n61762);
  assign n61764 = n41490 | n41853;
  assign n61765 = n61556 | n61764;
  assign n41856 = ~n61763 & n61765;
  assign n61561 = (n72893 & n72980) | (n72893 & n61560) | (n72980 & n61560);
  assign n61769 = n41655 | n41657;
  assign n73049 = n41294 | n41655;
  assign n73050 = (n41655 & n41657) | (n41655 & n73049) | (n41657 & n73049);
  assign n73051 = (n61442 & n61769) | (n61442 & n73050) | (n61769 & n73050);
  assign n73052 = (n61441 & n61769) | (n61441 & n73050) | (n61769 & n73050);
  assign n73053 = (n61140 & n73051) | (n61140 & n73052) | (n73051 & n73052);
  assign n61774 = n41634 | n41636;
  assign n73054 = n41273 | n41634;
  assign n73055 = (n41634 & n41636) | (n41634 & n73054) | (n41636 & n73054);
  assign n73056 = (n61432 & n61774) | (n61432 & n73055) | (n61774 & n73055);
  assign n73057 = (n61431 & n61774) | (n61431 & n73055) | (n61774 & n73055);
  assign n73058 = (n72835 & n73056) | (n72835 & n73057) | (n73056 & n73057);
  assign n41902 = x175 & x196;
  assign n61796 = n41902 & n73011;
  assign n61797 = (n41902 & n73020) | (n41902 & n61796) | (n73020 & n61796);
  assign n61798 = n41902 | n73011;
  assign n61799 = n73020 | n61798;
  assign n41905 = ~n61797 & n61799;
  assign n61794 = n41550 | n41552;
  assign n73067 = n41905 & n61794;
  assign n73065 = n41189 | n41550;
  assign n73066 = (n41550 & n41552) | (n41550 & n73065) | (n41552 & n73065);
  assign n73068 = n41905 & n73066;
  assign n73069 = (n61393 & n73067) | (n61393 & n73068) | (n73067 & n73068);
  assign n73070 = n41905 | n61794;
  assign n73071 = n41905 | n73066;
  assign n73072 = (n61393 & n73070) | (n61393 & n73071) | (n73070 & n73071);
  assign n41908 = ~n73069 & n73072;
  assign n41909 = x174 & x197;
  assign n41910 = n41908 & n41909;
  assign n41911 = n41908 | n41909;
  assign n41912 = ~n41910 & n41911;
  assign n61791 = n41557 | n41559;
  assign n61800 = n41912 & n61791;
  assign n61801 = n41557 & n41912;
  assign n61802 = (n73005 & n61800) | (n73005 & n61801) | (n61800 & n61801);
  assign n61803 = n41912 | n61791;
  assign n61804 = n41557 | n41912;
  assign n61805 = (n73005 & n61803) | (n73005 & n61804) | (n61803 & n61804);
  assign n41915 = ~n61802 & n61805;
  assign n41916 = x173 & x198;
  assign n41917 = n41915 & n41916;
  assign n41918 = n41915 | n41916;
  assign n41919 = ~n41917 & n41918;
  assign n61806 = n41564 & n41919;
  assign n73073 = (n41919 & n61609) | (n41919 & n61806) | (n61609 & n61806);
  assign n73074 = (n41919 & n61608) | (n41919 & n61806) | (n61608 & n61806);
  assign n73075 = (n61373 & n73073) | (n61373 & n73074) | (n73073 & n73074);
  assign n61808 = n41564 | n41919;
  assign n73076 = n61609 | n61808;
  assign n73077 = n61608 | n61808;
  assign n73078 = (n61373 & n73076) | (n61373 & n73077) | (n73076 & n73077);
  assign n41922 = ~n73075 & n73078;
  assign n41923 = x172 & x199;
  assign n41924 = n41922 & n41923;
  assign n41925 = n41922 | n41923;
  assign n41926 = ~n41924 & n41925;
  assign n61789 = n41571 | n41573;
  assign n73079 = n41926 & n61789;
  assign n73063 = n41210 | n41571;
  assign n73064 = (n41571 & n41573) | (n41571 & n73063) | (n41573 & n73063);
  assign n73080 = n41926 & n73064;
  assign n73081 = (n61403 & n73079) | (n61403 & n73080) | (n73079 & n73080);
  assign n73082 = n41926 | n61789;
  assign n73083 = n41926 | n73064;
  assign n73084 = (n61403 & n73082) | (n61403 & n73083) | (n73082 & n73083);
  assign n41929 = ~n73081 & n73084;
  assign n41930 = x171 & x200;
  assign n41931 = n41929 & n41930;
  assign n41932 = n41929 | n41930;
  assign n41933 = ~n41931 & n41932;
  assign n61786 = n41578 | n41580;
  assign n61810 = n41933 & n61786;
  assign n61811 = n41578 & n41933;
  assign n61812 = (n73000 & n61810) | (n73000 & n61811) | (n61810 & n61811);
  assign n61813 = n41933 | n61786;
  assign n61814 = n41578 | n41933;
  assign n61815 = (n73000 & n61813) | (n73000 & n61814) | (n61813 & n61814);
  assign n41936 = ~n61812 & n61815;
  assign n41937 = x170 & x201;
  assign n41938 = n41936 & n41937;
  assign n41939 = n41936 | n41937;
  assign n41940 = ~n41938 & n41939;
  assign n61816 = n41585 & n41940;
  assign n73085 = (n41940 & n61619) | (n41940 & n61816) | (n61619 & n61816);
  assign n73086 = (n41940 & n61618) | (n41940 & n61816) | (n61618 & n61816);
  assign n73087 = (n61368 & n73085) | (n61368 & n73086) | (n73085 & n73086);
  assign n61818 = n41585 | n41940;
  assign n73088 = n61619 | n61818;
  assign n73089 = n61618 | n61818;
  assign n73090 = (n61368 & n73088) | (n61368 & n73089) | (n73088 & n73089);
  assign n41943 = ~n73087 & n73090;
  assign n41944 = x169 & x202;
  assign n41945 = n41943 & n41944;
  assign n41946 = n41943 | n41944;
  assign n41947 = ~n41945 & n41946;
  assign n61784 = n41592 | n41594;
  assign n73091 = n41947 & n61784;
  assign n73061 = n41231 | n41592;
  assign n73062 = (n41592 & n41594) | (n41592 & n73061) | (n41594 & n73061);
  assign n73092 = n41947 & n73062;
  assign n73093 = (n61413 & n73091) | (n61413 & n73092) | (n73091 & n73092);
  assign n73094 = n41947 | n61784;
  assign n73095 = n41947 | n73062;
  assign n73096 = (n61413 & n73094) | (n61413 & n73095) | (n73094 & n73095);
  assign n41950 = ~n73093 & n73096;
  assign n41951 = x168 & x203;
  assign n41952 = n41950 & n41951;
  assign n41953 = n41950 | n41951;
  assign n41954 = ~n41952 & n41953;
  assign n61781 = n41599 | n41601;
  assign n61820 = n41954 & n61781;
  assign n61821 = n41599 & n41954;
  assign n61822 = (n72995 & n61820) | (n72995 & n61821) | (n61820 & n61821);
  assign n61823 = n41954 | n61781;
  assign n61824 = n41599 | n41954;
  assign n61825 = (n72995 & n61823) | (n72995 & n61824) | (n61823 & n61824);
  assign n41957 = ~n61822 & n61825;
  assign n41958 = x167 & x204;
  assign n41959 = n41957 & n41958;
  assign n41960 = n41957 | n41958;
  assign n41961 = ~n41959 & n41960;
  assign n61826 = n41606 & n41961;
  assign n73097 = (n41961 & n61629) | (n41961 & n61826) | (n61629 & n61826);
  assign n73098 = (n41961 & n61628) | (n41961 & n61826) | (n61628 & n61826);
  assign n73099 = (n61363 & n73097) | (n61363 & n73098) | (n73097 & n73098);
  assign n61828 = n41606 | n41961;
  assign n73100 = n61629 | n61828;
  assign n73101 = n61628 | n61828;
  assign n73102 = (n61363 & n73100) | (n61363 & n73101) | (n73100 & n73101);
  assign n41964 = ~n73099 & n73102;
  assign n41965 = x166 & x205;
  assign n41966 = n41964 & n41965;
  assign n41967 = n41964 | n41965;
  assign n41968 = ~n41966 & n41967;
  assign n61779 = n41613 | n41615;
  assign n73103 = n41968 & n61779;
  assign n73059 = n41252 | n41613;
  assign n73060 = (n41613 & n41615) | (n41613 & n73059) | (n41615 & n73059);
  assign n73104 = n41968 & n73060;
  assign n73105 = (n61423 & n73103) | (n61423 & n73104) | (n73103 & n73104);
  assign n73106 = n41968 | n61779;
  assign n73107 = n41968 | n73060;
  assign n73108 = (n61423 & n73106) | (n61423 & n73107) | (n73106 & n73107);
  assign n41971 = ~n73105 & n73108;
  assign n41972 = x165 & x206;
  assign n41973 = n41971 & n41972;
  assign n41974 = n41971 | n41972;
  assign n41975 = ~n41973 & n41974;
  assign n61776 = n41620 | n41622;
  assign n61830 = n41975 & n61776;
  assign n61831 = n41620 & n41975;
  assign n61832 = (n72990 & n61830) | (n72990 & n61831) | (n61830 & n61831);
  assign n61833 = n41975 | n61776;
  assign n61834 = n41620 | n41975;
  assign n61835 = (n72990 & n61833) | (n72990 & n61834) | (n61833 & n61834);
  assign n41978 = ~n61832 & n61835;
  assign n41979 = x164 & x207;
  assign n41980 = n41978 & n41979;
  assign n41981 = n41978 | n41979;
  assign n41982 = ~n41980 & n41981;
  assign n61836 = n41627 & n41982;
  assign n73109 = (n41982 & n61639) | (n41982 & n61836) | (n61639 & n61836);
  assign n73110 = (n41982 & n61638) | (n41982 & n61836) | (n61638 & n61836);
  assign n73111 = (n72906 & n73109) | (n72906 & n73110) | (n73109 & n73110);
  assign n61838 = n41627 | n41982;
  assign n73112 = n61639 | n61838;
  assign n73113 = n61638 | n61838;
  assign n73114 = (n72906 & n73112) | (n72906 & n73113) | (n73112 & n73113);
  assign n41985 = ~n73111 & n73114;
  assign n41986 = x163 & x208;
  assign n41987 = n41985 & n41986;
  assign n41988 = n41985 | n41986;
  assign n41989 = ~n41987 & n41988;
  assign n41990 = n73058 & n41989;
  assign n41991 = n73058 | n41989;
  assign n41992 = ~n41990 & n41991;
  assign n41993 = x162 & x209;
  assign n41994 = n41992 & n41993;
  assign n41995 = n41992 | n41993;
  assign n41996 = ~n41994 & n41995;
  assign n61771 = n41641 | n41643;
  assign n61840 = n41996 & n61771;
  assign n61841 = n41641 & n41996;
  assign n61842 = (n72985 & n61840) | (n72985 & n61841) | (n61840 & n61841);
  assign n61843 = n41996 | n61771;
  assign n61844 = n41641 | n41996;
  assign n61845 = (n72985 & n61843) | (n72985 & n61844) | (n61843 & n61844);
  assign n41999 = ~n61842 & n61845;
  assign n42000 = x161 & x210;
  assign n42001 = n41999 & n42000;
  assign n42002 = n41999 | n42000;
  assign n42003 = ~n42001 & n42002;
  assign n61846 = n41648 & n42003;
  assign n73115 = (n42003 & n61649) | (n42003 & n61846) | (n61649 & n61846);
  assign n73116 = (n42003 & n61648) | (n42003 & n61846) | (n61648 & n61846);
  assign n73117 = (n72901 & n73115) | (n72901 & n73116) | (n73115 & n73116);
  assign n61848 = n41648 | n42003;
  assign n73118 = n61649 | n61848;
  assign n73119 = n61648 | n61848;
  assign n73120 = (n72901 & n73118) | (n72901 & n73119) | (n73118 & n73119);
  assign n42006 = ~n73117 & n73120;
  assign n42007 = x160 & x211;
  assign n42008 = n42006 & n42007;
  assign n42009 = n42006 | n42007;
  assign n42010 = ~n42008 & n42009;
  assign n42011 = n73053 & n42010;
  assign n42012 = n73053 | n42010;
  assign n42013 = ~n42011 & n42012;
  assign n42014 = x159 & x212;
  assign n42015 = n42013 & n42014;
  assign n42016 = n42013 | n42014;
  assign n42017 = ~n42015 & n42016;
  assign n61766 = n41662 | n41664;
  assign n61850 = n42017 & n61766;
  assign n61851 = n41662 & n42017;
  assign n61852 = (n61561 & n61850) | (n61561 & n61851) | (n61850 & n61851);
  assign n61853 = n42017 | n61766;
  assign n61854 = n41662 | n42017;
  assign n61855 = (n61561 & n61853) | (n61561 & n61854) | (n61853 & n61854);
  assign n42020 = ~n61852 & n61855;
  assign n42021 = x158 & x213;
  assign n42022 = n42020 & n42021;
  assign n42023 = n42020 | n42021;
  assign n42024 = ~n42022 & n42023;
  assign n61856 = n41669 & n42024;
  assign n61857 = (n42024 & n73045) | (n42024 & n61856) | (n73045 & n61856);
  assign n61858 = n41669 | n42024;
  assign n61859 = n73045 | n61858;
  assign n42027 = ~n61857 & n61859;
  assign n42028 = x157 & x214;
  assign n42029 = n42027 & n42028;
  assign n42030 = n42027 | n42028;
  assign n42031 = ~n42029 & n42030;
  assign n61860 = n41676 & n42031;
  assign n61861 = (n42031 & n61663) | (n42031 & n61860) | (n61663 & n61860);
  assign n61862 = n41676 | n42031;
  assign n61863 = n61663 | n61862;
  assign n42034 = ~n61861 & n61863;
  assign n42035 = x156 & x215;
  assign n42036 = n42034 & n42035;
  assign n42037 = n42034 | n42035;
  assign n42038 = ~n42036 & n42037;
  assign n61864 = n41683 & n42038;
  assign n61865 = (n42038 & n61667) | (n42038 & n61864) | (n61667 & n61864);
  assign n61866 = n41683 | n42038;
  assign n61867 = n61667 | n61866;
  assign n42041 = ~n61865 & n61867;
  assign n42042 = x155 & x216;
  assign n42043 = n42041 & n42042;
  assign n42044 = n42041 | n42042;
  assign n42045 = ~n42043 & n42044;
  assign n61868 = n41690 & n42045;
  assign n61869 = (n42045 & n61671) | (n42045 & n61868) | (n61671 & n61868);
  assign n61870 = n41690 | n42045;
  assign n61871 = n61671 | n61870;
  assign n42048 = ~n61869 & n61871;
  assign n42049 = x154 & x217;
  assign n42050 = n42048 & n42049;
  assign n42051 = n42048 | n42049;
  assign n42052 = ~n42050 & n42051;
  assign n61872 = n41697 & n42052;
  assign n61873 = (n42052 & n61675) | (n42052 & n61872) | (n61675 & n61872);
  assign n61874 = n41697 | n42052;
  assign n61875 = n61675 | n61874;
  assign n42055 = ~n61873 & n61875;
  assign n42056 = x153 & x218;
  assign n42057 = n42055 & n42056;
  assign n42058 = n42055 | n42056;
  assign n42059 = ~n42057 & n42058;
  assign n61876 = n41704 & n42059;
  assign n61877 = (n42059 & n61679) | (n42059 & n61876) | (n61679 & n61876);
  assign n61878 = n41704 | n42059;
  assign n61879 = n61679 | n61878;
  assign n42062 = ~n61877 & n61879;
  assign n42063 = x152 & x219;
  assign n42064 = n42062 & n42063;
  assign n42065 = n42062 | n42063;
  assign n42066 = ~n42064 & n42065;
  assign n61880 = n41711 & n42066;
  assign n61881 = (n42066 & n61683) | (n42066 & n61880) | (n61683 & n61880);
  assign n61882 = n41711 | n42066;
  assign n61883 = n61683 | n61882;
  assign n42069 = ~n61881 & n61883;
  assign n42070 = x151 & x220;
  assign n42071 = n42069 & n42070;
  assign n42072 = n42069 | n42070;
  assign n42073 = ~n42071 & n42072;
  assign n61884 = n41718 & n42073;
  assign n61885 = (n42073 & n61687) | (n42073 & n61884) | (n61687 & n61884);
  assign n61886 = n41718 | n42073;
  assign n61887 = n61687 | n61886;
  assign n42076 = ~n61885 & n61887;
  assign n42077 = x150 & x221;
  assign n42078 = n42076 & n42077;
  assign n42079 = n42076 | n42077;
  assign n42080 = ~n42078 & n42079;
  assign n61888 = n41725 & n42080;
  assign n61889 = (n42080 & n61691) | (n42080 & n61888) | (n61691 & n61888);
  assign n61890 = n41725 | n42080;
  assign n61891 = n61691 | n61890;
  assign n42083 = ~n61889 & n61891;
  assign n42084 = x149 & x222;
  assign n42085 = n42083 & n42084;
  assign n42086 = n42083 | n42084;
  assign n42087 = ~n42085 & n42086;
  assign n61892 = n41732 & n42087;
  assign n61893 = (n42087 & n61695) | (n42087 & n61892) | (n61695 & n61892);
  assign n61894 = n41732 | n42087;
  assign n61895 = n61695 | n61894;
  assign n42090 = ~n61893 & n61895;
  assign n42091 = x148 & x223;
  assign n42092 = n42090 & n42091;
  assign n42093 = n42090 | n42091;
  assign n42094 = ~n42092 & n42093;
  assign n61896 = n41739 & n42094;
  assign n61897 = (n42094 & n61699) | (n42094 & n61896) | (n61699 & n61896);
  assign n61898 = n41739 | n42094;
  assign n61899 = n61699 | n61898;
  assign n42097 = ~n61897 & n61899;
  assign n42098 = x147 & x224;
  assign n42099 = n42097 & n42098;
  assign n42100 = n42097 | n42098;
  assign n42101 = ~n42099 & n42100;
  assign n61900 = n41746 & n42101;
  assign n61901 = (n42101 & n61703) | (n42101 & n61900) | (n61703 & n61900);
  assign n61902 = n41746 | n42101;
  assign n61903 = n61703 | n61902;
  assign n42104 = ~n61901 & n61903;
  assign n42105 = x146 & x225;
  assign n42106 = n42104 & n42105;
  assign n42107 = n42104 | n42105;
  assign n42108 = ~n42106 & n42107;
  assign n61904 = n41753 & n42108;
  assign n61905 = (n42108 & n61707) | (n42108 & n61904) | (n61707 & n61904);
  assign n61906 = n41753 | n42108;
  assign n61907 = n61707 | n61906;
  assign n42111 = ~n61905 & n61907;
  assign n42112 = x145 & x226;
  assign n42113 = n42111 & n42112;
  assign n42114 = n42111 | n42112;
  assign n42115 = ~n42113 & n42114;
  assign n61908 = n41760 & n42115;
  assign n61909 = (n42115 & n61711) | (n42115 & n61908) | (n61711 & n61908);
  assign n61910 = n41760 | n42115;
  assign n61911 = n61711 | n61910;
  assign n42118 = ~n61909 & n61911;
  assign n42119 = x144 & x227;
  assign n42120 = n42118 & n42119;
  assign n42121 = n42118 | n42119;
  assign n42122 = ~n42120 & n42121;
  assign n61912 = n41767 & n42122;
  assign n61913 = (n42122 & n61715) | (n42122 & n61912) | (n61715 & n61912);
  assign n61914 = n41767 | n42122;
  assign n61915 = n61715 | n61914;
  assign n42125 = ~n61913 & n61915;
  assign n42126 = x143 & x228;
  assign n42127 = n42125 & n42126;
  assign n42128 = n42125 | n42126;
  assign n42129 = ~n42127 & n42128;
  assign n61916 = n41774 & n42129;
  assign n61917 = (n42129 & n61719) | (n42129 & n61916) | (n61719 & n61916);
  assign n61918 = n41774 | n42129;
  assign n61919 = n61719 | n61918;
  assign n42132 = ~n61917 & n61919;
  assign n42133 = x142 & x229;
  assign n42134 = n42132 & n42133;
  assign n42135 = n42132 | n42133;
  assign n42136 = ~n42134 & n42135;
  assign n61920 = n41781 & n42136;
  assign n61921 = (n42136 & n61723) | (n42136 & n61920) | (n61723 & n61920);
  assign n61922 = n41781 | n42136;
  assign n61923 = n61723 | n61922;
  assign n42139 = ~n61921 & n61923;
  assign n42140 = x141 & x230;
  assign n42141 = n42139 & n42140;
  assign n42142 = n42139 | n42140;
  assign n42143 = ~n42141 & n42142;
  assign n61924 = n41788 & n42143;
  assign n61925 = (n42143 & n61727) | (n42143 & n61924) | (n61727 & n61924);
  assign n61926 = n41788 | n42143;
  assign n61927 = n61727 | n61926;
  assign n42146 = ~n61925 & n61927;
  assign n42147 = x140 & x231;
  assign n42148 = n42146 & n42147;
  assign n42149 = n42146 | n42147;
  assign n42150 = ~n42148 & n42149;
  assign n61928 = n41795 & n42150;
  assign n61929 = (n42150 & n61731) | (n42150 & n61928) | (n61731 & n61928);
  assign n61930 = n41795 | n42150;
  assign n61931 = n61731 | n61930;
  assign n42153 = ~n61929 & n61931;
  assign n42154 = x139 & x232;
  assign n42155 = n42153 & n42154;
  assign n42156 = n42153 | n42154;
  assign n42157 = ~n42155 & n42156;
  assign n61932 = n41802 & n42157;
  assign n61933 = (n42157 & n61735) | (n42157 & n61932) | (n61735 & n61932);
  assign n61934 = n41802 | n42157;
  assign n61935 = n61735 | n61934;
  assign n42160 = ~n61933 & n61935;
  assign n42161 = x138 & x233;
  assign n42162 = n42160 & n42161;
  assign n42163 = n42160 | n42161;
  assign n42164 = ~n42162 & n42163;
  assign n61936 = n41809 & n42164;
  assign n61937 = (n42164 & n61739) | (n42164 & n61936) | (n61739 & n61936);
  assign n61938 = n41809 | n42164;
  assign n61939 = n61739 | n61938;
  assign n42167 = ~n61937 & n61939;
  assign n42168 = x137 & x234;
  assign n42169 = n42167 & n42168;
  assign n42170 = n42167 | n42168;
  assign n42171 = ~n42169 & n42170;
  assign n61940 = n41816 & n42171;
  assign n61941 = (n42171 & n61743) | (n42171 & n61940) | (n61743 & n61940);
  assign n61942 = n41816 | n42171;
  assign n61943 = n61743 | n61942;
  assign n42174 = ~n61941 & n61943;
  assign n42175 = x136 & x235;
  assign n42176 = n42174 & n42175;
  assign n42177 = n42174 | n42175;
  assign n42178 = ~n42176 & n42177;
  assign n61944 = n41823 & n42178;
  assign n61945 = (n42178 & n61747) | (n42178 & n61944) | (n61747 & n61944);
  assign n61946 = n41823 | n42178;
  assign n61947 = n61747 | n61946;
  assign n42181 = ~n61945 & n61947;
  assign n42182 = x135 & x236;
  assign n42183 = n42181 & n42182;
  assign n42184 = n42181 | n42182;
  assign n42185 = ~n42183 & n42184;
  assign n61948 = n41830 & n42185;
  assign n61949 = (n42185 & n61751) | (n42185 & n61948) | (n61751 & n61948);
  assign n61950 = n41830 | n42185;
  assign n61951 = n61751 | n61950;
  assign n42188 = ~n61949 & n61951;
  assign n42189 = x134 & x237;
  assign n42190 = n42188 & n42189;
  assign n42191 = n42188 | n42189;
  assign n42192 = ~n42190 & n42191;
  assign n61952 = n41837 & n42192;
  assign n61953 = (n42192 & n61755) | (n42192 & n61952) | (n61755 & n61952);
  assign n61954 = n41837 | n42192;
  assign n61955 = n61755 | n61954;
  assign n42195 = ~n61953 & n61955;
  assign n42196 = x133 & x238;
  assign n42197 = n42195 & n42196;
  assign n42198 = n42195 | n42196;
  assign n42199 = ~n42197 & n42198;
  assign n61956 = n41844 & n42199;
  assign n61957 = (n42199 & n61759) | (n42199 & n61956) | (n61759 & n61956);
  assign n61958 = n41844 | n42199;
  assign n61959 = n61759 | n61958;
  assign n42202 = ~n61957 & n61959;
  assign n42203 = x132 & x239;
  assign n42204 = n42202 & n42203;
  assign n42205 = n42202 | n42203;
  assign n42206 = ~n42204 & n42205;
  assign n61960 = n41851 & n42206;
  assign n61961 = (n42206 & n61763) | (n42206 & n61960) | (n61763 & n61960);
  assign n61962 = n41851 | n42206;
  assign n61963 = n61763 | n61962;
  assign n42209 = ~n61961 & n61963;
  assign n61970 = n42001 | n42003;
  assign n73123 = n41648 | n42001;
  assign n73124 = (n42001 & n42003) | (n42001 & n73123) | (n42003 & n73123);
  assign n73125 = (n61649 & n61970) | (n61649 & n73124) | (n61970 & n73124);
  assign n73126 = (n61648 & n61970) | (n61648 & n73124) | (n61970 & n73124);
  assign n73127 = (n72901 & n73125) | (n72901 & n73126) | (n73125 & n73126);
  assign n61975 = n41980 | n41982;
  assign n73128 = n41627 | n41980;
  assign n73129 = (n41980 & n41982) | (n41980 & n73128) | (n41982 & n73128);
  assign n73130 = (n61639 & n61975) | (n61639 & n73129) | (n61975 & n73129);
  assign n73131 = (n61638 & n61975) | (n61638 & n73129) | (n61975 & n73129);
  assign n73132 = (n72906 & n73130) | (n72906 & n73131) | (n73130 & n73131);
  assign n61780 = (n61423 & n73060) | (n61423 & n61779) | (n73060 & n61779);
  assign n61980 = n41959 | n41961;
  assign n73133 = n41606 | n41959;
  assign n73134 = (n41959 & n41961) | (n41959 & n73133) | (n41961 & n73133);
  assign n73135 = (n61629 & n61980) | (n61629 & n73134) | (n61980 & n73134);
  assign n73136 = (n61628 & n61980) | (n61628 & n73134) | (n61980 & n73134);
  assign n73137 = (n61363 & n73135) | (n61363 & n73136) | (n73135 & n73136);
  assign n61785 = (n61413 & n73062) | (n61413 & n61784) | (n73062 & n61784);
  assign n61985 = n41938 | n41940;
  assign n73138 = n41585 | n41938;
  assign n73139 = (n41938 & n41940) | (n41938 & n73138) | (n41940 & n73138);
  assign n73140 = (n61619 & n61985) | (n61619 & n73139) | (n61985 & n73139);
  assign n73141 = (n61618 & n61985) | (n61618 & n73139) | (n61985 & n73139);
  assign n73142 = (n61368 & n73140) | (n61368 & n73141) | (n73140 & n73141);
  assign n61790 = (n61403 & n73064) | (n61403 & n61789) | (n73064 & n61789);
  assign n61990 = n41917 | n41919;
  assign n73143 = n41564 | n41917;
  assign n73144 = (n41917 & n41919) | (n41917 & n73143) | (n41919 & n73143);
  assign n73145 = (n61609 & n61990) | (n61609 & n73144) | (n61990 & n73144);
  assign n73146 = (n61608 & n61990) | (n61608 & n73144) | (n61990 & n73144);
  assign n73147 = (n61373 & n73145) | (n61373 & n73146) | (n73145 & n73146);
  assign n42254 = x175 & x197;
  assign n73149 = n42254 & n61796;
  assign n73150 = n41902 & n42254;
  assign n73151 = (n73020 & n73149) | (n73020 & n73150) | (n73149 & n73150);
  assign n73148 = (n41905 & n42254) | (n41905 & n73151) | (n42254 & n73151);
  assign n73152 = (n61794 & n73148) | (n61794 & n73151) | (n73148 & n73151);
  assign n73153 = (n73066 & n73148) | (n73066 & n73151) | (n73148 & n73151);
  assign n73154 = (n61393 & n73152) | (n61393 & n73153) | (n73152 & n73153);
  assign n73156 = n42254 | n61796;
  assign n73157 = n41902 | n42254;
  assign n73158 = (n73020 & n73156) | (n73020 & n73157) | (n73156 & n73157);
  assign n73155 = n41905 | n73158;
  assign n73159 = (n61794 & n73155) | (n61794 & n73158) | (n73155 & n73158);
  assign n73160 = (n73066 & n73155) | (n73066 & n73158) | (n73155 & n73158);
  assign n73161 = (n61393 & n73159) | (n61393 & n73160) | (n73159 & n73160);
  assign n42257 = ~n73154 & n73161;
  assign n62000 = n41910 & n42257;
  assign n62001 = (n42257 & n61802) | (n42257 & n62000) | (n61802 & n62000);
  assign n62002 = n41910 | n42257;
  assign n62003 = n61802 | n62002;
  assign n42260 = ~n62001 & n62003;
  assign n42261 = x174 & x198;
  assign n42262 = n42260 & n42261;
  assign n42263 = n42260 | n42261;
  assign n42264 = ~n42262 & n42263;
  assign n42265 = n73147 & n42264;
  assign n42266 = n73147 | n42264;
  assign n42267 = ~n42265 & n42266;
  assign n42268 = x173 & x199;
  assign n42269 = n42267 & n42268;
  assign n42270 = n42267 | n42268;
  assign n42271 = ~n42269 & n42270;
  assign n61987 = n41924 | n41926;
  assign n62004 = n42271 & n61987;
  assign n62005 = n41924 & n42271;
  assign n62006 = (n61790 & n62004) | (n61790 & n62005) | (n62004 & n62005);
  assign n62007 = n42271 | n61987;
  assign n62008 = n41924 | n42271;
  assign n62009 = (n61790 & n62007) | (n61790 & n62008) | (n62007 & n62008);
  assign n42274 = ~n62006 & n62009;
  assign n42275 = x172 & x200;
  assign n42276 = n42274 & n42275;
  assign n42277 = n42274 | n42275;
  assign n42278 = ~n42276 & n42277;
  assign n62010 = n41931 & n42278;
  assign n62011 = (n42278 & n61812) | (n42278 & n62010) | (n61812 & n62010);
  assign n62012 = n41931 | n42278;
  assign n62013 = n61812 | n62012;
  assign n42281 = ~n62011 & n62013;
  assign n42282 = x171 & x201;
  assign n42283 = n42281 & n42282;
  assign n42284 = n42281 | n42282;
  assign n42285 = ~n42283 & n42284;
  assign n42286 = n73142 & n42285;
  assign n42287 = n73142 | n42285;
  assign n42288 = ~n42286 & n42287;
  assign n42289 = x170 & x202;
  assign n42290 = n42288 & n42289;
  assign n42291 = n42288 | n42289;
  assign n42292 = ~n42290 & n42291;
  assign n61982 = n41945 | n41947;
  assign n62014 = n42292 & n61982;
  assign n62015 = n41945 & n42292;
  assign n62016 = (n61785 & n62014) | (n61785 & n62015) | (n62014 & n62015);
  assign n62017 = n42292 | n61982;
  assign n62018 = n41945 | n42292;
  assign n62019 = (n61785 & n62017) | (n61785 & n62018) | (n62017 & n62018);
  assign n42295 = ~n62016 & n62019;
  assign n42296 = x169 & x203;
  assign n42297 = n42295 & n42296;
  assign n42298 = n42295 | n42296;
  assign n42299 = ~n42297 & n42298;
  assign n62020 = n41952 & n42299;
  assign n62021 = (n42299 & n61822) | (n42299 & n62020) | (n61822 & n62020);
  assign n62022 = n41952 | n42299;
  assign n62023 = n61822 | n62022;
  assign n42302 = ~n62021 & n62023;
  assign n42303 = x168 & x204;
  assign n42304 = n42302 & n42303;
  assign n42305 = n42302 | n42303;
  assign n42306 = ~n42304 & n42305;
  assign n42307 = n73137 & n42306;
  assign n42308 = n73137 | n42306;
  assign n42309 = ~n42307 & n42308;
  assign n42310 = x167 & x205;
  assign n42311 = n42309 & n42310;
  assign n42312 = n42309 | n42310;
  assign n42313 = ~n42311 & n42312;
  assign n61977 = n41966 | n41968;
  assign n62024 = n42313 & n61977;
  assign n62025 = n41966 & n42313;
  assign n62026 = (n61780 & n62024) | (n61780 & n62025) | (n62024 & n62025);
  assign n62027 = n42313 | n61977;
  assign n62028 = n41966 | n42313;
  assign n62029 = (n61780 & n62027) | (n61780 & n62028) | (n62027 & n62028);
  assign n42316 = ~n62026 & n62029;
  assign n42317 = x166 & x206;
  assign n42318 = n42316 & n42317;
  assign n42319 = n42316 | n42317;
  assign n42320 = ~n42318 & n42319;
  assign n62030 = n41973 & n42320;
  assign n62031 = (n42320 & n61832) | (n42320 & n62030) | (n61832 & n62030);
  assign n62032 = n41973 | n42320;
  assign n62033 = n61832 | n62032;
  assign n42323 = ~n62031 & n62033;
  assign n42324 = x165 & x207;
  assign n42325 = n42323 & n42324;
  assign n42326 = n42323 | n42324;
  assign n42327 = ~n42325 & n42326;
  assign n42328 = n73132 & n42327;
  assign n42329 = n73132 | n42327;
  assign n42330 = ~n42328 & n42329;
  assign n42331 = x164 & x208;
  assign n42332 = n42330 & n42331;
  assign n42333 = n42330 | n42331;
  assign n42334 = ~n42332 & n42333;
  assign n61972 = n41987 | n41989;
  assign n62034 = n42334 & n61972;
  assign n62035 = n41987 & n42334;
  assign n62036 = (n73058 & n62034) | (n73058 & n62035) | (n62034 & n62035);
  assign n62037 = n42334 | n61972;
  assign n62038 = n41987 | n42334;
  assign n62039 = (n73058 & n62037) | (n73058 & n62038) | (n62037 & n62038);
  assign n42337 = ~n62036 & n62039;
  assign n42338 = x163 & x209;
  assign n42339 = n42337 & n42338;
  assign n42340 = n42337 | n42338;
  assign n42341 = ~n42339 & n42340;
  assign n62040 = n41994 & n42341;
  assign n73162 = (n42341 & n61841) | (n42341 & n62040) | (n61841 & n62040);
  assign n73163 = (n42341 & n61840) | (n42341 & n62040) | (n61840 & n62040);
  assign n73164 = (n72985 & n73162) | (n72985 & n73163) | (n73162 & n73163);
  assign n62042 = n41994 | n42341;
  assign n73165 = n61841 | n62042;
  assign n73166 = n61840 | n62042;
  assign n73167 = (n72985 & n73165) | (n72985 & n73166) | (n73165 & n73166);
  assign n42344 = ~n73164 & n73167;
  assign n42345 = x162 & x210;
  assign n42346 = n42344 & n42345;
  assign n42347 = n42344 | n42345;
  assign n42348 = ~n42346 & n42347;
  assign n42349 = n73127 & n42348;
  assign n42350 = n73127 | n42348;
  assign n42351 = ~n42349 & n42350;
  assign n42352 = x161 & x211;
  assign n42353 = n42351 & n42352;
  assign n42354 = n42351 | n42352;
  assign n42355 = ~n42353 & n42354;
  assign n61967 = n42008 | n42010;
  assign n62044 = n42355 & n61967;
  assign n62045 = n42008 & n42355;
  assign n62046 = (n73053 & n62044) | (n73053 & n62045) | (n62044 & n62045);
  assign n62047 = n42355 | n61967;
  assign n62048 = n42008 | n42355;
  assign n62049 = (n73053 & n62047) | (n73053 & n62048) | (n62047 & n62048);
  assign n42358 = ~n62046 & n62049;
  assign n42359 = x160 & x212;
  assign n42360 = n42358 & n42359;
  assign n42361 = n42358 | n42359;
  assign n42362 = ~n42360 & n42361;
  assign n62050 = n42015 & n42362;
  assign n73168 = (n42362 & n61851) | (n42362 & n62050) | (n61851 & n62050);
  assign n73169 = (n42362 & n61850) | (n42362 & n62050) | (n61850 & n62050);
  assign n73170 = (n61561 & n73168) | (n61561 & n73169) | (n73168 & n73169);
  assign n62052 = n42015 | n42362;
  assign n73171 = n61851 | n62052;
  assign n73172 = n61850 | n62052;
  assign n73173 = (n61561 & n73171) | (n61561 & n73172) | (n73171 & n73172);
  assign n42365 = ~n73170 & n73173;
  assign n42366 = x159 & x213;
  assign n42367 = n42365 & n42366;
  assign n42368 = n42365 | n42366;
  assign n42369 = ~n42367 & n42368;
  assign n61965 = n42022 | n42024;
  assign n73174 = n42369 & n61965;
  assign n73121 = n41669 | n42022;
  assign n73122 = (n42022 & n42024) | (n42022 & n73121) | (n42024 & n73121);
  assign n73175 = n42369 & n73122;
  assign n73176 = (n73045 & n73174) | (n73045 & n73175) | (n73174 & n73175);
  assign n73177 = n42369 | n61965;
  assign n73178 = n42369 | n73122;
  assign n73179 = (n73045 & n73177) | (n73045 & n73178) | (n73177 & n73178);
  assign n42372 = ~n73176 & n73179;
  assign n42373 = x158 & x214;
  assign n42374 = n42372 & n42373;
  assign n42375 = n42372 | n42373;
  assign n42376 = ~n42374 & n42375;
  assign n62054 = n42029 & n42376;
  assign n73180 = (n42376 & n61860) | (n42376 & n62054) | (n61860 & n62054);
  assign n73181 = (n42031 & n42376) | (n42031 & n62054) | (n42376 & n62054);
  assign n73182 = (n61663 & n73180) | (n61663 & n73181) | (n73180 & n73181);
  assign n62056 = n42029 | n42376;
  assign n73183 = n61860 | n62056;
  assign n73184 = n42031 | n62056;
  assign n73185 = (n61663 & n73183) | (n61663 & n73184) | (n73183 & n73184);
  assign n42379 = ~n73182 & n73185;
  assign n42380 = x157 & x215;
  assign n42381 = n42379 & n42380;
  assign n42382 = n42379 | n42380;
  assign n42383 = ~n42381 & n42382;
  assign n62058 = n42036 & n42383;
  assign n62059 = (n42383 & n61865) | (n42383 & n62058) | (n61865 & n62058);
  assign n62060 = n42036 | n42383;
  assign n62061 = n61865 | n62060;
  assign n42386 = ~n62059 & n62061;
  assign n42387 = x156 & x216;
  assign n42388 = n42386 & n42387;
  assign n42389 = n42386 | n42387;
  assign n42390 = ~n42388 & n42389;
  assign n62062 = n42043 & n42390;
  assign n62063 = (n42390 & n61869) | (n42390 & n62062) | (n61869 & n62062);
  assign n62064 = n42043 | n42390;
  assign n62065 = n61869 | n62064;
  assign n42393 = ~n62063 & n62065;
  assign n42394 = x155 & x217;
  assign n42395 = n42393 & n42394;
  assign n42396 = n42393 | n42394;
  assign n42397 = ~n42395 & n42396;
  assign n62066 = n42050 & n42397;
  assign n62067 = (n42397 & n61873) | (n42397 & n62066) | (n61873 & n62066);
  assign n62068 = n42050 | n42397;
  assign n62069 = n61873 | n62068;
  assign n42400 = ~n62067 & n62069;
  assign n42401 = x154 & x218;
  assign n42402 = n42400 & n42401;
  assign n42403 = n42400 | n42401;
  assign n42404 = ~n42402 & n42403;
  assign n62070 = n42057 & n42404;
  assign n62071 = (n42404 & n61877) | (n42404 & n62070) | (n61877 & n62070);
  assign n62072 = n42057 | n42404;
  assign n62073 = n61877 | n62072;
  assign n42407 = ~n62071 & n62073;
  assign n42408 = x153 & x219;
  assign n42409 = n42407 & n42408;
  assign n42410 = n42407 | n42408;
  assign n42411 = ~n42409 & n42410;
  assign n62074 = n42064 & n42411;
  assign n62075 = (n42411 & n61881) | (n42411 & n62074) | (n61881 & n62074);
  assign n62076 = n42064 | n42411;
  assign n62077 = n61881 | n62076;
  assign n42414 = ~n62075 & n62077;
  assign n42415 = x152 & x220;
  assign n42416 = n42414 & n42415;
  assign n42417 = n42414 | n42415;
  assign n42418 = ~n42416 & n42417;
  assign n62078 = n42071 & n42418;
  assign n62079 = (n42418 & n61885) | (n42418 & n62078) | (n61885 & n62078);
  assign n62080 = n42071 | n42418;
  assign n62081 = n61885 | n62080;
  assign n42421 = ~n62079 & n62081;
  assign n42422 = x151 & x221;
  assign n42423 = n42421 & n42422;
  assign n42424 = n42421 | n42422;
  assign n42425 = ~n42423 & n42424;
  assign n62082 = n42078 & n42425;
  assign n62083 = (n42425 & n61889) | (n42425 & n62082) | (n61889 & n62082);
  assign n62084 = n42078 | n42425;
  assign n62085 = n61889 | n62084;
  assign n42428 = ~n62083 & n62085;
  assign n42429 = x150 & x222;
  assign n42430 = n42428 & n42429;
  assign n42431 = n42428 | n42429;
  assign n42432 = ~n42430 & n42431;
  assign n62086 = n42085 & n42432;
  assign n62087 = (n42432 & n61893) | (n42432 & n62086) | (n61893 & n62086);
  assign n62088 = n42085 | n42432;
  assign n62089 = n61893 | n62088;
  assign n42435 = ~n62087 & n62089;
  assign n42436 = x149 & x223;
  assign n42437 = n42435 & n42436;
  assign n42438 = n42435 | n42436;
  assign n42439 = ~n42437 & n42438;
  assign n62090 = n42092 & n42439;
  assign n62091 = (n42439 & n61897) | (n42439 & n62090) | (n61897 & n62090);
  assign n62092 = n42092 | n42439;
  assign n62093 = n61897 | n62092;
  assign n42442 = ~n62091 & n62093;
  assign n42443 = x148 & x224;
  assign n42444 = n42442 & n42443;
  assign n42445 = n42442 | n42443;
  assign n42446 = ~n42444 & n42445;
  assign n62094 = n42099 & n42446;
  assign n62095 = (n42446 & n61901) | (n42446 & n62094) | (n61901 & n62094);
  assign n62096 = n42099 | n42446;
  assign n62097 = n61901 | n62096;
  assign n42449 = ~n62095 & n62097;
  assign n42450 = x147 & x225;
  assign n42451 = n42449 & n42450;
  assign n42452 = n42449 | n42450;
  assign n42453 = ~n42451 & n42452;
  assign n62098 = n42106 & n42453;
  assign n62099 = (n42453 & n61905) | (n42453 & n62098) | (n61905 & n62098);
  assign n62100 = n42106 | n42453;
  assign n62101 = n61905 | n62100;
  assign n42456 = ~n62099 & n62101;
  assign n42457 = x146 & x226;
  assign n42458 = n42456 & n42457;
  assign n42459 = n42456 | n42457;
  assign n42460 = ~n42458 & n42459;
  assign n62102 = n42113 & n42460;
  assign n62103 = (n42460 & n61909) | (n42460 & n62102) | (n61909 & n62102);
  assign n62104 = n42113 | n42460;
  assign n62105 = n61909 | n62104;
  assign n42463 = ~n62103 & n62105;
  assign n42464 = x145 & x227;
  assign n42465 = n42463 & n42464;
  assign n42466 = n42463 | n42464;
  assign n42467 = ~n42465 & n42466;
  assign n62106 = n42120 & n42467;
  assign n62107 = (n42467 & n61913) | (n42467 & n62106) | (n61913 & n62106);
  assign n62108 = n42120 | n42467;
  assign n62109 = n61913 | n62108;
  assign n42470 = ~n62107 & n62109;
  assign n42471 = x144 & x228;
  assign n42472 = n42470 & n42471;
  assign n42473 = n42470 | n42471;
  assign n42474 = ~n42472 & n42473;
  assign n62110 = n42127 & n42474;
  assign n62111 = (n42474 & n61917) | (n42474 & n62110) | (n61917 & n62110);
  assign n62112 = n42127 | n42474;
  assign n62113 = n61917 | n62112;
  assign n42477 = ~n62111 & n62113;
  assign n42478 = x143 & x229;
  assign n42479 = n42477 & n42478;
  assign n42480 = n42477 | n42478;
  assign n42481 = ~n42479 & n42480;
  assign n62114 = n42134 & n42481;
  assign n62115 = (n42481 & n61921) | (n42481 & n62114) | (n61921 & n62114);
  assign n62116 = n42134 | n42481;
  assign n62117 = n61921 | n62116;
  assign n42484 = ~n62115 & n62117;
  assign n42485 = x142 & x230;
  assign n42486 = n42484 & n42485;
  assign n42487 = n42484 | n42485;
  assign n42488 = ~n42486 & n42487;
  assign n62118 = n42141 & n42488;
  assign n62119 = (n42488 & n61925) | (n42488 & n62118) | (n61925 & n62118);
  assign n62120 = n42141 | n42488;
  assign n62121 = n61925 | n62120;
  assign n42491 = ~n62119 & n62121;
  assign n42492 = x141 & x231;
  assign n42493 = n42491 & n42492;
  assign n42494 = n42491 | n42492;
  assign n42495 = ~n42493 & n42494;
  assign n62122 = n42148 & n42495;
  assign n62123 = (n42495 & n61929) | (n42495 & n62122) | (n61929 & n62122);
  assign n62124 = n42148 | n42495;
  assign n62125 = n61929 | n62124;
  assign n42498 = ~n62123 & n62125;
  assign n42499 = x140 & x232;
  assign n42500 = n42498 & n42499;
  assign n42501 = n42498 | n42499;
  assign n42502 = ~n42500 & n42501;
  assign n62126 = n42155 & n42502;
  assign n62127 = (n42502 & n61933) | (n42502 & n62126) | (n61933 & n62126);
  assign n62128 = n42155 | n42502;
  assign n62129 = n61933 | n62128;
  assign n42505 = ~n62127 & n62129;
  assign n42506 = x139 & x233;
  assign n42507 = n42505 & n42506;
  assign n42508 = n42505 | n42506;
  assign n42509 = ~n42507 & n42508;
  assign n62130 = n42162 & n42509;
  assign n62131 = (n42509 & n61937) | (n42509 & n62130) | (n61937 & n62130);
  assign n62132 = n42162 | n42509;
  assign n62133 = n61937 | n62132;
  assign n42512 = ~n62131 & n62133;
  assign n42513 = x138 & x234;
  assign n42514 = n42512 & n42513;
  assign n42515 = n42512 | n42513;
  assign n42516 = ~n42514 & n42515;
  assign n62134 = n42169 & n42516;
  assign n62135 = (n42516 & n61941) | (n42516 & n62134) | (n61941 & n62134);
  assign n62136 = n42169 | n42516;
  assign n62137 = n61941 | n62136;
  assign n42519 = ~n62135 & n62137;
  assign n42520 = x137 & x235;
  assign n42521 = n42519 & n42520;
  assign n42522 = n42519 | n42520;
  assign n42523 = ~n42521 & n42522;
  assign n62138 = n42176 & n42523;
  assign n62139 = (n42523 & n61945) | (n42523 & n62138) | (n61945 & n62138);
  assign n62140 = n42176 | n42523;
  assign n62141 = n61945 | n62140;
  assign n42526 = ~n62139 & n62141;
  assign n42527 = x136 & x236;
  assign n42528 = n42526 & n42527;
  assign n42529 = n42526 | n42527;
  assign n42530 = ~n42528 & n42529;
  assign n62142 = n42183 & n42530;
  assign n62143 = (n42530 & n61949) | (n42530 & n62142) | (n61949 & n62142);
  assign n62144 = n42183 | n42530;
  assign n62145 = n61949 | n62144;
  assign n42533 = ~n62143 & n62145;
  assign n42534 = x135 & x237;
  assign n42535 = n42533 & n42534;
  assign n42536 = n42533 | n42534;
  assign n42537 = ~n42535 & n42536;
  assign n62146 = n42190 & n42537;
  assign n62147 = (n42537 & n61953) | (n42537 & n62146) | (n61953 & n62146);
  assign n62148 = n42190 | n42537;
  assign n62149 = n61953 | n62148;
  assign n42540 = ~n62147 & n62149;
  assign n42541 = x134 & x238;
  assign n42542 = n42540 & n42541;
  assign n42543 = n42540 | n42541;
  assign n42544 = ~n42542 & n42543;
  assign n62150 = n42197 & n42544;
  assign n62151 = (n42544 & n61957) | (n42544 & n62150) | (n61957 & n62150);
  assign n62152 = n42197 | n42544;
  assign n62153 = n61957 | n62152;
  assign n42547 = ~n62151 & n62153;
  assign n42548 = x133 & x239;
  assign n42549 = n42547 & n42548;
  assign n42550 = n42547 | n42548;
  assign n42551 = ~n42549 & n42550;
  assign n62154 = n42204 & n42551;
  assign n62155 = (n42551 & n61961) | (n42551 & n62154) | (n61961 & n62154);
  assign n62156 = n42204 | n42551;
  assign n62157 = n61961 | n62156;
  assign n42554 = ~n62155 & n62157;
  assign n61966 = (n73045 & n73122) | (n73045 & n61965) | (n73122 & n61965);
  assign n62161 = n42360 | n42362;
  assign n73186 = n42015 | n42360;
  assign n73187 = (n42360 & n42362) | (n42360 & n73186) | (n42362 & n73186);
  assign n73188 = (n61851 & n62161) | (n61851 & n73187) | (n62161 & n73187);
  assign n73189 = (n61850 & n62161) | (n61850 & n73187) | (n62161 & n73187);
  assign n73190 = (n61561 & n73188) | (n61561 & n73189) | (n73188 & n73189);
  assign n62166 = n42339 | n42341;
  assign n73191 = n41994 | n42339;
  assign n73192 = (n42339 & n42341) | (n42339 & n73191) | (n42341 & n73191);
  assign n73193 = (n61841 & n62166) | (n61841 & n73192) | (n62166 & n73192);
  assign n73194 = (n61840 & n62166) | (n61840 & n73192) | (n62166 & n73192);
  assign n73195 = (n72985 & n73193) | (n72985 & n73194) | (n73193 & n73194);
  assign n42598 = x175 & x198;
  assign n73202 = n42257 | n73154;
  assign n73203 = (n41910 & n73154) | (n41910 & n73202) | (n73154 & n73202);
  assign n62188 = n42598 & n73203;
  assign n73204 = n42598 & n73154;
  assign n73205 = (n42257 & n42598) | (n42257 & n73204) | (n42598 & n73204);
  assign n62190 = (n61802 & n62188) | (n61802 & n73205) | (n62188 & n73205);
  assign n62191 = n42598 | n73203;
  assign n73206 = n42598 | n73154;
  assign n73207 = n42257 | n73206;
  assign n62193 = (n61802 & n62191) | (n61802 & n73207) | (n62191 & n73207);
  assign n42601 = ~n62190 & n62193;
  assign n62195 = n42262 & n42601;
  assign n73208 = (n42264 & n42601) | (n42264 & n62195) | (n42601 & n62195);
  assign n62196 = (n73147 & n73208) | (n73147 & n62195) | (n73208 & n62195);
  assign n62198 = n42262 | n42601;
  assign n73209 = n42264 | n62198;
  assign n62199 = (n73147 & n73209) | (n73147 & n62198) | (n73209 & n62198);
  assign n42604 = ~n62196 & n62199;
  assign n42605 = x174 & x199;
  assign n42606 = n42604 & n42605;
  assign n42607 = n42604 | n42605;
  assign n42608 = ~n42606 & n42607;
  assign n62200 = n42269 & n42608;
  assign n73210 = (n42608 & n62005) | (n42608 & n62200) | (n62005 & n62200);
  assign n73211 = (n42608 & n62004) | (n42608 & n62200) | (n62004 & n62200);
  assign n73212 = (n61790 & n73210) | (n61790 & n73211) | (n73210 & n73211);
  assign n62202 = n42269 | n42608;
  assign n73213 = n62005 | n62202;
  assign n73214 = n62004 | n62202;
  assign n73215 = (n61790 & n73213) | (n61790 & n73214) | (n73213 & n73214);
  assign n42611 = ~n73212 & n73215;
  assign n42612 = x173 & x200;
  assign n42613 = n42611 & n42612;
  assign n42614 = n42611 | n42612;
  assign n42615 = ~n42613 & n42614;
  assign n62181 = n42276 | n42278;
  assign n73216 = n42615 & n62181;
  assign n73200 = n41931 | n42276;
  assign n73201 = (n42276 & n42278) | (n42276 & n73200) | (n42278 & n73200);
  assign n73217 = n42615 & n73201;
  assign n73218 = (n61812 & n73216) | (n61812 & n73217) | (n73216 & n73217);
  assign n73219 = n42615 | n62181;
  assign n73220 = n42615 | n73201;
  assign n73221 = (n61812 & n73219) | (n61812 & n73220) | (n73219 & n73220);
  assign n42618 = ~n73218 & n73221;
  assign n42619 = x172 & x201;
  assign n42620 = n42618 & n42619;
  assign n42621 = n42618 | n42619;
  assign n42622 = ~n42620 & n42621;
  assign n62178 = n42283 | n42285;
  assign n62204 = n42622 & n62178;
  assign n62205 = n42283 & n42622;
  assign n62206 = (n73142 & n62204) | (n73142 & n62205) | (n62204 & n62205);
  assign n62207 = n42622 | n62178;
  assign n62208 = n42283 | n42622;
  assign n62209 = (n73142 & n62207) | (n73142 & n62208) | (n62207 & n62208);
  assign n42625 = ~n62206 & n62209;
  assign n42626 = x171 & x202;
  assign n42627 = n42625 & n42626;
  assign n42628 = n42625 | n42626;
  assign n42629 = ~n42627 & n42628;
  assign n62210 = n42290 & n42629;
  assign n73222 = (n42629 & n62015) | (n42629 & n62210) | (n62015 & n62210);
  assign n73223 = (n42629 & n62014) | (n42629 & n62210) | (n62014 & n62210);
  assign n73224 = (n61785 & n73222) | (n61785 & n73223) | (n73222 & n73223);
  assign n62212 = n42290 | n42629;
  assign n73225 = n62015 | n62212;
  assign n73226 = n62014 | n62212;
  assign n73227 = (n61785 & n73225) | (n61785 & n73226) | (n73225 & n73226);
  assign n42632 = ~n73224 & n73227;
  assign n42633 = x170 & x203;
  assign n42634 = n42632 & n42633;
  assign n42635 = n42632 | n42633;
  assign n42636 = ~n42634 & n42635;
  assign n62176 = n42297 | n42299;
  assign n73228 = n42636 & n62176;
  assign n73198 = n41952 | n42297;
  assign n73199 = (n42297 & n42299) | (n42297 & n73198) | (n42299 & n73198);
  assign n73229 = n42636 & n73199;
  assign n73230 = (n61822 & n73228) | (n61822 & n73229) | (n73228 & n73229);
  assign n73231 = n42636 | n62176;
  assign n73232 = n42636 | n73199;
  assign n73233 = (n61822 & n73231) | (n61822 & n73232) | (n73231 & n73232);
  assign n42639 = ~n73230 & n73233;
  assign n42640 = x169 & x204;
  assign n42641 = n42639 & n42640;
  assign n42642 = n42639 | n42640;
  assign n42643 = ~n42641 & n42642;
  assign n62173 = n42304 | n42306;
  assign n62214 = n42643 & n62173;
  assign n62215 = n42304 & n42643;
  assign n62216 = (n73137 & n62214) | (n73137 & n62215) | (n62214 & n62215);
  assign n62217 = n42643 | n62173;
  assign n62218 = n42304 | n42643;
  assign n62219 = (n73137 & n62217) | (n73137 & n62218) | (n62217 & n62218);
  assign n42646 = ~n62216 & n62219;
  assign n42647 = x168 & x205;
  assign n42648 = n42646 & n42647;
  assign n42649 = n42646 | n42647;
  assign n42650 = ~n42648 & n42649;
  assign n62220 = n42311 & n42650;
  assign n73234 = (n42650 & n62025) | (n42650 & n62220) | (n62025 & n62220);
  assign n73235 = (n42650 & n62024) | (n42650 & n62220) | (n62024 & n62220);
  assign n73236 = (n61780 & n73234) | (n61780 & n73235) | (n73234 & n73235);
  assign n62222 = n42311 | n42650;
  assign n73237 = n62025 | n62222;
  assign n73238 = n62024 | n62222;
  assign n73239 = (n61780 & n73237) | (n61780 & n73238) | (n73237 & n73238);
  assign n42653 = ~n73236 & n73239;
  assign n42654 = x167 & x206;
  assign n42655 = n42653 & n42654;
  assign n42656 = n42653 | n42654;
  assign n42657 = ~n42655 & n42656;
  assign n62171 = n42318 | n42320;
  assign n73240 = n42657 & n62171;
  assign n73196 = n41973 | n42318;
  assign n73197 = (n42318 & n42320) | (n42318 & n73196) | (n42320 & n73196);
  assign n73241 = n42657 & n73197;
  assign n73242 = (n61832 & n73240) | (n61832 & n73241) | (n73240 & n73241);
  assign n73243 = n42657 | n62171;
  assign n73244 = n42657 | n73197;
  assign n73245 = (n61832 & n73243) | (n61832 & n73244) | (n73243 & n73244);
  assign n42660 = ~n73242 & n73245;
  assign n42661 = x166 & x207;
  assign n42662 = n42660 & n42661;
  assign n42663 = n42660 | n42661;
  assign n42664 = ~n42662 & n42663;
  assign n62168 = n42325 | n42327;
  assign n62224 = n42664 & n62168;
  assign n62225 = n42325 & n42664;
  assign n62226 = (n73132 & n62224) | (n73132 & n62225) | (n62224 & n62225);
  assign n62227 = n42664 | n62168;
  assign n62228 = n42325 | n42664;
  assign n62229 = (n73132 & n62227) | (n73132 & n62228) | (n62227 & n62228);
  assign n42667 = ~n62226 & n62229;
  assign n42668 = x165 & x208;
  assign n42669 = n42667 & n42668;
  assign n42670 = n42667 | n42668;
  assign n42671 = ~n42669 & n42670;
  assign n62230 = n42332 & n42671;
  assign n73246 = (n42671 & n62035) | (n42671 & n62230) | (n62035 & n62230);
  assign n73247 = (n42671 & n62034) | (n42671 & n62230) | (n62034 & n62230);
  assign n73248 = (n73058 & n73246) | (n73058 & n73247) | (n73246 & n73247);
  assign n62232 = n42332 | n42671;
  assign n73249 = n62035 | n62232;
  assign n73250 = n62034 | n62232;
  assign n73251 = (n73058 & n73249) | (n73058 & n73250) | (n73249 & n73250);
  assign n42674 = ~n73248 & n73251;
  assign n42675 = x164 & x209;
  assign n42676 = n42674 & n42675;
  assign n42677 = n42674 | n42675;
  assign n42678 = ~n42676 & n42677;
  assign n42679 = n73195 & n42678;
  assign n42680 = n73195 | n42678;
  assign n42681 = ~n42679 & n42680;
  assign n42682 = x163 & x210;
  assign n42683 = n42681 & n42682;
  assign n42684 = n42681 | n42682;
  assign n42685 = ~n42683 & n42684;
  assign n62163 = n42346 | n42348;
  assign n62234 = n42685 & n62163;
  assign n62235 = n42346 & n42685;
  assign n62236 = (n73127 & n62234) | (n73127 & n62235) | (n62234 & n62235);
  assign n62237 = n42685 | n62163;
  assign n62238 = n42346 | n42685;
  assign n62239 = (n73127 & n62237) | (n73127 & n62238) | (n62237 & n62238);
  assign n42688 = ~n62236 & n62239;
  assign n42689 = x162 & x211;
  assign n42690 = n42688 & n42689;
  assign n42691 = n42688 | n42689;
  assign n42692 = ~n42690 & n42691;
  assign n62240 = n42353 & n42692;
  assign n73252 = (n42692 & n62045) | (n42692 & n62240) | (n62045 & n62240);
  assign n73253 = (n42692 & n62044) | (n42692 & n62240) | (n62044 & n62240);
  assign n73254 = (n73053 & n73252) | (n73053 & n73253) | (n73252 & n73253);
  assign n62242 = n42353 | n42692;
  assign n73255 = n62045 | n62242;
  assign n73256 = n62044 | n62242;
  assign n73257 = (n73053 & n73255) | (n73053 & n73256) | (n73255 & n73256);
  assign n42695 = ~n73254 & n73257;
  assign n42696 = x161 & x212;
  assign n42697 = n42695 & n42696;
  assign n42698 = n42695 | n42696;
  assign n42699 = ~n42697 & n42698;
  assign n42700 = n73190 & n42699;
  assign n42701 = n73190 | n42699;
  assign n42702 = ~n42700 & n42701;
  assign n42703 = x160 & x213;
  assign n42704 = n42702 & n42703;
  assign n42705 = n42702 | n42703;
  assign n42706 = ~n42704 & n42705;
  assign n62158 = n42367 | n42369;
  assign n62244 = n42706 & n62158;
  assign n62245 = n42367 & n42706;
  assign n62246 = (n61966 & n62244) | (n61966 & n62245) | (n62244 & n62245);
  assign n62247 = n42706 | n62158;
  assign n62248 = n42367 | n42706;
  assign n62249 = (n61966 & n62247) | (n61966 & n62248) | (n62247 & n62248);
  assign n42709 = ~n62246 & n62249;
  assign n42710 = x159 & x214;
  assign n42711 = n42709 & n42710;
  assign n42712 = n42709 | n42710;
  assign n42713 = ~n42711 & n42712;
  assign n62250 = n42374 & n42713;
  assign n62251 = (n42713 & n73182) | (n42713 & n62250) | (n73182 & n62250);
  assign n62252 = n42374 | n42713;
  assign n62253 = n73182 | n62252;
  assign n42716 = ~n62251 & n62253;
  assign n42717 = x158 & x215;
  assign n42718 = n42716 & n42717;
  assign n42719 = n42716 | n42717;
  assign n42720 = ~n42718 & n42719;
  assign n62254 = n42381 & n42720;
  assign n62255 = (n42720 & n62059) | (n42720 & n62254) | (n62059 & n62254);
  assign n62256 = n42381 | n42720;
  assign n62257 = n62059 | n62256;
  assign n42723 = ~n62255 & n62257;
  assign n42724 = x157 & x216;
  assign n42725 = n42723 & n42724;
  assign n42726 = n42723 | n42724;
  assign n42727 = ~n42725 & n42726;
  assign n62258 = n42388 & n42727;
  assign n62259 = (n42727 & n62063) | (n42727 & n62258) | (n62063 & n62258);
  assign n62260 = n42388 | n42727;
  assign n62261 = n62063 | n62260;
  assign n42730 = ~n62259 & n62261;
  assign n42731 = x156 & x217;
  assign n42732 = n42730 & n42731;
  assign n42733 = n42730 | n42731;
  assign n42734 = ~n42732 & n42733;
  assign n62262 = n42395 & n42734;
  assign n62263 = (n42734 & n62067) | (n42734 & n62262) | (n62067 & n62262);
  assign n62264 = n42395 | n42734;
  assign n62265 = n62067 | n62264;
  assign n42737 = ~n62263 & n62265;
  assign n42738 = x155 & x218;
  assign n42739 = n42737 & n42738;
  assign n42740 = n42737 | n42738;
  assign n42741 = ~n42739 & n42740;
  assign n62266 = n42402 & n42741;
  assign n62267 = (n42741 & n62071) | (n42741 & n62266) | (n62071 & n62266);
  assign n62268 = n42402 | n42741;
  assign n62269 = n62071 | n62268;
  assign n42744 = ~n62267 & n62269;
  assign n42745 = x154 & x219;
  assign n42746 = n42744 & n42745;
  assign n42747 = n42744 | n42745;
  assign n42748 = ~n42746 & n42747;
  assign n62270 = n42409 & n42748;
  assign n62271 = (n42748 & n62075) | (n42748 & n62270) | (n62075 & n62270);
  assign n62272 = n42409 | n42748;
  assign n62273 = n62075 | n62272;
  assign n42751 = ~n62271 & n62273;
  assign n42752 = x153 & x220;
  assign n42753 = n42751 & n42752;
  assign n42754 = n42751 | n42752;
  assign n42755 = ~n42753 & n42754;
  assign n62274 = n42416 & n42755;
  assign n62275 = (n42755 & n62079) | (n42755 & n62274) | (n62079 & n62274);
  assign n62276 = n42416 | n42755;
  assign n62277 = n62079 | n62276;
  assign n42758 = ~n62275 & n62277;
  assign n42759 = x152 & x221;
  assign n42760 = n42758 & n42759;
  assign n42761 = n42758 | n42759;
  assign n42762 = ~n42760 & n42761;
  assign n62278 = n42423 & n42762;
  assign n62279 = (n42762 & n62083) | (n42762 & n62278) | (n62083 & n62278);
  assign n62280 = n42423 | n42762;
  assign n62281 = n62083 | n62280;
  assign n42765 = ~n62279 & n62281;
  assign n42766 = x151 & x222;
  assign n42767 = n42765 & n42766;
  assign n42768 = n42765 | n42766;
  assign n42769 = ~n42767 & n42768;
  assign n62282 = n42430 & n42769;
  assign n62283 = (n42769 & n62087) | (n42769 & n62282) | (n62087 & n62282);
  assign n62284 = n42430 | n42769;
  assign n62285 = n62087 | n62284;
  assign n42772 = ~n62283 & n62285;
  assign n42773 = x150 & x223;
  assign n42774 = n42772 & n42773;
  assign n42775 = n42772 | n42773;
  assign n42776 = ~n42774 & n42775;
  assign n62286 = n42437 & n42776;
  assign n62287 = (n42776 & n62091) | (n42776 & n62286) | (n62091 & n62286);
  assign n62288 = n42437 | n42776;
  assign n62289 = n62091 | n62288;
  assign n42779 = ~n62287 & n62289;
  assign n42780 = x149 & x224;
  assign n42781 = n42779 & n42780;
  assign n42782 = n42779 | n42780;
  assign n42783 = ~n42781 & n42782;
  assign n62290 = n42444 & n42783;
  assign n62291 = (n42783 & n62095) | (n42783 & n62290) | (n62095 & n62290);
  assign n62292 = n42444 | n42783;
  assign n62293 = n62095 | n62292;
  assign n42786 = ~n62291 & n62293;
  assign n42787 = x148 & x225;
  assign n42788 = n42786 & n42787;
  assign n42789 = n42786 | n42787;
  assign n42790 = ~n42788 & n42789;
  assign n62294 = n42451 & n42790;
  assign n62295 = (n42790 & n62099) | (n42790 & n62294) | (n62099 & n62294);
  assign n62296 = n42451 | n42790;
  assign n62297 = n62099 | n62296;
  assign n42793 = ~n62295 & n62297;
  assign n42794 = x147 & x226;
  assign n42795 = n42793 & n42794;
  assign n42796 = n42793 | n42794;
  assign n42797 = ~n42795 & n42796;
  assign n62298 = n42458 & n42797;
  assign n62299 = (n42797 & n62103) | (n42797 & n62298) | (n62103 & n62298);
  assign n62300 = n42458 | n42797;
  assign n62301 = n62103 | n62300;
  assign n42800 = ~n62299 & n62301;
  assign n42801 = x146 & x227;
  assign n42802 = n42800 & n42801;
  assign n42803 = n42800 | n42801;
  assign n42804 = ~n42802 & n42803;
  assign n62302 = n42465 & n42804;
  assign n62303 = (n42804 & n62107) | (n42804 & n62302) | (n62107 & n62302);
  assign n62304 = n42465 | n42804;
  assign n62305 = n62107 | n62304;
  assign n42807 = ~n62303 & n62305;
  assign n42808 = x145 & x228;
  assign n42809 = n42807 & n42808;
  assign n42810 = n42807 | n42808;
  assign n42811 = ~n42809 & n42810;
  assign n62306 = n42472 & n42811;
  assign n62307 = (n42811 & n62111) | (n42811 & n62306) | (n62111 & n62306);
  assign n62308 = n42472 | n42811;
  assign n62309 = n62111 | n62308;
  assign n42814 = ~n62307 & n62309;
  assign n42815 = x144 & x229;
  assign n42816 = n42814 & n42815;
  assign n42817 = n42814 | n42815;
  assign n42818 = ~n42816 & n42817;
  assign n62310 = n42479 & n42818;
  assign n62311 = (n42818 & n62115) | (n42818 & n62310) | (n62115 & n62310);
  assign n62312 = n42479 | n42818;
  assign n62313 = n62115 | n62312;
  assign n42821 = ~n62311 & n62313;
  assign n42822 = x143 & x230;
  assign n42823 = n42821 & n42822;
  assign n42824 = n42821 | n42822;
  assign n42825 = ~n42823 & n42824;
  assign n62314 = n42486 & n42825;
  assign n62315 = (n42825 & n62119) | (n42825 & n62314) | (n62119 & n62314);
  assign n62316 = n42486 | n42825;
  assign n62317 = n62119 | n62316;
  assign n42828 = ~n62315 & n62317;
  assign n42829 = x142 & x231;
  assign n42830 = n42828 & n42829;
  assign n42831 = n42828 | n42829;
  assign n42832 = ~n42830 & n42831;
  assign n62318 = n42493 & n42832;
  assign n62319 = (n42832 & n62123) | (n42832 & n62318) | (n62123 & n62318);
  assign n62320 = n42493 | n42832;
  assign n62321 = n62123 | n62320;
  assign n42835 = ~n62319 & n62321;
  assign n42836 = x141 & x232;
  assign n42837 = n42835 & n42836;
  assign n42838 = n42835 | n42836;
  assign n42839 = ~n42837 & n42838;
  assign n62322 = n42500 & n42839;
  assign n62323 = (n42839 & n62127) | (n42839 & n62322) | (n62127 & n62322);
  assign n62324 = n42500 | n42839;
  assign n62325 = n62127 | n62324;
  assign n42842 = ~n62323 & n62325;
  assign n42843 = x140 & x233;
  assign n42844 = n42842 & n42843;
  assign n42845 = n42842 | n42843;
  assign n42846 = ~n42844 & n42845;
  assign n62326 = n42507 & n42846;
  assign n62327 = (n42846 & n62131) | (n42846 & n62326) | (n62131 & n62326);
  assign n62328 = n42507 | n42846;
  assign n62329 = n62131 | n62328;
  assign n42849 = ~n62327 & n62329;
  assign n42850 = x139 & x234;
  assign n42851 = n42849 & n42850;
  assign n42852 = n42849 | n42850;
  assign n42853 = ~n42851 & n42852;
  assign n62330 = n42514 & n42853;
  assign n62331 = (n42853 & n62135) | (n42853 & n62330) | (n62135 & n62330);
  assign n62332 = n42514 | n42853;
  assign n62333 = n62135 | n62332;
  assign n42856 = ~n62331 & n62333;
  assign n42857 = x138 & x235;
  assign n42858 = n42856 & n42857;
  assign n42859 = n42856 | n42857;
  assign n42860 = ~n42858 & n42859;
  assign n62334 = n42521 & n42860;
  assign n62335 = (n42860 & n62139) | (n42860 & n62334) | (n62139 & n62334);
  assign n62336 = n42521 | n42860;
  assign n62337 = n62139 | n62336;
  assign n42863 = ~n62335 & n62337;
  assign n42864 = x137 & x236;
  assign n42865 = n42863 & n42864;
  assign n42866 = n42863 | n42864;
  assign n42867 = ~n42865 & n42866;
  assign n62338 = n42528 & n42867;
  assign n62339 = (n42867 & n62143) | (n42867 & n62338) | (n62143 & n62338);
  assign n62340 = n42528 | n42867;
  assign n62341 = n62143 | n62340;
  assign n42870 = ~n62339 & n62341;
  assign n42871 = x136 & x237;
  assign n42872 = n42870 & n42871;
  assign n42873 = n42870 | n42871;
  assign n42874 = ~n42872 & n42873;
  assign n62342 = n42535 & n42874;
  assign n62343 = (n42874 & n62147) | (n42874 & n62342) | (n62147 & n62342);
  assign n62344 = n42535 | n42874;
  assign n62345 = n62147 | n62344;
  assign n42877 = ~n62343 & n62345;
  assign n42878 = x135 & x238;
  assign n42879 = n42877 & n42878;
  assign n42880 = n42877 | n42878;
  assign n42881 = ~n42879 & n42880;
  assign n62346 = n42542 & n42881;
  assign n62347 = (n42881 & n62151) | (n42881 & n62346) | (n62151 & n62346);
  assign n62348 = n42542 | n42881;
  assign n62349 = n62151 | n62348;
  assign n42884 = ~n62347 & n62349;
  assign n42885 = x134 & x239;
  assign n42886 = n42884 & n42885;
  assign n42887 = n42884 | n42885;
  assign n42888 = ~n42886 & n42887;
  assign n62350 = n42549 & n42888;
  assign n62351 = (n42888 & n62155) | (n42888 & n62350) | (n62155 & n62350);
  assign n62352 = n42549 | n42888;
  assign n62353 = n62155 | n62352;
  assign n42891 = ~n62351 & n62353;
  assign n62360 = n42690 | n42692;
  assign n73260 = n42353 | n42690;
  assign n73261 = (n42690 & n42692) | (n42690 & n73260) | (n42692 & n73260);
  assign n73262 = (n62045 & n62360) | (n62045 & n73261) | (n62360 & n73261);
  assign n73263 = (n62044 & n62360) | (n62044 & n73261) | (n62360 & n73261);
  assign n73264 = (n73053 & n73262) | (n73053 & n73263) | (n73262 & n73263);
  assign n62365 = n42669 | n42671;
  assign n73265 = n42332 | n42669;
  assign n73266 = (n42669 & n42671) | (n42669 & n73265) | (n42671 & n73265);
  assign n73267 = (n62035 & n62365) | (n62035 & n73266) | (n62365 & n73266);
  assign n73268 = (n62034 & n62365) | (n62034 & n73266) | (n62365 & n73266);
  assign n73269 = (n73058 & n73267) | (n73058 & n73268) | (n73267 & n73268);
  assign n62172 = (n61832 & n73197) | (n61832 & n62171) | (n73197 & n62171);
  assign n62370 = n42648 | n42650;
  assign n73270 = n42311 | n42648;
  assign n73271 = (n42648 & n42650) | (n42648 & n73270) | (n42650 & n73270);
  assign n73272 = (n62025 & n62370) | (n62025 & n73271) | (n62370 & n73271);
  assign n73273 = (n62024 & n62370) | (n62024 & n73271) | (n62370 & n73271);
  assign n73274 = (n61780 & n73272) | (n61780 & n73273) | (n73272 & n73273);
  assign n62177 = (n61822 & n73199) | (n61822 & n62176) | (n73199 & n62176);
  assign n62375 = n42627 | n42629;
  assign n73275 = n42290 | n42627;
  assign n73276 = (n42627 & n42629) | (n42627 & n73275) | (n42629 & n73275);
  assign n73277 = (n62015 & n62375) | (n62015 & n73276) | (n62375 & n73276);
  assign n73278 = (n62014 & n62375) | (n62014 & n73276) | (n62375 & n73276);
  assign n73279 = (n61785 & n73277) | (n61785 & n73278) | (n73277 & n73278);
  assign n62182 = (n61812 & n73201) | (n61812 & n62181) | (n73201 & n62181);
  assign n62380 = n42606 | n42608;
  assign n73280 = n42269 | n42606;
  assign n73281 = (n42606 & n42608) | (n42606 & n73280) | (n42608 & n73280);
  assign n73282 = (n62005 & n62380) | (n62005 & n73281) | (n62380 & n73281);
  assign n73283 = (n62004 & n62380) | (n62004 & n73281) | (n62380 & n73281);
  assign n73284 = (n61790 & n73282) | (n61790 & n73283) | (n73282 & n73283);
  assign n42934 = x175 & x199;
  assign n73285 = n42934 & n62188;
  assign n73286 = n42934 & n73205;
  assign n73287 = (n61802 & n73285) | (n61802 & n73286) | (n73285 & n73286);
  assign n73288 = (n42934 & n73208) | (n42934 & n73287) | (n73208 & n73287);
  assign n73289 = (n42934 & n62195) | (n42934 & n73287) | (n62195 & n73287);
  assign n73290 = (n73147 & n73288) | (n73147 & n73289) | (n73288 & n73289);
  assign n73291 = n42934 | n62188;
  assign n73292 = n42934 | n73205;
  assign n73293 = (n61802 & n73291) | (n61802 & n73292) | (n73291 & n73292);
  assign n73294 = n73208 | n73293;
  assign n73295 = n62195 | n73293;
  assign n73296 = (n73147 & n73294) | (n73147 & n73295) | (n73294 & n73295);
  assign n42937 = ~n73290 & n73296;
  assign n42938 = n73284 & n42937;
  assign n42939 = n73284 | n42937;
  assign n42940 = ~n42938 & n42939;
  assign n42941 = x174 & x200;
  assign n42942 = n42940 & n42941;
  assign n42943 = n42940 | n42941;
  assign n42944 = ~n42942 & n42943;
  assign n62377 = n42613 | n42615;
  assign n62386 = n42944 & n62377;
  assign n62387 = n42613 & n42944;
  assign n62388 = (n62182 & n62386) | (n62182 & n62387) | (n62386 & n62387);
  assign n62389 = n42944 | n62377;
  assign n62390 = n42613 | n42944;
  assign n62391 = (n62182 & n62389) | (n62182 & n62390) | (n62389 & n62390);
  assign n42947 = ~n62388 & n62391;
  assign n42948 = x173 & x201;
  assign n42949 = n42947 & n42948;
  assign n42950 = n42947 | n42948;
  assign n42951 = ~n42949 & n42950;
  assign n62392 = n42620 & n42951;
  assign n62393 = (n42951 & n62206) | (n42951 & n62392) | (n62206 & n62392);
  assign n62394 = n42620 | n42951;
  assign n62395 = n62206 | n62394;
  assign n42954 = ~n62393 & n62395;
  assign n42955 = x172 & x202;
  assign n42956 = n42954 & n42955;
  assign n42957 = n42954 | n42955;
  assign n42958 = ~n42956 & n42957;
  assign n42959 = n73279 & n42958;
  assign n42960 = n73279 | n42958;
  assign n42961 = ~n42959 & n42960;
  assign n42962 = x171 & x203;
  assign n42963 = n42961 & n42962;
  assign n42964 = n42961 | n42962;
  assign n42965 = ~n42963 & n42964;
  assign n62372 = n42634 | n42636;
  assign n62396 = n42965 & n62372;
  assign n62397 = n42634 & n42965;
  assign n62398 = (n62177 & n62396) | (n62177 & n62397) | (n62396 & n62397);
  assign n62399 = n42965 | n62372;
  assign n62400 = n42634 | n42965;
  assign n62401 = (n62177 & n62399) | (n62177 & n62400) | (n62399 & n62400);
  assign n42968 = ~n62398 & n62401;
  assign n42969 = x170 & x204;
  assign n42970 = n42968 & n42969;
  assign n42971 = n42968 | n42969;
  assign n42972 = ~n42970 & n42971;
  assign n62402 = n42641 & n42972;
  assign n62403 = (n42972 & n62216) | (n42972 & n62402) | (n62216 & n62402);
  assign n62404 = n42641 | n42972;
  assign n62405 = n62216 | n62404;
  assign n42975 = ~n62403 & n62405;
  assign n42976 = x169 & x205;
  assign n42977 = n42975 & n42976;
  assign n42978 = n42975 | n42976;
  assign n42979 = ~n42977 & n42978;
  assign n42980 = n73274 & n42979;
  assign n42981 = n73274 | n42979;
  assign n42982 = ~n42980 & n42981;
  assign n42983 = x168 & x206;
  assign n42984 = n42982 & n42983;
  assign n42985 = n42982 | n42983;
  assign n42986 = ~n42984 & n42985;
  assign n62367 = n42655 | n42657;
  assign n62406 = n42986 & n62367;
  assign n62407 = n42655 & n42986;
  assign n62408 = (n62172 & n62406) | (n62172 & n62407) | (n62406 & n62407);
  assign n62409 = n42986 | n62367;
  assign n62410 = n42655 | n42986;
  assign n62411 = (n62172 & n62409) | (n62172 & n62410) | (n62409 & n62410);
  assign n42989 = ~n62408 & n62411;
  assign n42990 = x167 & x207;
  assign n42991 = n42989 & n42990;
  assign n42992 = n42989 | n42990;
  assign n42993 = ~n42991 & n42992;
  assign n62412 = n42662 & n42993;
  assign n62413 = (n42993 & n62226) | (n42993 & n62412) | (n62226 & n62412);
  assign n62414 = n42662 | n42993;
  assign n62415 = n62226 | n62414;
  assign n42996 = ~n62413 & n62415;
  assign n42997 = x166 & x208;
  assign n42998 = n42996 & n42997;
  assign n42999 = n42996 | n42997;
  assign n43000 = ~n42998 & n42999;
  assign n43001 = n73269 & n43000;
  assign n43002 = n73269 | n43000;
  assign n43003 = ~n43001 & n43002;
  assign n43004 = x165 & x209;
  assign n43005 = n43003 & n43004;
  assign n43006 = n43003 | n43004;
  assign n43007 = ~n43005 & n43006;
  assign n62362 = n42676 | n42678;
  assign n62416 = n43007 & n62362;
  assign n62417 = n42676 & n43007;
  assign n62418 = (n73195 & n62416) | (n73195 & n62417) | (n62416 & n62417);
  assign n62419 = n43007 | n62362;
  assign n62420 = n42676 | n43007;
  assign n62421 = (n73195 & n62419) | (n73195 & n62420) | (n62419 & n62420);
  assign n43010 = ~n62418 & n62421;
  assign n43011 = x164 & x210;
  assign n43012 = n43010 & n43011;
  assign n43013 = n43010 | n43011;
  assign n43014 = ~n43012 & n43013;
  assign n62422 = n42683 & n43014;
  assign n73297 = (n43014 & n62235) | (n43014 & n62422) | (n62235 & n62422);
  assign n73298 = (n43014 & n62234) | (n43014 & n62422) | (n62234 & n62422);
  assign n73299 = (n73127 & n73297) | (n73127 & n73298) | (n73297 & n73298);
  assign n62424 = n42683 | n43014;
  assign n73300 = n62235 | n62424;
  assign n73301 = n62234 | n62424;
  assign n73302 = (n73127 & n73300) | (n73127 & n73301) | (n73300 & n73301);
  assign n43017 = ~n73299 & n73302;
  assign n43018 = x163 & x211;
  assign n43019 = n43017 & n43018;
  assign n43020 = n43017 | n43018;
  assign n43021 = ~n43019 & n43020;
  assign n43022 = n73264 & n43021;
  assign n43023 = n73264 | n43021;
  assign n43024 = ~n43022 & n43023;
  assign n43025 = x162 & x212;
  assign n43026 = n43024 & n43025;
  assign n43027 = n43024 | n43025;
  assign n43028 = ~n43026 & n43027;
  assign n62357 = n42697 | n42699;
  assign n62426 = n43028 & n62357;
  assign n62427 = n42697 & n43028;
  assign n62428 = (n73190 & n62426) | (n73190 & n62427) | (n62426 & n62427);
  assign n62429 = n43028 | n62357;
  assign n62430 = n42697 | n43028;
  assign n62431 = (n73190 & n62429) | (n73190 & n62430) | (n62429 & n62430);
  assign n43031 = ~n62428 & n62431;
  assign n43032 = x161 & x213;
  assign n43033 = n43031 & n43032;
  assign n43034 = n43031 | n43032;
  assign n43035 = ~n43033 & n43034;
  assign n62432 = n42704 & n43035;
  assign n73303 = (n43035 & n62245) | (n43035 & n62432) | (n62245 & n62432);
  assign n73304 = (n43035 & n62244) | (n43035 & n62432) | (n62244 & n62432);
  assign n73305 = (n61966 & n73303) | (n61966 & n73304) | (n73303 & n73304);
  assign n62434 = n42704 | n43035;
  assign n73306 = n62245 | n62434;
  assign n73307 = n62244 | n62434;
  assign n73308 = (n61966 & n73306) | (n61966 & n73307) | (n73306 & n73307);
  assign n43038 = ~n73305 & n73308;
  assign n43039 = x160 & x214;
  assign n43040 = n43038 & n43039;
  assign n43041 = n43038 | n43039;
  assign n43042 = ~n43040 & n43041;
  assign n62355 = n42711 | n42713;
  assign n73309 = n43042 & n62355;
  assign n73258 = n42374 | n42711;
  assign n73259 = (n42711 & n42713) | (n42711 & n73258) | (n42713 & n73258);
  assign n73310 = n43042 & n73259;
  assign n73311 = (n73182 & n73309) | (n73182 & n73310) | (n73309 & n73310);
  assign n73312 = n43042 | n62355;
  assign n73313 = n43042 | n73259;
  assign n73314 = (n73182 & n73312) | (n73182 & n73313) | (n73312 & n73313);
  assign n43045 = ~n73311 & n73314;
  assign n43046 = x159 & x215;
  assign n43047 = n43045 & n43046;
  assign n43048 = n43045 | n43046;
  assign n43049 = ~n43047 & n43048;
  assign n62436 = n42718 & n43049;
  assign n73315 = (n43049 & n62254) | (n43049 & n62436) | (n62254 & n62436);
  assign n73316 = (n42720 & n43049) | (n42720 & n62436) | (n43049 & n62436);
  assign n73317 = (n62059 & n73315) | (n62059 & n73316) | (n73315 & n73316);
  assign n62438 = n42718 | n43049;
  assign n73318 = n62254 | n62438;
  assign n73319 = n42720 | n62438;
  assign n73320 = (n62059 & n73318) | (n62059 & n73319) | (n73318 & n73319);
  assign n43052 = ~n73317 & n73320;
  assign n43053 = x158 & x216;
  assign n43054 = n43052 & n43053;
  assign n43055 = n43052 | n43053;
  assign n43056 = ~n43054 & n43055;
  assign n62440 = n42725 & n43056;
  assign n62441 = (n43056 & n62259) | (n43056 & n62440) | (n62259 & n62440);
  assign n62442 = n42725 | n43056;
  assign n62443 = n62259 | n62442;
  assign n43059 = ~n62441 & n62443;
  assign n43060 = x157 & x217;
  assign n43061 = n43059 & n43060;
  assign n43062 = n43059 | n43060;
  assign n43063 = ~n43061 & n43062;
  assign n62444 = n42732 & n43063;
  assign n62445 = (n43063 & n62263) | (n43063 & n62444) | (n62263 & n62444);
  assign n62446 = n42732 | n43063;
  assign n62447 = n62263 | n62446;
  assign n43066 = ~n62445 & n62447;
  assign n43067 = x156 & x218;
  assign n43068 = n43066 & n43067;
  assign n43069 = n43066 | n43067;
  assign n43070 = ~n43068 & n43069;
  assign n62448 = n42739 & n43070;
  assign n62449 = (n43070 & n62267) | (n43070 & n62448) | (n62267 & n62448);
  assign n62450 = n42739 | n43070;
  assign n62451 = n62267 | n62450;
  assign n43073 = ~n62449 & n62451;
  assign n43074 = x155 & x219;
  assign n43075 = n43073 & n43074;
  assign n43076 = n43073 | n43074;
  assign n43077 = ~n43075 & n43076;
  assign n62452 = n42746 & n43077;
  assign n62453 = (n43077 & n62271) | (n43077 & n62452) | (n62271 & n62452);
  assign n62454 = n42746 | n43077;
  assign n62455 = n62271 | n62454;
  assign n43080 = ~n62453 & n62455;
  assign n43081 = x154 & x220;
  assign n43082 = n43080 & n43081;
  assign n43083 = n43080 | n43081;
  assign n43084 = ~n43082 & n43083;
  assign n62456 = n42753 & n43084;
  assign n62457 = (n43084 & n62275) | (n43084 & n62456) | (n62275 & n62456);
  assign n62458 = n42753 | n43084;
  assign n62459 = n62275 | n62458;
  assign n43087 = ~n62457 & n62459;
  assign n43088 = x153 & x221;
  assign n43089 = n43087 & n43088;
  assign n43090 = n43087 | n43088;
  assign n43091 = ~n43089 & n43090;
  assign n62460 = n42760 & n43091;
  assign n62461 = (n43091 & n62279) | (n43091 & n62460) | (n62279 & n62460);
  assign n62462 = n42760 | n43091;
  assign n62463 = n62279 | n62462;
  assign n43094 = ~n62461 & n62463;
  assign n43095 = x152 & x222;
  assign n43096 = n43094 & n43095;
  assign n43097 = n43094 | n43095;
  assign n43098 = ~n43096 & n43097;
  assign n62464 = n42767 & n43098;
  assign n62465 = (n43098 & n62283) | (n43098 & n62464) | (n62283 & n62464);
  assign n62466 = n42767 | n43098;
  assign n62467 = n62283 | n62466;
  assign n43101 = ~n62465 & n62467;
  assign n43102 = x151 & x223;
  assign n43103 = n43101 & n43102;
  assign n43104 = n43101 | n43102;
  assign n43105 = ~n43103 & n43104;
  assign n62468 = n42774 & n43105;
  assign n62469 = (n43105 & n62287) | (n43105 & n62468) | (n62287 & n62468);
  assign n62470 = n42774 | n43105;
  assign n62471 = n62287 | n62470;
  assign n43108 = ~n62469 & n62471;
  assign n43109 = x150 & x224;
  assign n43110 = n43108 & n43109;
  assign n43111 = n43108 | n43109;
  assign n43112 = ~n43110 & n43111;
  assign n62472 = n42781 & n43112;
  assign n62473 = (n43112 & n62291) | (n43112 & n62472) | (n62291 & n62472);
  assign n62474 = n42781 | n43112;
  assign n62475 = n62291 | n62474;
  assign n43115 = ~n62473 & n62475;
  assign n43116 = x149 & x225;
  assign n43117 = n43115 & n43116;
  assign n43118 = n43115 | n43116;
  assign n43119 = ~n43117 & n43118;
  assign n62476 = n42788 & n43119;
  assign n62477 = (n43119 & n62295) | (n43119 & n62476) | (n62295 & n62476);
  assign n62478 = n42788 | n43119;
  assign n62479 = n62295 | n62478;
  assign n43122 = ~n62477 & n62479;
  assign n43123 = x148 & x226;
  assign n43124 = n43122 & n43123;
  assign n43125 = n43122 | n43123;
  assign n43126 = ~n43124 & n43125;
  assign n62480 = n42795 & n43126;
  assign n62481 = (n43126 & n62299) | (n43126 & n62480) | (n62299 & n62480);
  assign n62482 = n42795 | n43126;
  assign n62483 = n62299 | n62482;
  assign n43129 = ~n62481 & n62483;
  assign n43130 = x147 & x227;
  assign n43131 = n43129 & n43130;
  assign n43132 = n43129 | n43130;
  assign n43133 = ~n43131 & n43132;
  assign n62484 = n42802 & n43133;
  assign n62485 = (n43133 & n62303) | (n43133 & n62484) | (n62303 & n62484);
  assign n62486 = n42802 | n43133;
  assign n62487 = n62303 | n62486;
  assign n43136 = ~n62485 & n62487;
  assign n43137 = x146 & x228;
  assign n43138 = n43136 & n43137;
  assign n43139 = n43136 | n43137;
  assign n43140 = ~n43138 & n43139;
  assign n62488 = n42809 & n43140;
  assign n62489 = (n43140 & n62307) | (n43140 & n62488) | (n62307 & n62488);
  assign n62490 = n42809 | n43140;
  assign n62491 = n62307 | n62490;
  assign n43143 = ~n62489 & n62491;
  assign n43144 = x145 & x229;
  assign n43145 = n43143 & n43144;
  assign n43146 = n43143 | n43144;
  assign n43147 = ~n43145 & n43146;
  assign n62492 = n42816 & n43147;
  assign n62493 = (n43147 & n62311) | (n43147 & n62492) | (n62311 & n62492);
  assign n62494 = n42816 | n43147;
  assign n62495 = n62311 | n62494;
  assign n43150 = ~n62493 & n62495;
  assign n43151 = x144 & x230;
  assign n43152 = n43150 & n43151;
  assign n43153 = n43150 | n43151;
  assign n43154 = ~n43152 & n43153;
  assign n62496 = n42823 & n43154;
  assign n62497 = (n43154 & n62315) | (n43154 & n62496) | (n62315 & n62496);
  assign n62498 = n42823 | n43154;
  assign n62499 = n62315 | n62498;
  assign n43157 = ~n62497 & n62499;
  assign n43158 = x143 & x231;
  assign n43159 = n43157 & n43158;
  assign n43160 = n43157 | n43158;
  assign n43161 = ~n43159 & n43160;
  assign n62500 = n42830 & n43161;
  assign n62501 = (n43161 & n62319) | (n43161 & n62500) | (n62319 & n62500);
  assign n62502 = n42830 | n43161;
  assign n62503 = n62319 | n62502;
  assign n43164 = ~n62501 & n62503;
  assign n43165 = x142 & x232;
  assign n43166 = n43164 & n43165;
  assign n43167 = n43164 | n43165;
  assign n43168 = ~n43166 & n43167;
  assign n62504 = n42837 & n43168;
  assign n62505 = (n43168 & n62323) | (n43168 & n62504) | (n62323 & n62504);
  assign n62506 = n42837 | n43168;
  assign n62507 = n62323 | n62506;
  assign n43171 = ~n62505 & n62507;
  assign n43172 = x141 & x233;
  assign n43173 = n43171 & n43172;
  assign n43174 = n43171 | n43172;
  assign n43175 = ~n43173 & n43174;
  assign n62508 = n42844 & n43175;
  assign n62509 = (n43175 & n62327) | (n43175 & n62508) | (n62327 & n62508);
  assign n62510 = n42844 | n43175;
  assign n62511 = n62327 | n62510;
  assign n43178 = ~n62509 & n62511;
  assign n43179 = x140 & x234;
  assign n43180 = n43178 & n43179;
  assign n43181 = n43178 | n43179;
  assign n43182 = ~n43180 & n43181;
  assign n62512 = n42851 & n43182;
  assign n62513 = (n43182 & n62331) | (n43182 & n62512) | (n62331 & n62512);
  assign n62514 = n42851 | n43182;
  assign n62515 = n62331 | n62514;
  assign n43185 = ~n62513 & n62515;
  assign n43186 = x139 & x235;
  assign n43187 = n43185 & n43186;
  assign n43188 = n43185 | n43186;
  assign n43189 = ~n43187 & n43188;
  assign n62516 = n42858 & n43189;
  assign n62517 = (n43189 & n62335) | (n43189 & n62516) | (n62335 & n62516);
  assign n62518 = n42858 | n43189;
  assign n62519 = n62335 | n62518;
  assign n43192 = ~n62517 & n62519;
  assign n43193 = x138 & x236;
  assign n43194 = n43192 & n43193;
  assign n43195 = n43192 | n43193;
  assign n43196 = ~n43194 & n43195;
  assign n62520 = n42865 & n43196;
  assign n62521 = (n43196 & n62339) | (n43196 & n62520) | (n62339 & n62520);
  assign n62522 = n42865 | n43196;
  assign n62523 = n62339 | n62522;
  assign n43199 = ~n62521 & n62523;
  assign n43200 = x137 & x237;
  assign n43201 = n43199 & n43200;
  assign n43202 = n43199 | n43200;
  assign n43203 = ~n43201 & n43202;
  assign n62524 = n42872 & n43203;
  assign n62525 = (n43203 & n62343) | (n43203 & n62524) | (n62343 & n62524);
  assign n62526 = n42872 | n43203;
  assign n62527 = n62343 | n62526;
  assign n43206 = ~n62525 & n62527;
  assign n43207 = x136 & x238;
  assign n43208 = n43206 & n43207;
  assign n43209 = n43206 | n43207;
  assign n43210 = ~n43208 & n43209;
  assign n62528 = n42879 & n43210;
  assign n62529 = (n43210 & n62347) | (n43210 & n62528) | (n62347 & n62528);
  assign n62530 = n42879 | n43210;
  assign n62531 = n62347 | n62530;
  assign n43213 = ~n62529 & n62531;
  assign n43214 = x135 & x239;
  assign n43215 = n43213 & n43214;
  assign n43216 = n43213 | n43214;
  assign n43217 = ~n43215 & n43216;
  assign n62532 = n42886 & n43217;
  assign n62533 = (n43217 & n62351) | (n43217 & n62532) | (n62351 & n62532);
  assign n62534 = n42886 | n43217;
  assign n62535 = n62351 | n62534;
  assign n43220 = ~n62533 & n62535;
  assign n62356 = (n73182 & n73259) | (n73182 & n62355) | (n73259 & n62355);
  assign n62539 = n43033 | n43035;
  assign n73321 = n42704 | n43033;
  assign n73322 = (n43033 & n43035) | (n43033 & n73321) | (n43035 & n73321);
  assign n73323 = (n62245 & n62539) | (n62245 & n73322) | (n62539 & n73322);
  assign n73324 = (n62244 & n62539) | (n62244 & n73322) | (n62539 & n73322);
  assign n73325 = (n61966 & n73323) | (n61966 & n73324) | (n73323 & n73324);
  assign n62544 = n43012 | n43014;
  assign n73326 = n42683 | n43012;
  assign n73327 = (n43012 & n43014) | (n43012 & n73326) | (n43014 & n73326);
  assign n73328 = (n62235 & n62544) | (n62235 & n73327) | (n62544 & n73327);
  assign n73329 = (n62234 & n62544) | (n62234 & n73327) | (n62544 & n73327);
  assign n73330 = (n73127 & n73328) | (n73127 & n73329) | (n73328 & n73329);
  assign n43262 = x175 & x200;
  assign n73337 = n43262 & n73290;
  assign n73338 = (n42937 & n43262) | (n42937 & n73337) | (n43262 & n73337);
  assign n62564 = n43262 & n73290;
  assign n62565 = (n73284 & n73338) | (n73284 & n62564) | (n73338 & n62564);
  assign n73339 = n43262 | n73290;
  assign n73340 = n42937 | n73339;
  assign n62567 = n43262 | n73290;
  assign n62568 = (n73284 & n73340) | (n73284 & n62567) | (n73340 & n62567);
  assign n43265 = ~n62565 & n62568;
  assign n62569 = n42942 & n43265;
  assign n73341 = (n43265 & n62387) | (n43265 & n62569) | (n62387 & n62569);
  assign n73342 = (n43265 & n62386) | (n43265 & n62569) | (n62386 & n62569);
  assign n73343 = (n62182 & n73341) | (n62182 & n73342) | (n73341 & n73342);
  assign n62571 = n42942 | n43265;
  assign n73344 = n62387 | n62571;
  assign n73345 = n62386 | n62571;
  assign n73346 = (n62182 & n73344) | (n62182 & n73345) | (n73344 & n73345);
  assign n43268 = ~n73343 & n73346;
  assign n43269 = x174 & x201;
  assign n43270 = n43268 & n43269;
  assign n43271 = n43268 | n43269;
  assign n43272 = ~n43270 & n43271;
  assign n62559 = n42949 | n42951;
  assign n73347 = n43272 & n62559;
  assign n73335 = n42620 | n42949;
  assign n73336 = (n42949 & n42951) | (n42949 & n73335) | (n42951 & n73335);
  assign n73348 = n43272 & n73336;
  assign n73349 = (n62206 & n73347) | (n62206 & n73348) | (n73347 & n73348);
  assign n73350 = n43272 | n62559;
  assign n73351 = n43272 | n73336;
  assign n73352 = (n62206 & n73350) | (n62206 & n73351) | (n73350 & n73351);
  assign n43275 = ~n73349 & n73352;
  assign n43276 = x173 & x202;
  assign n43277 = n43275 & n43276;
  assign n43278 = n43275 | n43276;
  assign n43279 = ~n43277 & n43278;
  assign n62556 = n42956 | n42958;
  assign n62573 = n43279 & n62556;
  assign n62574 = n42956 & n43279;
  assign n62575 = (n73279 & n62573) | (n73279 & n62574) | (n62573 & n62574);
  assign n62576 = n43279 | n62556;
  assign n62577 = n42956 | n43279;
  assign n62578 = (n73279 & n62576) | (n73279 & n62577) | (n62576 & n62577);
  assign n43282 = ~n62575 & n62578;
  assign n43283 = x172 & x203;
  assign n43284 = n43282 & n43283;
  assign n43285 = n43282 | n43283;
  assign n43286 = ~n43284 & n43285;
  assign n62579 = n42963 & n43286;
  assign n73353 = (n43286 & n62397) | (n43286 & n62579) | (n62397 & n62579);
  assign n73354 = (n43286 & n62396) | (n43286 & n62579) | (n62396 & n62579);
  assign n73355 = (n62177 & n73353) | (n62177 & n73354) | (n73353 & n73354);
  assign n62581 = n42963 | n43286;
  assign n73356 = n62397 | n62581;
  assign n73357 = n62396 | n62581;
  assign n73358 = (n62177 & n73356) | (n62177 & n73357) | (n73356 & n73357);
  assign n43289 = ~n73355 & n73358;
  assign n43290 = x171 & x204;
  assign n43291 = n43289 & n43290;
  assign n43292 = n43289 | n43290;
  assign n43293 = ~n43291 & n43292;
  assign n62554 = n42970 | n42972;
  assign n73359 = n43293 & n62554;
  assign n73333 = n42641 | n42970;
  assign n73334 = (n42970 & n42972) | (n42970 & n73333) | (n42972 & n73333);
  assign n73360 = n43293 & n73334;
  assign n73361 = (n62216 & n73359) | (n62216 & n73360) | (n73359 & n73360);
  assign n73362 = n43293 | n62554;
  assign n73363 = n43293 | n73334;
  assign n73364 = (n62216 & n73362) | (n62216 & n73363) | (n73362 & n73363);
  assign n43296 = ~n73361 & n73364;
  assign n43297 = x170 & x205;
  assign n43298 = n43296 & n43297;
  assign n43299 = n43296 | n43297;
  assign n43300 = ~n43298 & n43299;
  assign n62551 = n42977 | n42979;
  assign n62583 = n43300 & n62551;
  assign n62584 = n42977 & n43300;
  assign n62585 = (n73274 & n62583) | (n73274 & n62584) | (n62583 & n62584);
  assign n62586 = n43300 | n62551;
  assign n62587 = n42977 | n43300;
  assign n62588 = (n73274 & n62586) | (n73274 & n62587) | (n62586 & n62587);
  assign n43303 = ~n62585 & n62588;
  assign n43304 = x169 & x206;
  assign n43305 = n43303 & n43304;
  assign n43306 = n43303 | n43304;
  assign n43307 = ~n43305 & n43306;
  assign n62589 = n42984 & n43307;
  assign n73365 = (n43307 & n62407) | (n43307 & n62589) | (n62407 & n62589);
  assign n73366 = (n43307 & n62406) | (n43307 & n62589) | (n62406 & n62589);
  assign n73367 = (n62172 & n73365) | (n62172 & n73366) | (n73365 & n73366);
  assign n62591 = n42984 | n43307;
  assign n73368 = n62407 | n62591;
  assign n73369 = n62406 | n62591;
  assign n73370 = (n62172 & n73368) | (n62172 & n73369) | (n73368 & n73369);
  assign n43310 = ~n73367 & n73370;
  assign n43311 = x168 & x207;
  assign n43312 = n43310 & n43311;
  assign n43313 = n43310 | n43311;
  assign n43314 = ~n43312 & n43313;
  assign n62549 = n42991 | n42993;
  assign n73371 = n43314 & n62549;
  assign n73331 = n42662 | n42991;
  assign n73332 = (n42991 & n42993) | (n42991 & n73331) | (n42993 & n73331);
  assign n73372 = n43314 & n73332;
  assign n73373 = (n62226 & n73371) | (n62226 & n73372) | (n73371 & n73372);
  assign n73374 = n43314 | n62549;
  assign n73375 = n43314 | n73332;
  assign n73376 = (n62226 & n73374) | (n62226 & n73375) | (n73374 & n73375);
  assign n43317 = ~n73373 & n73376;
  assign n43318 = x167 & x208;
  assign n43319 = n43317 & n43318;
  assign n43320 = n43317 | n43318;
  assign n43321 = ~n43319 & n43320;
  assign n62546 = n42998 | n43000;
  assign n62593 = n43321 & n62546;
  assign n62594 = n42998 & n43321;
  assign n62595 = (n73269 & n62593) | (n73269 & n62594) | (n62593 & n62594);
  assign n62596 = n43321 | n62546;
  assign n62597 = n42998 | n43321;
  assign n62598 = (n73269 & n62596) | (n73269 & n62597) | (n62596 & n62597);
  assign n43324 = ~n62595 & n62598;
  assign n43325 = x166 & x209;
  assign n43326 = n43324 & n43325;
  assign n43327 = n43324 | n43325;
  assign n43328 = ~n43326 & n43327;
  assign n62599 = n43005 & n43328;
  assign n73377 = (n43328 & n62417) | (n43328 & n62599) | (n62417 & n62599);
  assign n73378 = (n43328 & n62416) | (n43328 & n62599) | (n62416 & n62599);
  assign n73379 = (n73195 & n73377) | (n73195 & n73378) | (n73377 & n73378);
  assign n62601 = n43005 | n43328;
  assign n73380 = n62417 | n62601;
  assign n73381 = n62416 | n62601;
  assign n73382 = (n73195 & n73380) | (n73195 & n73381) | (n73380 & n73381);
  assign n43331 = ~n73379 & n73382;
  assign n43332 = x165 & x210;
  assign n43333 = n43331 & n43332;
  assign n43334 = n43331 | n43332;
  assign n43335 = ~n43333 & n43334;
  assign n43336 = n73330 & n43335;
  assign n43337 = n73330 | n43335;
  assign n43338 = ~n43336 & n43337;
  assign n43339 = x164 & x211;
  assign n43340 = n43338 & n43339;
  assign n43341 = n43338 | n43339;
  assign n43342 = ~n43340 & n43341;
  assign n62541 = n43019 | n43021;
  assign n62603 = n43342 & n62541;
  assign n62604 = n43019 & n43342;
  assign n62605 = (n73264 & n62603) | (n73264 & n62604) | (n62603 & n62604);
  assign n62606 = n43342 | n62541;
  assign n62607 = n43019 | n43342;
  assign n62608 = (n73264 & n62606) | (n73264 & n62607) | (n62606 & n62607);
  assign n43345 = ~n62605 & n62608;
  assign n43346 = x163 & x212;
  assign n43347 = n43345 & n43346;
  assign n43348 = n43345 | n43346;
  assign n43349 = ~n43347 & n43348;
  assign n62609 = n43026 & n43349;
  assign n73383 = (n43349 & n62427) | (n43349 & n62609) | (n62427 & n62609);
  assign n73384 = (n43349 & n62426) | (n43349 & n62609) | (n62426 & n62609);
  assign n73385 = (n73190 & n73383) | (n73190 & n73384) | (n73383 & n73384);
  assign n62611 = n43026 | n43349;
  assign n73386 = n62427 | n62611;
  assign n73387 = n62426 | n62611;
  assign n73388 = (n73190 & n73386) | (n73190 & n73387) | (n73386 & n73387);
  assign n43352 = ~n73385 & n73388;
  assign n43353 = x162 & x213;
  assign n43354 = n43352 & n43353;
  assign n43355 = n43352 | n43353;
  assign n43356 = ~n43354 & n43355;
  assign n43357 = n73325 & n43356;
  assign n43358 = n73325 | n43356;
  assign n43359 = ~n43357 & n43358;
  assign n43360 = x161 & x214;
  assign n43361 = n43359 & n43360;
  assign n43362 = n43359 | n43360;
  assign n43363 = ~n43361 & n43362;
  assign n62536 = n43040 | n43042;
  assign n62613 = n43363 & n62536;
  assign n62614 = n43040 & n43363;
  assign n62615 = (n62356 & n62613) | (n62356 & n62614) | (n62613 & n62614);
  assign n62616 = n43363 | n62536;
  assign n62617 = n43040 | n43363;
  assign n62618 = (n62356 & n62616) | (n62356 & n62617) | (n62616 & n62617);
  assign n43366 = ~n62615 & n62618;
  assign n43367 = x160 & x215;
  assign n43368 = n43366 & n43367;
  assign n43369 = n43366 | n43367;
  assign n43370 = ~n43368 & n43369;
  assign n62619 = n43047 & n43370;
  assign n62620 = (n43370 & n73317) | (n43370 & n62619) | (n73317 & n62619);
  assign n62621 = n43047 | n43370;
  assign n62622 = n73317 | n62621;
  assign n43373 = ~n62620 & n62622;
  assign n43374 = x159 & x216;
  assign n43375 = n43373 & n43374;
  assign n43376 = n43373 | n43374;
  assign n43377 = ~n43375 & n43376;
  assign n62623 = n43054 & n43377;
  assign n62624 = (n43377 & n62441) | (n43377 & n62623) | (n62441 & n62623);
  assign n62625 = n43054 | n43377;
  assign n62626 = n62441 | n62625;
  assign n43380 = ~n62624 & n62626;
  assign n43381 = x158 & x217;
  assign n43382 = n43380 & n43381;
  assign n43383 = n43380 | n43381;
  assign n43384 = ~n43382 & n43383;
  assign n62627 = n43061 & n43384;
  assign n62628 = (n43384 & n62445) | (n43384 & n62627) | (n62445 & n62627);
  assign n62629 = n43061 | n43384;
  assign n62630 = n62445 | n62629;
  assign n43387 = ~n62628 & n62630;
  assign n43388 = x157 & x218;
  assign n43389 = n43387 & n43388;
  assign n43390 = n43387 | n43388;
  assign n43391 = ~n43389 & n43390;
  assign n62631 = n43068 & n43391;
  assign n62632 = (n43391 & n62449) | (n43391 & n62631) | (n62449 & n62631);
  assign n62633 = n43068 | n43391;
  assign n62634 = n62449 | n62633;
  assign n43394 = ~n62632 & n62634;
  assign n43395 = x156 & x219;
  assign n43396 = n43394 & n43395;
  assign n43397 = n43394 | n43395;
  assign n43398 = ~n43396 & n43397;
  assign n62635 = n43075 & n43398;
  assign n62636 = (n43398 & n62453) | (n43398 & n62635) | (n62453 & n62635);
  assign n62637 = n43075 | n43398;
  assign n62638 = n62453 | n62637;
  assign n43401 = ~n62636 & n62638;
  assign n43402 = x155 & x220;
  assign n43403 = n43401 & n43402;
  assign n43404 = n43401 | n43402;
  assign n43405 = ~n43403 & n43404;
  assign n62639 = n43082 & n43405;
  assign n62640 = (n43405 & n62457) | (n43405 & n62639) | (n62457 & n62639);
  assign n62641 = n43082 | n43405;
  assign n62642 = n62457 | n62641;
  assign n43408 = ~n62640 & n62642;
  assign n43409 = x154 & x221;
  assign n43410 = n43408 & n43409;
  assign n43411 = n43408 | n43409;
  assign n43412 = ~n43410 & n43411;
  assign n62643 = n43089 & n43412;
  assign n62644 = (n43412 & n62461) | (n43412 & n62643) | (n62461 & n62643);
  assign n62645 = n43089 | n43412;
  assign n62646 = n62461 | n62645;
  assign n43415 = ~n62644 & n62646;
  assign n43416 = x153 & x222;
  assign n43417 = n43415 & n43416;
  assign n43418 = n43415 | n43416;
  assign n43419 = ~n43417 & n43418;
  assign n62647 = n43096 & n43419;
  assign n62648 = (n43419 & n62465) | (n43419 & n62647) | (n62465 & n62647);
  assign n62649 = n43096 | n43419;
  assign n62650 = n62465 | n62649;
  assign n43422 = ~n62648 & n62650;
  assign n43423 = x152 & x223;
  assign n43424 = n43422 & n43423;
  assign n43425 = n43422 | n43423;
  assign n43426 = ~n43424 & n43425;
  assign n62651 = n43103 & n43426;
  assign n62652 = (n43426 & n62469) | (n43426 & n62651) | (n62469 & n62651);
  assign n62653 = n43103 | n43426;
  assign n62654 = n62469 | n62653;
  assign n43429 = ~n62652 & n62654;
  assign n43430 = x151 & x224;
  assign n43431 = n43429 & n43430;
  assign n43432 = n43429 | n43430;
  assign n43433 = ~n43431 & n43432;
  assign n62655 = n43110 & n43433;
  assign n62656 = (n43433 & n62473) | (n43433 & n62655) | (n62473 & n62655);
  assign n62657 = n43110 | n43433;
  assign n62658 = n62473 | n62657;
  assign n43436 = ~n62656 & n62658;
  assign n43437 = x150 & x225;
  assign n43438 = n43436 & n43437;
  assign n43439 = n43436 | n43437;
  assign n43440 = ~n43438 & n43439;
  assign n62659 = n43117 & n43440;
  assign n62660 = (n43440 & n62477) | (n43440 & n62659) | (n62477 & n62659);
  assign n62661 = n43117 | n43440;
  assign n62662 = n62477 | n62661;
  assign n43443 = ~n62660 & n62662;
  assign n43444 = x149 & x226;
  assign n43445 = n43443 & n43444;
  assign n43446 = n43443 | n43444;
  assign n43447 = ~n43445 & n43446;
  assign n62663 = n43124 & n43447;
  assign n62664 = (n43447 & n62481) | (n43447 & n62663) | (n62481 & n62663);
  assign n62665 = n43124 | n43447;
  assign n62666 = n62481 | n62665;
  assign n43450 = ~n62664 & n62666;
  assign n43451 = x148 & x227;
  assign n43452 = n43450 & n43451;
  assign n43453 = n43450 | n43451;
  assign n43454 = ~n43452 & n43453;
  assign n62667 = n43131 & n43454;
  assign n62668 = (n43454 & n62485) | (n43454 & n62667) | (n62485 & n62667);
  assign n62669 = n43131 | n43454;
  assign n62670 = n62485 | n62669;
  assign n43457 = ~n62668 & n62670;
  assign n43458 = x147 & x228;
  assign n43459 = n43457 & n43458;
  assign n43460 = n43457 | n43458;
  assign n43461 = ~n43459 & n43460;
  assign n62671 = n43138 & n43461;
  assign n62672 = (n43461 & n62489) | (n43461 & n62671) | (n62489 & n62671);
  assign n62673 = n43138 | n43461;
  assign n62674 = n62489 | n62673;
  assign n43464 = ~n62672 & n62674;
  assign n43465 = x146 & x229;
  assign n43466 = n43464 & n43465;
  assign n43467 = n43464 | n43465;
  assign n43468 = ~n43466 & n43467;
  assign n62675 = n43145 & n43468;
  assign n62676 = (n43468 & n62493) | (n43468 & n62675) | (n62493 & n62675);
  assign n62677 = n43145 | n43468;
  assign n62678 = n62493 | n62677;
  assign n43471 = ~n62676 & n62678;
  assign n43472 = x145 & x230;
  assign n43473 = n43471 & n43472;
  assign n43474 = n43471 | n43472;
  assign n43475 = ~n43473 & n43474;
  assign n62679 = n43152 & n43475;
  assign n62680 = (n43475 & n62497) | (n43475 & n62679) | (n62497 & n62679);
  assign n62681 = n43152 | n43475;
  assign n62682 = n62497 | n62681;
  assign n43478 = ~n62680 & n62682;
  assign n43479 = x144 & x231;
  assign n43480 = n43478 & n43479;
  assign n43481 = n43478 | n43479;
  assign n43482 = ~n43480 & n43481;
  assign n62683 = n43159 & n43482;
  assign n62684 = (n43482 & n62501) | (n43482 & n62683) | (n62501 & n62683);
  assign n62685 = n43159 | n43482;
  assign n62686 = n62501 | n62685;
  assign n43485 = ~n62684 & n62686;
  assign n43486 = x143 & x232;
  assign n43487 = n43485 & n43486;
  assign n43488 = n43485 | n43486;
  assign n43489 = ~n43487 & n43488;
  assign n62687 = n43166 & n43489;
  assign n62688 = (n43489 & n62505) | (n43489 & n62687) | (n62505 & n62687);
  assign n62689 = n43166 | n43489;
  assign n62690 = n62505 | n62689;
  assign n43492 = ~n62688 & n62690;
  assign n43493 = x142 & x233;
  assign n43494 = n43492 & n43493;
  assign n43495 = n43492 | n43493;
  assign n43496 = ~n43494 & n43495;
  assign n62691 = n43173 & n43496;
  assign n62692 = (n43496 & n62509) | (n43496 & n62691) | (n62509 & n62691);
  assign n62693 = n43173 | n43496;
  assign n62694 = n62509 | n62693;
  assign n43499 = ~n62692 & n62694;
  assign n43500 = x141 & x234;
  assign n43501 = n43499 & n43500;
  assign n43502 = n43499 | n43500;
  assign n43503 = ~n43501 & n43502;
  assign n62695 = n43180 & n43503;
  assign n62696 = (n43503 & n62513) | (n43503 & n62695) | (n62513 & n62695);
  assign n62697 = n43180 | n43503;
  assign n62698 = n62513 | n62697;
  assign n43506 = ~n62696 & n62698;
  assign n43507 = x140 & x235;
  assign n43508 = n43506 & n43507;
  assign n43509 = n43506 | n43507;
  assign n43510 = ~n43508 & n43509;
  assign n62699 = n43187 & n43510;
  assign n62700 = (n43510 & n62517) | (n43510 & n62699) | (n62517 & n62699);
  assign n62701 = n43187 | n43510;
  assign n62702 = n62517 | n62701;
  assign n43513 = ~n62700 & n62702;
  assign n43514 = x139 & x236;
  assign n43515 = n43513 & n43514;
  assign n43516 = n43513 | n43514;
  assign n43517 = ~n43515 & n43516;
  assign n62703 = n43194 & n43517;
  assign n62704 = (n43517 & n62521) | (n43517 & n62703) | (n62521 & n62703);
  assign n62705 = n43194 | n43517;
  assign n62706 = n62521 | n62705;
  assign n43520 = ~n62704 & n62706;
  assign n43521 = x138 & x237;
  assign n43522 = n43520 & n43521;
  assign n43523 = n43520 | n43521;
  assign n43524 = ~n43522 & n43523;
  assign n62707 = n43201 & n43524;
  assign n62708 = (n43524 & n62525) | (n43524 & n62707) | (n62525 & n62707);
  assign n62709 = n43201 | n43524;
  assign n62710 = n62525 | n62709;
  assign n43527 = ~n62708 & n62710;
  assign n43528 = x137 & x238;
  assign n43529 = n43527 & n43528;
  assign n43530 = n43527 | n43528;
  assign n43531 = ~n43529 & n43530;
  assign n62711 = n43208 & n43531;
  assign n62712 = (n43531 & n62529) | (n43531 & n62711) | (n62529 & n62711);
  assign n62713 = n43208 | n43531;
  assign n62714 = n62529 | n62713;
  assign n43534 = ~n62712 & n62714;
  assign n43535 = x136 & x239;
  assign n43536 = n43534 & n43535;
  assign n43537 = n43534 | n43535;
  assign n43538 = ~n43536 & n43537;
  assign n62715 = n43215 & n43538;
  assign n62716 = (n43538 & n62533) | (n43538 & n62715) | (n62533 & n62715);
  assign n62717 = n43215 | n43538;
  assign n62718 = n62533 | n62717;
  assign n43541 = ~n62716 & n62718;
  assign n62725 = n43347 | n43349;
  assign n73391 = n43026 | n43347;
  assign n73392 = (n43347 & n43349) | (n43347 & n73391) | (n43349 & n73391);
  assign n73393 = (n62427 & n62725) | (n62427 & n73392) | (n62725 & n73392);
  assign n73394 = (n62426 & n62725) | (n62426 & n73392) | (n62725 & n73392);
  assign n73395 = (n73190 & n73393) | (n73190 & n73394) | (n73393 & n73394);
  assign n62730 = n43326 | n43328;
  assign n73396 = n43005 | n43326;
  assign n73397 = (n43326 & n43328) | (n43326 & n73396) | (n43328 & n73396);
  assign n73398 = (n62417 & n62730) | (n62417 & n73397) | (n62730 & n73397);
  assign n73399 = (n62416 & n62730) | (n62416 & n73397) | (n62730 & n73397);
  assign n73400 = (n73195 & n73398) | (n73195 & n73399) | (n73398 & n73399);
  assign n62550 = (n62226 & n73332) | (n62226 & n62549) | (n73332 & n62549);
  assign n62735 = n43305 | n43307;
  assign n73401 = n42984 | n43305;
  assign n73402 = (n43305 & n43307) | (n43305 & n73401) | (n43307 & n73401);
  assign n73403 = (n62407 & n62735) | (n62407 & n73402) | (n62735 & n73402);
  assign n73404 = (n62406 & n62735) | (n62406 & n73402) | (n62735 & n73402);
  assign n73405 = (n62172 & n73403) | (n62172 & n73404) | (n73403 & n73404);
  assign n62555 = (n62216 & n73334) | (n62216 & n62554) | (n73334 & n62554);
  assign n62740 = n43284 | n43286;
  assign n73406 = n42963 | n43284;
  assign n73407 = (n43284 & n43286) | (n43284 & n73406) | (n43286 & n73406);
  assign n73408 = (n62397 & n62740) | (n62397 & n73407) | (n62740 & n73407);
  assign n73409 = (n62396 & n62740) | (n62396 & n73407) | (n62740 & n73407);
  assign n73410 = (n62177 & n73408) | (n62177 & n73409) | (n73408 & n73409);
  assign n43582 = x175 & x201;
  assign n62745 = n43265 | n62565;
  assign n73411 = (n42942 & n62565) | (n42942 & n62745) | (n62565 & n62745);
  assign n62747 = n43582 & n73411;
  assign n73412 = n43582 & n62565;
  assign n73413 = (n43265 & n43582) | (n43265 & n73412) | (n43582 & n73412);
  assign n73414 = (n62387 & n62747) | (n62387 & n73413) | (n62747 & n73413);
  assign n73415 = (n62386 & n62747) | (n62386 & n73413) | (n62747 & n73413);
  assign n73416 = (n62182 & n73414) | (n62182 & n73415) | (n73414 & n73415);
  assign n62750 = n43582 | n73411;
  assign n73417 = n43582 | n62565;
  assign n73418 = n43265 | n73417;
  assign n73419 = (n62387 & n62750) | (n62387 & n73418) | (n62750 & n73418);
  assign n73420 = (n62386 & n62750) | (n62386 & n73418) | (n62750 & n73418);
  assign n73421 = (n62182 & n73419) | (n62182 & n73420) | (n73419 & n73420);
  assign n43585 = ~n73416 & n73421;
  assign n62754 = n43270 & n43585;
  assign n73422 = (n43272 & n43585) | (n43272 & n62754) | (n43585 & n62754);
  assign n73423 = (n62559 & n62754) | (n62559 & n73422) | (n62754 & n73422);
  assign n73424 = (n62754 & n73336) | (n62754 & n73422) | (n73336 & n73422);
  assign n73425 = (n62206 & n73423) | (n62206 & n73424) | (n73423 & n73424);
  assign n62757 = n43270 | n43585;
  assign n73426 = n43272 | n62757;
  assign n73427 = (n62559 & n62757) | (n62559 & n73426) | (n62757 & n73426);
  assign n73428 = (n62757 & n73336) | (n62757 & n73426) | (n73336 & n73426);
  assign n73429 = (n62206 & n73427) | (n62206 & n73428) | (n73427 & n73428);
  assign n43588 = ~n73425 & n73429;
  assign n43589 = x174 & x202;
  assign n43590 = n43588 & n43589;
  assign n43591 = n43588 | n43589;
  assign n43592 = ~n43590 & n43591;
  assign n62759 = n43277 & n43592;
  assign n62760 = (n43592 & n62575) | (n43592 & n62759) | (n62575 & n62759);
  assign n62761 = n43277 | n43592;
  assign n62762 = n62575 | n62761;
  assign n43595 = ~n62760 & n62762;
  assign n43596 = x173 & x203;
  assign n43597 = n43595 & n43596;
  assign n43598 = n43595 | n43596;
  assign n43599 = ~n43597 & n43598;
  assign n43600 = n73410 & n43599;
  assign n43601 = n73410 | n43599;
  assign n43602 = ~n43600 & n43601;
  assign n43603 = x172 & x204;
  assign n43604 = n43602 & n43603;
  assign n43605 = n43602 | n43603;
  assign n43606 = ~n43604 & n43605;
  assign n62737 = n43291 | n43293;
  assign n62763 = n43606 & n62737;
  assign n62764 = n43291 & n43606;
  assign n62765 = (n62555 & n62763) | (n62555 & n62764) | (n62763 & n62764);
  assign n62766 = n43606 | n62737;
  assign n62767 = n43291 | n43606;
  assign n62768 = (n62555 & n62766) | (n62555 & n62767) | (n62766 & n62767);
  assign n43609 = ~n62765 & n62768;
  assign n43610 = x171 & x205;
  assign n43611 = n43609 & n43610;
  assign n43612 = n43609 | n43610;
  assign n43613 = ~n43611 & n43612;
  assign n62769 = n43298 & n43613;
  assign n62770 = (n43613 & n62585) | (n43613 & n62769) | (n62585 & n62769);
  assign n62771 = n43298 | n43613;
  assign n62772 = n62585 | n62771;
  assign n43616 = ~n62770 & n62772;
  assign n43617 = x170 & x206;
  assign n43618 = n43616 & n43617;
  assign n43619 = n43616 | n43617;
  assign n43620 = ~n43618 & n43619;
  assign n43621 = n73405 & n43620;
  assign n43622 = n73405 | n43620;
  assign n43623 = ~n43621 & n43622;
  assign n43624 = x169 & x207;
  assign n43625 = n43623 & n43624;
  assign n43626 = n43623 | n43624;
  assign n43627 = ~n43625 & n43626;
  assign n62732 = n43312 | n43314;
  assign n62773 = n43627 & n62732;
  assign n62774 = n43312 & n43627;
  assign n62775 = (n62550 & n62773) | (n62550 & n62774) | (n62773 & n62774);
  assign n62776 = n43627 | n62732;
  assign n62777 = n43312 | n43627;
  assign n62778 = (n62550 & n62776) | (n62550 & n62777) | (n62776 & n62777);
  assign n43630 = ~n62775 & n62778;
  assign n43631 = x168 & x208;
  assign n43632 = n43630 & n43631;
  assign n43633 = n43630 | n43631;
  assign n43634 = ~n43632 & n43633;
  assign n62779 = n43319 & n43634;
  assign n62780 = (n43634 & n62595) | (n43634 & n62779) | (n62595 & n62779);
  assign n62781 = n43319 | n43634;
  assign n62782 = n62595 | n62781;
  assign n43637 = ~n62780 & n62782;
  assign n43638 = x167 & x209;
  assign n43639 = n43637 & n43638;
  assign n43640 = n43637 | n43638;
  assign n43641 = ~n43639 & n43640;
  assign n43642 = n73400 & n43641;
  assign n43643 = n73400 | n43641;
  assign n43644 = ~n43642 & n43643;
  assign n43645 = x166 & x210;
  assign n43646 = n43644 & n43645;
  assign n43647 = n43644 | n43645;
  assign n43648 = ~n43646 & n43647;
  assign n62727 = n43333 | n43335;
  assign n62783 = n43648 & n62727;
  assign n62784 = n43333 & n43648;
  assign n62785 = (n73330 & n62783) | (n73330 & n62784) | (n62783 & n62784);
  assign n62786 = n43648 | n62727;
  assign n62787 = n43333 | n43648;
  assign n62788 = (n73330 & n62786) | (n73330 & n62787) | (n62786 & n62787);
  assign n43651 = ~n62785 & n62788;
  assign n43652 = x165 & x211;
  assign n43653 = n43651 & n43652;
  assign n43654 = n43651 | n43652;
  assign n43655 = ~n43653 & n43654;
  assign n62789 = n43340 & n43655;
  assign n73430 = (n43655 & n62604) | (n43655 & n62789) | (n62604 & n62789);
  assign n73431 = (n43655 & n62603) | (n43655 & n62789) | (n62603 & n62789);
  assign n73432 = (n73264 & n73430) | (n73264 & n73431) | (n73430 & n73431);
  assign n62791 = n43340 | n43655;
  assign n73433 = n62604 | n62791;
  assign n73434 = n62603 | n62791;
  assign n73435 = (n73264 & n73433) | (n73264 & n73434) | (n73433 & n73434);
  assign n43658 = ~n73432 & n73435;
  assign n43659 = x164 & x212;
  assign n43660 = n43658 & n43659;
  assign n43661 = n43658 | n43659;
  assign n43662 = ~n43660 & n43661;
  assign n43663 = n73395 & n43662;
  assign n43664 = n73395 | n43662;
  assign n43665 = ~n43663 & n43664;
  assign n43666 = x163 & x213;
  assign n43667 = n43665 & n43666;
  assign n43668 = n43665 | n43666;
  assign n43669 = ~n43667 & n43668;
  assign n62722 = n43354 | n43356;
  assign n62793 = n43669 & n62722;
  assign n62794 = n43354 & n43669;
  assign n62795 = (n73325 & n62793) | (n73325 & n62794) | (n62793 & n62794);
  assign n62796 = n43669 | n62722;
  assign n62797 = n43354 | n43669;
  assign n62798 = (n73325 & n62796) | (n73325 & n62797) | (n62796 & n62797);
  assign n43672 = ~n62795 & n62798;
  assign n43673 = x162 & x214;
  assign n43674 = n43672 & n43673;
  assign n43675 = n43672 | n43673;
  assign n43676 = ~n43674 & n43675;
  assign n62799 = n43361 & n43676;
  assign n73436 = (n43676 & n62614) | (n43676 & n62799) | (n62614 & n62799);
  assign n73437 = (n43676 & n62613) | (n43676 & n62799) | (n62613 & n62799);
  assign n73438 = (n62356 & n73436) | (n62356 & n73437) | (n73436 & n73437);
  assign n62801 = n43361 | n43676;
  assign n73439 = n62614 | n62801;
  assign n73440 = n62613 | n62801;
  assign n73441 = (n62356 & n73439) | (n62356 & n73440) | (n73439 & n73440);
  assign n43679 = ~n73438 & n73441;
  assign n43680 = x161 & x215;
  assign n43681 = n43679 & n43680;
  assign n43682 = n43679 | n43680;
  assign n43683 = ~n43681 & n43682;
  assign n62720 = n43368 | n43370;
  assign n73442 = n43683 & n62720;
  assign n73389 = n43047 | n43368;
  assign n73390 = (n43368 & n43370) | (n43368 & n73389) | (n43370 & n73389);
  assign n73443 = n43683 & n73390;
  assign n73444 = (n73317 & n73442) | (n73317 & n73443) | (n73442 & n73443);
  assign n73445 = n43683 | n62720;
  assign n73446 = n43683 | n73390;
  assign n73447 = (n73317 & n73445) | (n73317 & n73446) | (n73445 & n73446);
  assign n43686 = ~n73444 & n73447;
  assign n43687 = x160 & x216;
  assign n43688 = n43686 & n43687;
  assign n43689 = n43686 | n43687;
  assign n43690 = ~n43688 & n43689;
  assign n62803 = n43375 & n43690;
  assign n73448 = (n43690 & n62623) | (n43690 & n62803) | (n62623 & n62803);
  assign n73449 = (n43377 & n43690) | (n43377 & n62803) | (n43690 & n62803);
  assign n73450 = (n62441 & n73448) | (n62441 & n73449) | (n73448 & n73449);
  assign n62805 = n43375 | n43690;
  assign n73451 = n62623 | n62805;
  assign n73452 = n43377 | n62805;
  assign n73453 = (n62441 & n73451) | (n62441 & n73452) | (n73451 & n73452);
  assign n43693 = ~n73450 & n73453;
  assign n43694 = x159 & x217;
  assign n43695 = n43693 & n43694;
  assign n43696 = n43693 | n43694;
  assign n43697 = ~n43695 & n43696;
  assign n62807 = n43382 & n43697;
  assign n62808 = (n43697 & n62628) | (n43697 & n62807) | (n62628 & n62807);
  assign n62809 = n43382 | n43697;
  assign n62810 = n62628 | n62809;
  assign n43700 = ~n62808 & n62810;
  assign n43701 = x158 & x218;
  assign n43702 = n43700 & n43701;
  assign n43703 = n43700 | n43701;
  assign n43704 = ~n43702 & n43703;
  assign n62811 = n43389 & n43704;
  assign n62812 = (n43704 & n62632) | (n43704 & n62811) | (n62632 & n62811);
  assign n62813 = n43389 | n43704;
  assign n62814 = n62632 | n62813;
  assign n43707 = ~n62812 & n62814;
  assign n43708 = x157 & x219;
  assign n43709 = n43707 & n43708;
  assign n43710 = n43707 | n43708;
  assign n43711 = ~n43709 & n43710;
  assign n62815 = n43396 & n43711;
  assign n62816 = (n43711 & n62636) | (n43711 & n62815) | (n62636 & n62815);
  assign n62817 = n43396 | n43711;
  assign n62818 = n62636 | n62817;
  assign n43714 = ~n62816 & n62818;
  assign n43715 = x156 & x220;
  assign n43716 = n43714 & n43715;
  assign n43717 = n43714 | n43715;
  assign n43718 = ~n43716 & n43717;
  assign n62819 = n43403 & n43718;
  assign n62820 = (n43718 & n62640) | (n43718 & n62819) | (n62640 & n62819);
  assign n62821 = n43403 | n43718;
  assign n62822 = n62640 | n62821;
  assign n43721 = ~n62820 & n62822;
  assign n43722 = x155 & x221;
  assign n43723 = n43721 & n43722;
  assign n43724 = n43721 | n43722;
  assign n43725 = ~n43723 & n43724;
  assign n62823 = n43410 & n43725;
  assign n62824 = (n43725 & n62644) | (n43725 & n62823) | (n62644 & n62823);
  assign n62825 = n43410 | n43725;
  assign n62826 = n62644 | n62825;
  assign n43728 = ~n62824 & n62826;
  assign n43729 = x154 & x222;
  assign n43730 = n43728 & n43729;
  assign n43731 = n43728 | n43729;
  assign n43732 = ~n43730 & n43731;
  assign n62827 = n43417 & n43732;
  assign n62828 = (n43732 & n62648) | (n43732 & n62827) | (n62648 & n62827);
  assign n62829 = n43417 | n43732;
  assign n62830 = n62648 | n62829;
  assign n43735 = ~n62828 & n62830;
  assign n43736 = x153 & x223;
  assign n43737 = n43735 & n43736;
  assign n43738 = n43735 | n43736;
  assign n43739 = ~n43737 & n43738;
  assign n62831 = n43424 & n43739;
  assign n62832 = (n43739 & n62652) | (n43739 & n62831) | (n62652 & n62831);
  assign n62833 = n43424 | n43739;
  assign n62834 = n62652 | n62833;
  assign n43742 = ~n62832 & n62834;
  assign n43743 = x152 & x224;
  assign n43744 = n43742 & n43743;
  assign n43745 = n43742 | n43743;
  assign n43746 = ~n43744 & n43745;
  assign n62835 = n43431 & n43746;
  assign n62836 = (n43746 & n62656) | (n43746 & n62835) | (n62656 & n62835);
  assign n62837 = n43431 | n43746;
  assign n62838 = n62656 | n62837;
  assign n43749 = ~n62836 & n62838;
  assign n43750 = x151 & x225;
  assign n43751 = n43749 & n43750;
  assign n43752 = n43749 | n43750;
  assign n43753 = ~n43751 & n43752;
  assign n62839 = n43438 & n43753;
  assign n62840 = (n43753 & n62660) | (n43753 & n62839) | (n62660 & n62839);
  assign n62841 = n43438 | n43753;
  assign n62842 = n62660 | n62841;
  assign n43756 = ~n62840 & n62842;
  assign n43757 = x150 & x226;
  assign n43758 = n43756 & n43757;
  assign n43759 = n43756 | n43757;
  assign n43760 = ~n43758 & n43759;
  assign n62843 = n43445 & n43760;
  assign n62844 = (n43760 & n62664) | (n43760 & n62843) | (n62664 & n62843);
  assign n62845 = n43445 | n43760;
  assign n62846 = n62664 | n62845;
  assign n43763 = ~n62844 & n62846;
  assign n43764 = x149 & x227;
  assign n43765 = n43763 & n43764;
  assign n43766 = n43763 | n43764;
  assign n43767 = ~n43765 & n43766;
  assign n62847 = n43452 & n43767;
  assign n62848 = (n43767 & n62668) | (n43767 & n62847) | (n62668 & n62847);
  assign n62849 = n43452 | n43767;
  assign n62850 = n62668 | n62849;
  assign n43770 = ~n62848 & n62850;
  assign n43771 = x148 & x228;
  assign n43772 = n43770 & n43771;
  assign n43773 = n43770 | n43771;
  assign n43774 = ~n43772 & n43773;
  assign n62851 = n43459 & n43774;
  assign n62852 = (n43774 & n62672) | (n43774 & n62851) | (n62672 & n62851);
  assign n62853 = n43459 | n43774;
  assign n62854 = n62672 | n62853;
  assign n43777 = ~n62852 & n62854;
  assign n43778 = x147 & x229;
  assign n43779 = n43777 & n43778;
  assign n43780 = n43777 | n43778;
  assign n43781 = ~n43779 & n43780;
  assign n62855 = n43466 & n43781;
  assign n62856 = (n43781 & n62676) | (n43781 & n62855) | (n62676 & n62855);
  assign n62857 = n43466 | n43781;
  assign n62858 = n62676 | n62857;
  assign n43784 = ~n62856 & n62858;
  assign n43785 = x146 & x230;
  assign n43786 = n43784 & n43785;
  assign n43787 = n43784 | n43785;
  assign n43788 = ~n43786 & n43787;
  assign n62859 = n43473 & n43788;
  assign n62860 = (n43788 & n62680) | (n43788 & n62859) | (n62680 & n62859);
  assign n62861 = n43473 | n43788;
  assign n62862 = n62680 | n62861;
  assign n43791 = ~n62860 & n62862;
  assign n43792 = x145 & x231;
  assign n43793 = n43791 & n43792;
  assign n43794 = n43791 | n43792;
  assign n43795 = ~n43793 & n43794;
  assign n62863 = n43480 & n43795;
  assign n62864 = (n43795 & n62684) | (n43795 & n62863) | (n62684 & n62863);
  assign n62865 = n43480 | n43795;
  assign n62866 = n62684 | n62865;
  assign n43798 = ~n62864 & n62866;
  assign n43799 = x144 & x232;
  assign n43800 = n43798 & n43799;
  assign n43801 = n43798 | n43799;
  assign n43802 = ~n43800 & n43801;
  assign n62867 = n43487 & n43802;
  assign n62868 = (n43802 & n62688) | (n43802 & n62867) | (n62688 & n62867);
  assign n62869 = n43487 | n43802;
  assign n62870 = n62688 | n62869;
  assign n43805 = ~n62868 & n62870;
  assign n43806 = x143 & x233;
  assign n43807 = n43805 & n43806;
  assign n43808 = n43805 | n43806;
  assign n43809 = ~n43807 & n43808;
  assign n62871 = n43494 & n43809;
  assign n62872 = (n43809 & n62692) | (n43809 & n62871) | (n62692 & n62871);
  assign n62873 = n43494 | n43809;
  assign n62874 = n62692 | n62873;
  assign n43812 = ~n62872 & n62874;
  assign n43813 = x142 & x234;
  assign n43814 = n43812 & n43813;
  assign n43815 = n43812 | n43813;
  assign n43816 = ~n43814 & n43815;
  assign n62875 = n43501 & n43816;
  assign n62876 = (n43816 & n62696) | (n43816 & n62875) | (n62696 & n62875);
  assign n62877 = n43501 | n43816;
  assign n62878 = n62696 | n62877;
  assign n43819 = ~n62876 & n62878;
  assign n43820 = x141 & x235;
  assign n43821 = n43819 & n43820;
  assign n43822 = n43819 | n43820;
  assign n43823 = ~n43821 & n43822;
  assign n62879 = n43508 & n43823;
  assign n62880 = (n43823 & n62700) | (n43823 & n62879) | (n62700 & n62879);
  assign n62881 = n43508 | n43823;
  assign n62882 = n62700 | n62881;
  assign n43826 = ~n62880 & n62882;
  assign n43827 = x140 & x236;
  assign n43828 = n43826 & n43827;
  assign n43829 = n43826 | n43827;
  assign n43830 = ~n43828 & n43829;
  assign n62883 = n43515 & n43830;
  assign n62884 = (n43830 & n62704) | (n43830 & n62883) | (n62704 & n62883);
  assign n62885 = n43515 | n43830;
  assign n62886 = n62704 | n62885;
  assign n43833 = ~n62884 & n62886;
  assign n43834 = x139 & x237;
  assign n43835 = n43833 & n43834;
  assign n43836 = n43833 | n43834;
  assign n43837 = ~n43835 & n43836;
  assign n62887 = n43522 & n43837;
  assign n62888 = (n43837 & n62708) | (n43837 & n62887) | (n62708 & n62887);
  assign n62889 = n43522 | n43837;
  assign n62890 = n62708 | n62889;
  assign n43840 = ~n62888 & n62890;
  assign n43841 = x138 & x238;
  assign n43842 = n43840 & n43841;
  assign n43843 = n43840 | n43841;
  assign n43844 = ~n43842 & n43843;
  assign n62891 = n43529 & n43844;
  assign n62892 = (n43844 & n62712) | (n43844 & n62891) | (n62712 & n62891);
  assign n62893 = n43529 | n43844;
  assign n62894 = n62712 | n62893;
  assign n43847 = ~n62892 & n62894;
  assign n43848 = x137 & x239;
  assign n43849 = n43847 & n43848;
  assign n43850 = n43847 | n43848;
  assign n43851 = ~n43849 & n43850;
  assign n62895 = n43536 & n43851;
  assign n62896 = (n43851 & n62716) | (n43851 & n62895) | (n62716 & n62895);
  assign n62897 = n43536 | n43851;
  assign n62898 = n62716 | n62897;
  assign n43854 = ~n62896 & n62898;
  assign n62721 = (n73317 & n73390) | (n73317 & n62720) | (n73390 & n62720);
  assign n62902 = n43674 | n43676;
  assign n73454 = n43361 | n43674;
  assign n73455 = (n43674 & n43676) | (n43674 & n73454) | (n43676 & n73454);
  assign n73456 = (n62614 & n62902) | (n62614 & n73455) | (n62902 & n73455);
  assign n73457 = (n62613 & n62902) | (n62613 & n73455) | (n62902 & n73455);
  assign n73458 = (n62356 & n73456) | (n62356 & n73457) | (n73456 & n73457);
  assign n62907 = n43653 | n43655;
  assign n73459 = n43340 | n43653;
  assign n73460 = (n43653 & n43655) | (n43653 & n73459) | (n43655 & n73459);
  assign n73461 = (n62604 & n62907) | (n62604 & n73460) | (n62907 & n73460);
  assign n73462 = (n62603 & n62907) | (n62603 & n73460) | (n62907 & n73460);
  assign n73463 = (n73264 & n73461) | (n73264 & n73462) | (n73461 & n73462);
  assign n43894 = x175 & x202;
  assign n62924 = n43894 & n73416;
  assign n62925 = (n43894 & n73425) | (n43894 & n62924) | (n73425 & n62924);
  assign n62926 = n43894 | n73416;
  assign n62927 = n73425 | n62926;
  assign n43897 = ~n62925 & n62927;
  assign n62922 = n43590 | n43592;
  assign n73470 = n43897 & n62922;
  assign n73468 = n43277 | n43590;
  assign n73469 = (n43590 & n43592) | (n43590 & n73468) | (n43592 & n73468);
  assign n73471 = n43897 & n73469;
  assign n73472 = (n62575 & n73470) | (n62575 & n73471) | (n73470 & n73471);
  assign n73473 = n43897 | n62922;
  assign n73474 = n43897 | n73469;
  assign n73475 = (n62575 & n73473) | (n62575 & n73474) | (n73473 & n73474);
  assign n43900 = ~n73472 & n73475;
  assign n43901 = x174 & x203;
  assign n43902 = n43900 & n43901;
  assign n43903 = n43900 | n43901;
  assign n43904 = ~n43902 & n43903;
  assign n62919 = n43597 | n43599;
  assign n62928 = n43904 & n62919;
  assign n62929 = n43597 & n43904;
  assign n62930 = (n73410 & n62928) | (n73410 & n62929) | (n62928 & n62929);
  assign n62931 = n43904 | n62919;
  assign n62932 = n43597 | n43904;
  assign n62933 = (n73410 & n62931) | (n73410 & n62932) | (n62931 & n62932);
  assign n43907 = ~n62930 & n62933;
  assign n43908 = x173 & x204;
  assign n43909 = n43907 & n43908;
  assign n43910 = n43907 | n43908;
  assign n43911 = ~n43909 & n43910;
  assign n62934 = n43604 & n43911;
  assign n73476 = (n43911 & n62764) | (n43911 & n62934) | (n62764 & n62934);
  assign n73477 = (n43911 & n62763) | (n43911 & n62934) | (n62763 & n62934);
  assign n73478 = (n62555 & n73476) | (n62555 & n73477) | (n73476 & n73477);
  assign n62936 = n43604 | n43911;
  assign n73479 = n62764 | n62936;
  assign n73480 = n62763 | n62936;
  assign n73481 = (n62555 & n73479) | (n62555 & n73480) | (n73479 & n73480);
  assign n43914 = ~n73478 & n73481;
  assign n43915 = x172 & x205;
  assign n43916 = n43914 & n43915;
  assign n43917 = n43914 | n43915;
  assign n43918 = ~n43916 & n43917;
  assign n62917 = n43611 | n43613;
  assign n73482 = n43918 & n62917;
  assign n73466 = n43298 | n43611;
  assign n73467 = (n43611 & n43613) | (n43611 & n73466) | (n43613 & n73466);
  assign n73483 = n43918 & n73467;
  assign n73484 = (n62585 & n73482) | (n62585 & n73483) | (n73482 & n73483);
  assign n73485 = n43918 | n62917;
  assign n73486 = n43918 | n73467;
  assign n73487 = (n62585 & n73485) | (n62585 & n73486) | (n73485 & n73486);
  assign n43921 = ~n73484 & n73487;
  assign n43922 = x171 & x206;
  assign n43923 = n43921 & n43922;
  assign n43924 = n43921 | n43922;
  assign n43925 = ~n43923 & n43924;
  assign n62914 = n43618 | n43620;
  assign n62938 = n43925 & n62914;
  assign n62939 = n43618 & n43925;
  assign n62940 = (n73405 & n62938) | (n73405 & n62939) | (n62938 & n62939);
  assign n62941 = n43925 | n62914;
  assign n62942 = n43618 | n43925;
  assign n62943 = (n73405 & n62941) | (n73405 & n62942) | (n62941 & n62942);
  assign n43928 = ~n62940 & n62943;
  assign n43929 = x170 & x207;
  assign n43930 = n43928 & n43929;
  assign n43931 = n43928 | n43929;
  assign n43932 = ~n43930 & n43931;
  assign n62944 = n43625 & n43932;
  assign n73488 = (n43932 & n62774) | (n43932 & n62944) | (n62774 & n62944);
  assign n73489 = (n43932 & n62773) | (n43932 & n62944) | (n62773 & n62944);
  assign n73490 = (n62550 & n73488) | (n62550 & n73489) | (n73488 & n73489);
  assign n62946 = n43625 | n43932;
  assign n73491 = n62774 | n62946;
  assign n73492 = n62773 | n62946;
  assign n73493 = (n62550 & n73491) | (n62550 & n73492) | (n73491 & n73492);
  assign n43935 = ~n73490 & n73493;
  assign n43936 = x169 & x208;
  assign n43937 = n43935 & n43936;
  assign n43938 = n43935 | n43936;
  assign n43939 = ~n43937 & n43938;
  assign n62912 = n43632 | n43634;
  assign n73494 = n43939 & n62912;
  assign n73464 = n43319 | n43632;
  assign n73465 = (n43632 & n43634) | (n43632 & n73464) | (n43634 & n73464);
  assign n73495 = n43939 & n73465;
  assign n73496 = (n62595 & n73494) | (n62595 & n73495) | (n73494 & n73495);
  assign n73497 = n43939 | n62912;
  assign n73498 = n43939 | n73465;
  assign n73499 = (n62595 & n73497) | (n62595 & n73498) | (n73497 & n73498);
  assign n43942 = ~n73496 & n73499;
  assign n43943 = x168 & x209;
  assign n43944 = n43942 & n43943;
  assign n43945 = n43942 | n43943;
  assign n43946 = ~n43944 & n43945;
  assign n62909 = n43639 | n43641;
  assign n62948 = n43946 & n62909;
  assign n62949 = n43639 & n43946;
  assign n62950 = (n73400 & n62948) | (n73400 & n62949) | (n62948 & n62949);
  assign n62951 = n43946 | n62909;
  assign n62952 = n43639 | n43946;
  assign n62953 = (n73400 & n62951) | (n73400 & n62952) | (n62951 & n62952);
  assign n43949 = ~n62950 & n62953;
  assign n43950 = x167 & x210;
  assign n43951 = n43949 & n43950;
  assign n43952 = n43949 | n43950;
  assign n43953 = ~n43951 & n43952;
  assign n62954 = n43646 & n43953;
  assign n73500 = (n43953 & n62784) | (n43953 & n62954) | (n62784 & n62954);
  assign n73501 = (n43953 & n62783) | (n43953 & n62954) | (n62783 & n62954);
  assign n73502 = (n73330 & n73500) | (n73330 & n73501) | (n73500 & n73501);
  assign n62956 = n43646 | n43953;
  assign n73503 = n62784 | n62956;
  assign n73504 = n62783 | n62956;
  assign n73505 = (n73330 & n73503) | (n73330 & n73504) | (n73503 & n73504);
  assign n43956 = ~n73502 & n73505;
  assign n43957 = x166 & x211;
  assign n43958 = n43956 & n43957;
  assign n43959 = n43956 | n43957;
  assign n43960 = ~n43958 & n43959;
  assign n43961 = n73463 & n43960;
  assign n43962 = n73463 | n43960;
  assign n43963 = ~n43961 & n43962;
  assign n43964 = x165 & x212;
  assign n43965 = n43963 & n43964;
  assign n43966 = n43963 | n43964;
  assign n43967 = ~n43965 & n43966;
  assign n62904 = n43660 | n43662;
  assign n62958 = n43967 & n62904;
  assign n62959 = n43660 & n43967;
  assign n62960 = (n73395 & n62958) | (n73395 & n62959) | (n62958 & n62959);
  assign n62961 = n43967 | n62904;
  assign n62962 = n43660 | n43967;
  assign n62963 = (n73395 & n62961) | (n73395 & n62962) | (n62961 & n62962);
  assign n43970 = ~n62960 & n62963;
  assign n43971 = x164 & x213;
  assign n43972 = n43970 & n43971;
  assign n43973 = n43970 | n43971;
  assign n43974 = ~n43972 & n43973;
  assign n62964 = n43667 & n43974;
  assign n73506 = (n43974 & n62794) | (n43974 & n62964) | (n62794 & n62964);
  assign n73507 = (n43974 & n62793) | (n43974 & n62964) | (n62793 & n62964);
  assign n73508 = (n73325 & n73506) | (n73325 & n73507) | (n73506 & n73507);
  assign n62966 = n43667 | n43974;
  assign n73509 = n62794 | n62966;
  assign n73510 = n62793 | n62966;
  assign n73511 = (n73325 & n73509) | (n73325 & n73510) | (n73509 & n73510);
  assign n43977 = ~n73508 & n73511;
  assign n43978 = x163 & x214;
  assign n43979 = n43977 & n43978;
  assign n43980 = n43977 | n43978;
  assign n43981 = ~n43979 & n43980;
  assign n43982 = n73458 & n43981;
  assign n43983 = n73458 | n43981;
  assign n43984 = ~n43982 & n43983;
  assign n43985 = x162 & x215;
  assign n43986 = n43984 & n43985;
  assign n43987 = n43984 | n43985;
  assign n43988 = ~n43986 & n43987;
  assign n62899 = n43681 | n43683;
  assign n62968 = n43988 & n62899;
  assign n62969 = n43681 & n43988;
  assign n62970 = (n62721 & n62968) | (n62721 & n62969) | (n62968 & n62969);
  assign n62971 = n43988 | n62899;
  assign n62972 = n43681 | n43988;
  assign n62973 = (n62721 & n62971) | (n62721 & n62972) | (n62971 & n62972);
  assign n43991 = ~n62970 & n62973;
  assign n43992 = x161 & x216;
  assign n43993 = n43991 & n43992;
  assign n43994 = n43991 | n43992;
  assign n43995 = ~n43993 & n43994;
  assign n62974 = n43688 & n43995;
  assign n62975 = (n43995 & n73450) | (n43995 & n62974) | (n73450 & n62974);
  assign n62976 = n43688 | n43995;
  assign n62977 = n73450 | n62976;
  assign n43998 = ~n62975 & n62977;
  assign n43999 = x160 & x217;
  assign n44000 = n43998 & n43999;
  assign n44001 = n43998 | n43999;
  assign n44002 = ~n44000 & n44001;
  assign n62978 = n43695 & n44002;
  assign n62979 = (n44002 & n62808) | (n44002 & n62978) | (n62808 & n62978);
  assign n62980 = n43695 | n44002;
  assign n62981 = n62808 | n62980;
  assign n44005 = ~n62979 & n62981;
  assign n44006 = x159 & x218;
  assign n44007 = n44005 & n44006;
  assign n44008 = n44005 | n44006;
  assign n44009 = ~n44007 & n44008;
  assign n62982 = n43702 & n44009;
  assign n62983 = (n44009 & n62812) | (n44009 & n62982) | (n62812 & n62982);
  assign n62984 = n43702 | n44009;
  assign n62985 = n62812 | n62984;
  assign n44012 = ~n62983 & n62985;
  assign n44013 = x158 & x219;
  assign n44014 = n44012 & n44013;
  assign n44015 = n44012 | n44013;
  assign n44016 = ~n44014 & n44015;
  assign n62986 = n43709 & n44016;
  assign n62987 = (n44016 & n62816) | (n44016 & n62986) | (n62816 & n62986);
  assign n62988 = n43709 | n44016;
  assign n62989 = n62816 | n62988;
  assign n44019 = ~n62987 & n62989;
  assign n44020 = x157 & x220;
  assign n44021 = n44019 & n44020;
  assign n44022 = n44019 | n44020;
  assign n44023 = ~n44021 & n44022;
  assign n62990 = n43716 & n44023;
  assign n62991 = (n44023 & n62820) | (n44023 & n62990) | (n62820 & n62990);
  assign n62992 = n43716 | n44023;
  assign n62993 = n62820 | n62992;
  assign n44026 = ~n62991 & n62993;
  assign n44027 = x156 & x221;
  assign n44028 = n44026 & n44027;
  assign n44029 = n44026 | n44027;
  assign n44030 = ~n44028 & n44029;
  assign n62994 = n43723 & n44030;
  assign n62995 = (n44030 & n62824) | (n44030 & n62994) | (n62824 & n62994);
  assign n62996 = n43723 | n44030;
  assign n62997 = n62824 | n62996;
  assign n44033 = ~n62995 & n62997;
  assign n44034 = x155 & x222;
  assign n44035 = n44033 & n44034;
  assign n44036 = n44033 | n44034;
  assign n44037 = ~n44035 & n44036;
  assign n62998 = n43730 & n44037;
  assign n62999 = (n44037 & n62828) | (n44037 & n62998) | (n62828 & n62998);
  assign n63000 = n43730 | n44037;
  assign n63001 = n62828 | n63000;
  assign n44040 = ~n62999 & n63001;
  assign n44041 = x154 & x223;
  assign n44042 = n44040 & n44041;
  assign n44043 = n44040 | n44041;
  assign n44044 = ~n44042 & n44043;
  assign n63002 = n43737 & n44044;
  assign n63003 = (n44044 & n62832) | (n44044 & n63002) | (n62832 & n63002);
  assign n63004 = n43737 | n44044;
  assign n63005 = n62832 | n63004;
  assign n44047 = ~n63003 & n63005;
  assign n44048 = x153 & x224;
  assign n44049 = n44047 & n44048;
  assign n44050 = n44047 | n44048;
  assign n44051 = ~n44049 & n44050;
  assign n63006 = n43744 & n44051;
  assign n63007 = (n44051 & n62836) | (n44051 & n63006) | (n62836 & n63006);
  assign n63008 = n43744 | n44051;
  assign n63009 = n62836 | n63008;
  assign n44054 = ~n63007 & n63009;
  assign n44055 = x152 & x225;
  assign n44056 = n44054 & n44055;
  assign n44057 = n44054 | n44055;
  assign n44058 = ~n44056 & n44057;
  assign n63010 = n43751 & n44058;
  assign n63011 = (n44058 & n62840) | (n44058 & n63010) | (n62840 & n63010);
  assign n63012 = n43751 | n44058;
  assign n63013 = n62840 | n63012;
  assign n44061 = ~n63011 & n63013;
  assign n44062 = x151 & x226;
  assign n44063 = n44061 & n44062;
  assign n44064 = n44061 | n44062;
  assign n44065 = ~n44063 & n44064;
  assign n63014 = n43758 & n44065;
  assign n63015 = (n44065 & n62844) | (n44065 & n63014) | (n62844 & n63014);
  assign n63016 = n43758 | n44065;
  assign n63017 = n62844 | n63016;
  assign n44068 = ~n63015 & n63017;
  assign n44069 = x150 & x227;
  assign n44070 = n44068 & n44069;
  assign n44071 = n44068 | n44069;
  assign n44072 = ~n44070 & n44071;
  assign n63018 = n43765 & n44072;
  assign n63019 = (n44072 & n62848) | (n44072 & n63018) | (n62848 & n63018);
  assign n63020 = n43765 | n44072;
  assign n63021 = n62848 | n63020;
  assign n44075 = ~n63019 & n63021;
  assign n44076 = x149 & x228;
  assign n44077 = n44075 & n44076;
  assign n44078 = n44075 | n44076;
  assign n44079 = ~n44077 & n44078;
  assign n63022 = n43772 & n44079;
  assign n63023 = (n44079 & n62852) | (n44079 & n63022) | (n62852 & n63022);
  assign n63024 = n43772 | n44079;
  assign n63025 = n62852 | n63024;
  assign n44082 = ~n63023 & n63025;
  assign n44083 = x148 & x229;
  assign n44084 = n44082 & n44083;
  assign n44085 = n44082 | n44083;
  assign n44086 = ~n44084 & n44085;
  assign n63026 = n43779 & n44086;
  assign n63027 = (n44086 & n62856) | (n44086 & n63026) | (n62856 & n63026);
  assign n63028 = n43779 | n44086;
  assign n63029 = n62856 | n63028;
  assign n44089 = ~n63027 & n63029;
  assign n44090 = x147 & x230;
  assign n44091 = n44089 & n44090;
  assign n44092 = n44089 | n44090;
  assign n44093 = ~n44091 & n44092;
  assign n63030 = n43786 & n44093;
  assign n63031 = (n44093 & n62860) | (n44093 & n63030) | (n62860 & n63030);
  assign n63032 = n43786 | n44093;
  assign n63033 = n62860 | n63032;
  assign n44096 = ~n63031 & n63033;
  assign n44097 = x146 & x231;
  assign n44098 = n44096 & n44097;
  assign n44099 = n44096 | n44097;
  assign n44100 = ~n44098 & n44099;
  assign n63034 = n43793 & n44100;
  assign n63035 = (n44100 & n62864) | (n44100 & n63034) | (n62864 & n63034);
  assign n63036 = n43793 | n44100;
  assign n63037 = n62864 | n63036;
  assign n44103 = ~n63035 & n63037;
  assign n44104 = x145 & x232;
  assign n44105 = n44103 & n44104;
  assign n44106 = n44103 | n44104;
  assign n44107 = ~n44105 & n44106;
  assign n63038 = n43800 & n44107;
  assign n63039 = (n44107 & n62868) | (n44107 & n63038) | (n62868 & n63038);
  assign n63040 = n43800 | n44107;
  assign n63041 = n62868 | n63040;
  assign n44110 = ~n63039 & n63041;
  assign n44111 = x144 & x233;
  assign n44112 = n44110 & n44111;
  assign n44113 = n44110 | n44111;
  assign n44114 = ~n44112 & n44113;
  assign n63042 = n43807 & n44114;
  assign n63043 = (n44114 & n62872) | (n44114 & n63042) | (n62872 & n63042);
  assign n63044 = n43807 | n44114;
  assign n63045 = n62872 | n63044;
  assign n44117 = ~n63043 & n63045;
  assign n44118 = x143 & x234;
  assign n44119 = n44117 & n44118;
  assign n44120 = n44117 | n44118;
  assign n44121 = ~n44119 & n44120;
  assign n63046 = n43814 & n44121;
  assign n63047 = (n44121 & n62876) | (n44121 & n63046) | (n62876 & n63046);
  assign n63048 = n43814 | n44121;
  assign n63049 = n62876 | n63048;
  assign n44124 = ~n63047 & n63049;
  assign n44125 = x142 & x235;
  assign n44126 = n44124 & n44125;
  assign n44127 = n44124 | n44125;
  assign n44128 = ~n44126 & n44127;
  assign n63050 = n43821 & n44128;
  assign n63051 = (n44128 & n62880) | (n44128 & n63050) | (n62880 & n63050);
  assign n63052 = n43821 | n44128;
  assign n63053 = n62880 | n63052;
  assign n44131 = ~n63051 & n63053;
  assign n44132 = x141 & x236;
  assign n44133 = n44131 & n44132;
  assign n44134 = n44131 | n44132;
  assign n44135 = ~n44133 & n44134;
  assign n63054 = n43828 & n44135;
  assign n63055 = (n44135 & n62884) | (n44135 & n63054) | (n62884 & n63054);
  assign n63056 = n43828 | n44135;
  assign n63057 = n62884 | n63056;
  assign n44138 = ~n63055 & n63057;
  assign n44139 = x140 & x237;
  assign n44140 = n44138 & n44139;
  assign n44141 = n44138 | n44139;
  assign n44142 = ~n44140 & n44141;
  assign n63058 = n43835 & n44142;
  assign n63059 = (n44142 & n62888) | (n44142 & n63058) | (n62888 & n63058);
  assign n63060 = n43835 | n44142;
  assign n63061 = n62888 | n63060;
  assign n44145 = ~n63059 & n63061;
  assign n44146 = x139 & x238;
  assign n44147 = n44145 & n44146;
  assign n44148 = n44145 | n44146;
  assign n44149 = ~n44147 & n44148;
  assign n63062 = n43842 & n44149;
  assign n63063 = (n44149 & n62892) | (n44149 & n63062) | (n62892 & n63062);
  assign n63064 = n43842 | n44149;
  assign n63065 = n62892 | n63064;
  assign n44152 = ~n63063 & n63065;
  assign n44153 = x138 & x239;
  assign n44154 = n44152 & n44153;
  assign n44155 = n44152 | n44153;
  assign n44156 = ~n44154 & n44155;
  assign n63066 = n43849 & n44156;
  assign n63067 = (n44156 & n62896) | (n44156 & n63066) | (n62896 & n63066);
  assign n63068 = n43849 | n44156;
  assign n63069 = n62896 | n63068;
  assign n44159 = ~n63067 & n63069;
  assign n63076 = n43972 | n43974;
  assign n73514 = n43667 | n43972;
  assign n73515 = (n43972 & n43974) | (n43972 & n73514) | (n43974 & n73514);
  assign n73516 = (n62794 & n63076) | (n62794 & n73515) | (n63076 & n73515);
  assign n73517 = (n62793 & n63076) | (n62793 & n73515) | (n63076 & n73515);
  assign n73518 = (n73325 & n73516) | (n73325 & n73517) | (n73516 & n73517);
  assign n63081 = n43951 | n43953;
  assign n73519 = n43646 | n43951;
  assign n73520 = (n43951 & n43953) | (n43951 & n73519) | (n43953 & n73519);
  assign n73521 = (n62784 & n63081) | (n62784 & n73520) | (n63081 & n73520);
  assign n73522 = (n62783 & n63081) | (n62783 & n73520) | (n63081 & n73520);
  assign n73523 = (n73330 & n73521) | (n73330 & n73522) | (n73521 & n73522);
  assign n62913 = (n62595 & n73465) | (n62595 & n62912) | (n73465 & n62912);
  assign n63086 = n43930 | n43932;
  assign n73524 = n43625 | n43930;
  assign n73525 = (n43930 & n43932) | (n43930 & n73524) | (n43932 & n73524);
  assign n73526 = (n62774 & n63086) | (n62774 & n73525) | (n63086 & n73525);
  assign n73527 = (n62773 & n63086) | (n62773 & n73525) | (n63086 & n73525);
  assign n73528 = (n62550 & n73526) | (n62550 & n73527) | (n73526 & n73527);
  assign n62918 = (n62585 & n73467) | (n62585 & n62917) | (n73467 & n62917);
  assign n63091 = n43909 | n43911;
  assign n73529 = n43604 | n43909;
  assign n73530 = (n43909 & n43911) | (n43909 & n73529) | (n43911 & n73529);
  assign n73531 = (n62764 & n63091) | (n62764 & n73530) | (n63091 & n73530);
  assign n73532 = (n62763 & n63091) | (n62763 & n73530) | (n63091 & n73530);
  assign n73533 = (n62555 & n73531) | (n62555 & n73532) | (n73531 & n73532);
  assign n44198 = x175 & x203;
  assign n73535 = n44198 & n62924;
  assign n73536 = n43894 & n44198;
  assign n73537 = (n73425 & n73535) | (n73425 & n73536) | (n73535 & n73536);
  assign n73534 = (n43897 & n44198) | (n43897 & n73537) | (n44198 & n73537);
  assign n73538 = (n62922 & n73534) | (n62922 & n73537) | (n73534 & n73537);
  assign n73539 = (n73469 & n73534) | (n73469 & n73537) | (n73534 & n73537);
  assign n73540 = (n62575 & n73538) | (n62575 & n73539) | (n73538 & n73539);
  assign n73542 = n44198 | n62924;
  assign n73543 = n43894 | n44198;
  assign n73544 = (n73425 & n73542) | (n73425 & n73543) | (n73542 & n73543);
  assign n73541 = n43897 | n73544;
  assign n73545 = (n62922 & n73541) | (n62922 & n73544) | (n73541 & n73544);
  assign n73546 = (n73469 & n73541) | (n73469 & n73544) | (n73541 & n73544);
  assign n73547 = (n62575 & n73545) | (n62575 & n73546) | (n73545 & n73546);
  assign n44201 = ~n73540 & n73547;
  assign n63101 = n43902 & n44201;
  assign n63102 = (n44201 & n62930) | (n44201 & n63101) | (n62930 & n63101);
  assign n63103 = n43902 | n44201;
  assign n63104 = n62930 | n63103;
  assign n44204 = ~n63102 & n63104;
  assign n44205 = x174 & x204;
  assign n44206 = n44204 & n44205;
  assign n44207 = n44204 | n44205;
  assign n44208 = ~n44206 & n44207;
  assign n44209 = n73533 & n44208;
  assign n44210 = n73533 | n44208;
  assign n44211 = ~n44209 & n44210;
  assign n44212 = x173 & x205;
  assign n44213 = n44211 & n44212;
  assign n44214 = n44211 | n44212;
  assign n44215 = ~n44213 & n44214;
  assign n63088 = n43916 | n43918;
  assign n63105 = n44215 & n63088;
  assign n63106 = n43916 & n44215;
  assign n63107 = (n62918 & n63105) | (n62918 & n63106) | (n63105 & n63106);
  assign n63108 = n44215 | n63088;
  assign n63109 = n43916 | n44215;
  assign n63110 = (n62918 & n63108) | (n62918 & n63109) | (n63108 & n63109);
  assign n44218 = ~n63107 & n63110;
  assign n44219 = x172 & x206;
  assign n44220 = n44218 & n44219;
  assign n44221 = n44218 | n44219;
  assign n44222 = ~n44220 & n44221;
  assign n63111 = n43923 & n44222;
  assign n63112 = (n44222 & n62940) | (n44222 & n63111) | (n62940 & n63111);
  assign n63113 = n43923 | n44222;
  assign n63114 = n62940 | n63113;
  assign n44225 = ~n63112 & n63114;
  assign n44226 = x171 & x207;
  assign n44227 = n44225 & n44226;
  assign n44228 = n44225 | n44226;
  assign n44229 = ~n44227 & n44228;
  assign n44230 = n73528 & n44229;
  assign n44231 = n73528 | n44229;
  assign n44232 = ~n44230 & n44231;
  assign n44233 = x170 & x208;
  assign n44234 = n44232 & n44233;
  assign n44235 = n44232 | n44233;
  assign n44236 = ~n44234 & n44235;
  assign n63083 = n43937 | n43939;
  assign n63115 = n44236 & n63083;
  assign n63116 = n43937 & n44236;
  assign n63117 = (n62913 & n63115) | (n62913 & n63116) | (n63115 & n63116);
  assign n63118 = n44236 | n63083;
  assign n63119 = n43937 | n44236;
  assign n63120 = (n62913 & n63118) | (n62913 & n63119) | (n63118 & n63119);
  assign n44239 = ~n63117 & n63120;
  assign n44240 = x169 & x209;
  assign n44241 = n44239 & n44240;
  assign n44242 = n44239 | n44240;
  assign n44243 = ~n44241 & n44242;
  assign n63121 = n43944 & n44243;
  assign n63122 = (n44243 & n62950) | (n44243 & n63121) | (n62950 & n63121);
  assign n63123 = n43944 | n44243;
  assign n63124 = n62950 | n63123;
  assign n44246 = ~n63122 & n63124;
  assign n44247 = x168 & x210;
  assign n44248 = n44246 & n44247;
  assign n44249 = n44246 | n44247;
  assign n44250 = ~n44248 & n44249;
  assign n44251 = n73523 & n44250;
  assign n44252 = n73523 | n44250;
  assign n44253 = ~n44251 & n44252;
  assign n44254 = x167 & x211;
  assign n44255 = n44253 & n44254;
  assign n44256 = n44253 | n44254;
  assign n44257 = ~n44255 & n44256;
  assign n63078 = n43958 | n43960;
  assign n63125 = n44257 & n63078;
  assign n63126 = n43958 & n44257;
  assign n63127 = (n73463 & n63125) | (n73463 & n63126) | (n63125 & n63126);
  assign n63128 = n44257 | n63078;
  assign n63129 = n43958 | n44257;
  assign n63130 = (n73463 & n63128) | (n73463 & n63129) | (n63128 & n63129);
  assign n44260 = ~n63127 & n63130;
  assign n44261 = x166 & x212;
  assign n44262 = n44260 & n44261;
  assign n44263 = n44260 | n44261;
  assign n44264 = ~n44262 & n44263;
  assign n63131 = n43965 & n44264;
  assign n73548 = (n44264 & n62959) | (n44264 & n63131) | (n62959 & n63131);
  assign n73549 = (n44264 & n62958) | (n44264 & n63131) | (n62958 & n63131);
  assign n73550 = (n73395 & n73548) | (n73395 & n73549) | (n73548 & n73549);
  assign n63133 = n43965 | n44264;
  assign n73551 = n62959 | n63133;
  assign n73552 = n62958 | n63133;
  assign n73553 = (n73395 & n73551) | (n73395 & n73552) | (n73551 & n73552);
  assign n44267 = ~n73550 & n73553;
  assign n44268 = x165 & x213;
  assign n44269 = n44267 & n44268;
  assign n44270 = n44267 | n44268;
  assign n44271 = ~n44269 & n44270;
  assign n44272 = n73518 & n44271;
  assign n44273 = n73518 | n44271;
  assign n44274 = ~n44272 & n44273;
  assign n44275 = x164 & x214;
  assign n44276 = n44274 & n44275;
  assign n44277 = n44274 | n44275;
  assign n44278 = ~n44276 & n44277;
  assign n63073 = n43979 | n43981;
  assign n63135 = n44278 & n63073;
  assign n63136 = n43979 & n44278;
  assign n63137 = (n73458 & n63135) | (n73458 & n63136) | (n63135 & n63136);
  assign n63138 = n44278 | n63073;
  assign n63139 = n43979 | n44278;
  assign n63140 = (n73458 & n63138) | (n73458 & n63139) | (n63138 & n63139);
  assign n44281 = ~n63137 & n63140;
  assign n44282 = x163 & x215;
  assign n44283 = n44281 & n44282;
  assign n44284 = n44281 | n44282;
  assign n44285 = ~n44283 & n44284;
  assign n63141 = n43986 & n44285;
  assign n73554 = (n44285 & n62969) | (n44285 & n63141) | (n62969 & n63141);
  assign n73555 = (n44285 & n62968) | (n44285 & n63141) | (n62968 & n63141);
  assign n73556 = (n62721 & n73554) | (n62721 & n73555) | (n73554 & n73555);
  assign n63143 = n43986 | n44285;
  assign n73557 = n62969 | n63143;
  assign n73558 = n62968 | n63143;
  assign n73559 = (n62721 & n73557) | (n62721 & n73558) | (n73557 & n73558);
  assign n44288 = ~n73556 & n73559;
  assign n44289 = x162 & x216;
  assign n44290 = n44288 & n44289;
  assign n44291 = n44288 | n44289;
  assign n44292 = ~n44290 & n44291;
  assign n63071 = n43993 | n43995;
  assign n73560 = n44292 & n63071;
  assign n73512 = n43688 | n43993;
  assign n73513 = (n43993 & n43995) | (n43993 & n73512) | (n43995 & n73512);
  assign n73561 = n44292 & n73513;
  assign n73562 = (n73450 & n73560) | (n73450 & n73561) | (n73560 & n73561);
  assign n73563 = n44292 | n63071;
  assign n73564 = n44292 | n73513;
  assign n73565 = (n73450 & n73563) | (n73450 & n73564) | (n73563 & n73564);
  assign n44295 = ~n73562 & n73565;
  assign n44296 = x161 & x217;
  assign n44297 = n44295 & n44296;
  assign n44298 = n44295 | n44296;
  assign n44299 = ~n44297 & n44298;
  assign n63145 = n44000 & n44299;
  assign n73566 = (n44299 & n62978) | (n44299 & n63145) | (n62978 & n63145);
  assign n73567 = (n44002 & n44299) | (n44002 & n63145) | (n44299 & n63145);
  assign n73568 = (n62808 & n73566) | (n62808 & n73567) | (n73566 & n73567);
  assign n63147 = n44000 | n44299;
  assign n73569 = n62978 | n63147;
  assign n73570 = n44002 | n63147;
  assign n73571 = (n62808 & n73569) | (n62808 & n73570) | (n73569 & n73570);
  assign n44302 = ~n73568 & n73571;
  assign n44303 = x160 & x218;
  assign n44304 = n44302 & n44303;
  assign n44305 = n44302 | n44303;
  assign n44306 = ~n44304 & n44305;
  assign n63149 = n44007 & n44306;
  assign n63150 = (n44306 & n62983) | (n44306 & n63149) | (n62983 & n63149);
  assign n63151 = n44007 | n44306;
  assign n63152 = n62983 | n63151;
  assign n44309 = ~n63150 & n63152;
  assign n44310 = x159 & x219;
  assign n44311 = n44309 & n44310;
  assign n44312 = n44309 | n44310;
  assign n44313 = ~n44311 & n44312;
  assign n63153 = n44014 & n44313;
  assign n63154 = (n44313 & n62987) | (n44313 & n63153) | (n62987 & n63153);
  assign n63155 = n44014 | n44313;
  assign n63156 = n62987 | n63155;
  assign n44316 = ~n63154 & n63156;
  assign n44317 = x158 & x220;
  assign n44318 = n44316 & n44317;
  assign n44319 = n44316 | n44317;
  assign n44320 = ~n44318 & n44319;
  assign n63157 = n44021 & n44320;
  assign n63158 = (n44320 & n62991) | (n44320 & n63157) | (n62991 & n63157);
  assign n63159 = n44021 | n44320;
  assign n63160 = n62991 | n63159;
  assign n44323 = ~n63158 & n63160;
  assign n44324 = x157 & x221;
  assign n44325 = n44323 & n44324;
  assign n44326 = n44323 | n44324;
  assign n44327 = ~n44325 & n44326;
  assign n63161 = n44028 & n44327;
  assign n63162 = (n44327 & n62995) | (n44327 & n63161) | (n62995 & n63161);
  assign n63163 = n44028 | n44327;
  assign n63164 = n62995 | n63163;
  assign n44330 = ~n63162 & n63164;
  assign n44331 = x156 & x222;
  assign n44332 = n44330 & n44331;
  assign n44333 = n44330 | n44331;
  assign n44334 = ~n44332 & n44333;
  assign n63165 = n44035 & n44334;
  assign n63166 = (n44334 & n62999) | (n44334 & n63165) | (n62999 & n63165);
  assign n63167 = n44035 | n44334;
  assign n63168 = n62999 | n63167;
  assign n44337 = ~n63166 & n63168;
  assign n44338 = x155 & x223;
  assign n44339 = n44337 & n44338;
  assign n44340 = n44337 | n44338;
  assign n44341 = ~n44339 & n44340;
  assign n63169 = n44042 & n44341;
  assign n63170 = (n44341 & n63003) | (n44341 & n63169) | (n63003 & n63169);
  assign n63171 = n44042 | n44341;
  assign n63172 = n63003 | n63171;
  assign n44344 = ~n63170 & n63172;
  assign n44345 = x154 & x224;
  assign n44346 = n44344 & n44345;
  assign n44347 = n44344 | n44345;
  assign n44348 = ~n44346 & n44347;
  assign n63173 = n44049 & n44348;
  assign n63174 = (n44348 & n63007) | (n44348 & n63173) | (n63007 & n63173);
  assign n63175 = n44049 | n44348;
  assign n63176 = n63007 | n63175;
  assign n44351 = ~n63174 & n63176;
  assign n44352 = x153 & x225;
  assign n44353 = n44351 & n44352;
  assign n44354 = n44351 | n44352;
  assign n44355 = ~n44353 & n44354;
  assign n63177 = n44056 & n44355;
  assign n63178 = (n44355 & n63011) | (n44355 & n63177) | (n63011 & n63177);
  assign n63179 = n44056 | n44355;
  assign n63180 = n63011 | n63179;
  assign n44358 = ~n63178 & n63180;
  assign n44359 = x152 & x226;
  assign n44360 = n44358 & n44359;
  assign n44361 = n44358 | n44359;
  assign n44362 = ~n44360 & n44361;
  assign n63181 = n44063 & n44362;
  assign n63182 = (n44362 & n63015) | (n44362 & n63181) | (n63015 & n63181);
  assign n63183 = n44063 | n44362;
  assign n63184 = n63015 | n63183;
  assign n44365 = ~n63182 & n63184;
  assign n44366 = x151 & x227;
  assign n44367 = n44365 & n44366;
  assign n44368 = n44365 | n44366;
  assign n44369 = ~n44367 & n44368;
  assign n63185 = n44070 & n44369;
  assign n63186 = (n44369 & n63019) | (n44369 & n63185) | (n63019 & n63185);
  assign n63187 = n44070 | n44369;
  assign n63188 = n63019 | n63187;
  assign n44372 = ~n63186 & n63188;
  assign n44373 = x150 & x228;
  assign n44374 = n44372 & n44373;
  assign n44375 = n44372 | n44373;
  assign n44376 = ~n44374 & n44375;
  assign n63189 = n44077 & n44376;
  assign n63190 = (n44376 & n63023) | (n44376 & n63189) | (n63023 & n63189);
  assign n63191 = n44077 | n44376;
  assign n63192 = n63023 | n63191;
  assign n44379 = ~n63190 & n63192;
  assign n44380 = x149 & x229;
  assign n44381 = n44379 & n44380;
  assign n44382 = n44379 | n44380;
  assign n44383 = ~n44381 & n44382;
  assign n63193 = n44084 & n44383;
  assign n63194 = (n44383 & n63027) | (n44383 & n63193) | (n63027 & n63193);
  assign n63195 = n44084 | n44383;
  assign n63196 = n63027 | n63195;
  assign n44386 = ~n63194 & n63196;
  assign n44387 = x148 & x230;
  assign n44388 = n44386 & n44387;
  assign n44389 = n44386 | n44387;
  assign n44390 = ~n44388 & n44389;
  assign n63197 = n44091 & n44390;
  assign n63198 = (n44390 & n63031) | (n44390 & n63197) | (n63031 & n63197);
  assign n63199 = n44091 | n44390;
  assign n63200 = n63031 | n63199;
  assign n44393 = ~n63198 & n63200;
  assign n44394 = x147 & x231;
  assign n44395 = n44393 & n44394;
  assign n44396 = n44393 | n44394;
  assign n44397 = ~n44395 & n44396;
  assign n63201 = n44098 & n44397;
  assign n63202 = (n44397 & n63035) | (n44397 & n63201) | (n63035 & n63201);
  assign n63203 = n44098 | n44397;
  assign n63204 = n63035 | n63203;
  assign n44400 = ~n63202 & n63204;
  assign n44401 = x146 & x232;
  assign n44402 = n44400 & n44401;
  assign n44403 = n44400 | n44401;
  assign n44404 = ~n44402 & n44403;
  assign n63205 = n44105 & n44404;
  assign n63206 = (n44404 & n63039) | (n44404 & n63205) | (n63039 & n63205);
  assign n63207 = n44105 | n44404;
  assign n63208 = n63039 | n63207;
  assign n44407 = ~n63206 & n63208;
  assign n44408 = x145 & x233;
  assign n44409 = n44407 & n44408;
  assign n44410 = n44407 | n44408;
  assign n44411 = ~n44409 & n44410;
  assign n63209 = n44112 & n44411;
  assign n63210 = (n44411 & n63043) | (n44411 & n63209) | (n63043 & n63209);
  assign n63211 = n44112 | n44411;
  assign n63212 = n63043 | n63211;
  assign n44414 = ~n63210 & n63212;
  assign n44415 = x144 & x234;
  assign n44416 = n44414 & n44415;
  assign n44417 = n44414 | n44415;
  assign n44418 = ~n44416 & n44417;
  assign n63213 = n44119 & n44418;
  assign n63214 = (n44418 & n63047) | (n44418 & n63213) | (n63047 & n63213);
  assign n63215 = n44119 | n44418;
  assign n63216 = n63047 | n63215;
  assign n44421 = ~n63214 & n63216;
  assign n44422 = x143 & x235;
  assign n44423 = n44421 & n44422;
  assign n44424 = n44421 | n44422;
  assign n44425 = ~n44423 & n44424;
  assign n63217 = n44126 & n44425;
  assign n63218 = (n44425 & n63051) | (n44425 & n63217) | (n63051 & n63217);
  assign n63219 = n44126 | n44425;
  assign n63220 = n63051 | n63219;
  assign n44428 = ~n63218 & n63220;
  assign n44429 = x142 & x236;
  assign n44430 = n44428 & n44429;
  assign n44431 = n44428 | n44429;
  assign n44432 = ~n44430 & n44431;
  assign n63221 = n44133 & n44432;
  assign n63222 = (n44432 & n63055) | (n44432 & n63221) | (n63055 & n63221);
  assign n63223 = n44133 | n44432;
  assign n63224 = n63055 | n63223;
  assign n44435 = ~n63222 & n63224;
  assign n44436 = x141 & x237;
  assign n44437 = n44435 & n44436;
  assign n44438 = n44435 | n44436;
  assign n44439 = ~n44437 & n44438;
  assign n63225 = n44140 & n44439;
  assign n63226 = (n44439 & n63059) | (n44439 & n63225) | (n63059 & n63225);
  assign n63227 = n44140 | n44439;
  assign n63228 = n63059 | n63227;
  assign n44442 = ~n63226 & n63228;
  assign n44443 = x140 & x238;
  assign n44444 = n44442 & n44443;
  assign n44445 = n44442 | n44443;
  assign n44446 = ~n44444 & n44445;
  assign n63229 = n44147 & n44446;
  assign n63230 = (n44446 & n63063) | (n44446 & n63229) | (n63063 & n63229);
  assign n63231 = n44147 | n44446;
  assign n63232 = n63063 | n63231;
  assign n44449 = ~n63230 & n63232;
  assign n44450 = x139 & x239;
  assign n44451 = n44449 & n44450;
  assign n44452 = n44449 | n44450;
  assign n44453 = ~n44451 & n44452;
  assign n63233 = n44154 & n44453;
  assign n63234 = (n44453 & n63067) | (n44453 & n63233) | (n63067 & n63233);
  assign n63235 = n44154 | n44453;
  assign n63236 = n63067 | n63235;
  assign n44456 = ~n63234 & n63236;
  assign n63072 = (n73450 & n73513) | (n73450 & n63071) | (n73513 & n63071);
  assign n63240 = n44283 | n44285;
  assign n73572 = n43986 | n44283;
  assign n73573 = (n44283 & n44285) | (n44283 & n73572) | (n44285 & n73572);
  assign n73574 = (n62969 & n63240) | (n62969 & n73573) | (n63240 & n73573);
  assign n73575 = (n62968 & n63240) | (n62968 & n73573) | (n63240 & n73573);
  assign n73576 = (n62721 & n73574) | (n62721 & n73575) | (n73574 & n73575);
  assign n63245 = n44262 | n44264;
  assign n73577 = n43965 | n44262;
  assign n73578 = (n44262 & n44264) | (n44262 & n73577) | (n44264 & n73577);
  assign n73579 = (n62959 & n63245) | (n62959 & n73578) | (n63245 & n73578);
  assign n73580 = (n62958 & n63245) | (n62958 & n73578) | (n63245 & n73578);
  assign n73581 = (n73395 & n73579) | (n73395 & n73580) | (n73579 & n73580);
  assign n44494 = x175 & x204;
  assign n73586 = n44201 | n73540;
  assign n73587 = (n43902 & n73540) | (n43902 & n73586) | (n73540 & n73586);
  assign n63262 = n44494 & n73587;
  assign n73588 = n44494 & n73540;
  assign n73589 = (n44201 & n44494) | (n44201 & n73588) | (n44494 & n73588);
  assign n63264 = (n62930 & n63262) | (n62930 & n73589) | (n63262 & n73589);
  assign n63265 = n44494 | n73587;
  assign n73590 = n44494 | n73540;
  assign n73591 = n44201 | n73590;
  assign n63267 = (n62930 & n63265) | (n62930 & n73591) | (n63265 & n73591);
  assign n44497 = ~n63264 & n63267;
  assign n63269 = n44206 & n44497;
  assign n73592 = (n44208 & n44497) | (n44208 & n63269) | (n44497 & n63269);
  assign n63270 = (n73533 & n73592) | (n73533 & n63269) | (n73592 & n63269);
  assign n63272 = n44206 | n44497;
  assign n73593 = n44208 | n63272;
  assign n63273 = (n73533 & n73593) | (n73533 & n63272) | (n73593 & n63272);
  assign n44500 = ~n63270 & n63273;
  assign n44501 = x174 & x205;
  assign n44502 = n44500 & n44501;
  assign n44503 = n44500 | n44501;
  assign n44504 = ~n44502 & n44503;
  assign n63274 = n44213 & n44504;
  assign n73594 = (n44504 & n63106) | (n44504 & n63274) | (n63106 & n63274);
  assign n73595 = (n44504 & n63105) | (n44504 & n63274) | (n63105 & n63274);
  assign n73596 = (n62918 & n73594) | (n62918 & n73595) | (n73594 & n73595);
  assign n63276 = n44213 | n44504;
  assign n73597 = n63106 | n63276;
  assign n73598 = n63105 | n63276;
  assign n73599 = (n62918 & n73597) | (n62918 & n73598) | (n73597 & n73598);
  assign n44507 = ~n73596 & n73599;
  assign n44508 = x173 & x206;
  assign n44509 = n44507 & n44508;
  assign n44510 = n44507 | n44508;
  assign n44511 = ~n44509 & n44510;
  assign n63255 = n44220 | n44222;
  assign n73600 = n44511 & n63255;
  assign n73584 = n43923 | n44220;
  assign n73585 = (n44220 & n44222) | (n44220 & n73584) | (n44222 & n73584);
  assign n73601 = n44511 & n73585;
  assign n73602 = (n62940 & n73600) | (n62940 & n73601) | (n73600 & n73601);
  assign n73603 = n44511 | n63255;
  assign n73604 = n44511 | n73585;
  assign n73605 = (n62940 & n73603) | (n62940 & n73604) | (n73603 & n73604);
  assign n44514 = ~n73602 & n73605;
  assign n44515 = x172 & x207;
  assign n44516 = n44514 & n44515;
  assign n44517 = n44514 | n44515;
  assign n44518 = ~n44516 & n44517;
  assign n63252 = n44227 | n44229;
  assign n63278 = n44518 & n63252;
  assign n63279 = n44227 & n44518;
  assign n63280 = (n73528 & n63278) | (n73528 & n63279) | (n63278 & n63279);
  assign n63281 = n44518 | n63252;
  assign n63282 = n44227 | n44518;
  assign n63283 = (n73528 & n63281) | (n73528 & n63282) | (n63281 & n63282);
  assign n44521 = ~n63280 & n63283;
  assign n44522 = x171 & x208;
  assign n44523 = n44521 & n44522;
  assign n44524 = n44521 | n44522;
  assign n44525 = ~n44523 & n44524;
  assign n63284 = n44234 & n44525;
  assign n73606 = (n44525 & n63116) | (n44525 & n63284) | (n63116 & n63284);
  assign n73607 = (n44525 & n63115) | (n44525 & n63284) | (n63115 & n63284);
  assign n73608 = (n62913 & n73606) | (n62913 & n73607) | (n73606 & n73607);
  assign n63286 = n44234 | n44525;
  assign n73609 = n63116 | n63286;
  assign n73610 = n63115 | n63286;
  assign n73611 = (n62913 & n73609) | (n62913 & n73610) | (n73609 & n73610);
  assign n44528 = ~n73608 & n73611;
  assign n44529 = x170 & x209;
  assign n44530 = n44528 & n44529;
  assign n44531 = n44528 | n44529;
  assign n44532 = ~n44530 & n44531;
  assign n63250 = n44241 | n44243;
  assign n73612 = n44532 & n63250;
  assign n73582 = n43944 | n44241;
  assign n73583 = (n44241 & n44243) | (n44241 & n73582) | (n44243 & n73582);
  assign n73613 = n44532 & n73583;
  assign n73614 = (n62950 & n73612) | (n62950 & n73613) | (n73612 & n73613);
  assign n73615 = n44532 | n63250;
  assign n73616 = n44532 | n73583;
  assign n73617 = (n62950 & n73615) | (n62950 & n73616) | (n73615 & n73616);
  assign n44535 = ~n73614 & n73617;
  assign n44536 = x169 & x210;
  assign n44537 = n44535 & n44536;
  assign n44538 = n44535 | n44536;
  assign n44539 = ~n44537 & n44538;
  assign n63247 = n44248 | n44250;
  assign n63288 = n44539 & n63247;
  assign n63289 = n44248 & n44539;
  assign n63290 = (n73523 & n63288) | (n73523 & n63289) | (n63288 & n63289);
  assign n63291 = n44539 | n63247;
  assign n63292 = n44248 | n44539;
  assign n63293 = (n73523 & n63291) | (n73523 & n63292) | (n63291 & n63292);
  assign n44542 = ~n63290 & n63293;
  assign n44543 = x168 & x211;
  assign n44544 = n44542 & n44543;
  assign n44545 = n44542 | n44543;
  assign n44546 = ~n44544 & n44545;
  assign n63294 = n44255 & n44546;
  assign n73618 = (n44546 & n63126) | (n44546 & n63294) | (n63126 & n63294);
  assign n73619 = (n44546 & n63125) | (n44546 & n63294) | (n63125 & n63294);
  assign n73620 = (n73463 & n73618) | (n73463 & n73619) | (n73618 & n73619);
  assign n63296 = n44255 | n44546;
  assign n73621 = n63126 | n63296;
  assign n73622 = n63125 | n63296;
  assign n73623 = (n73463 & n73621) | (n73463 & n73622) | (n73621 & n73622);
  assign n44549 = ~n73620 & n73623;
  assign n44550 = x167 & x212;
  assign n44551 = n44549 & n44550;
  assign n44552 = n44549 | n44550;
  assign n44553 = ~n44551 & n44552;
  assign n44554 = n73581 & n44553;
  assign n44555 = n73581 | n44553;
  assign n44556 = ~n44554 & n44555;
  assign n44557 = x166 & x213;
  assign n44558 = n44556 & n44557;
  assign n44559 = n44556 | n44557;
  assign n44560 = ~n44558 & n44559;
  assign n63242 = n44269 | n44271;
  assign n63298 = n44560 & n63242;
  assign n63299 = n44269 & n44560;
  assign n63300 = (n73518 & n63298) | (n73518 & n63299) | (n63298 & n63299);
  assign n63301 = n44560 | n63242;
  assign n63302 = n44269 | n44560;
  assign n63303 = (n73518 & n63301) | (n73518 & n63302) | (n63301 & n63302);
  assign n44563 = ~n63300 & n63303;
  assign n44564 = x165 & x214;
  assign n44565 = n44563 & n44564;
  assign n44566 = n44563 | n44564;
  assign n44567 = ~n44565 & n44566;
  assign n63304 = n44276 & n44567;
  assign n73624 = (n44567 & n63136) | (n44567 & n63304) | (n63136 & n63304);
  assign n73625 = (n44567 & n63135) | (n44567 & n63304) | (n63135 & n63304);
  assign n73626 = (n73458 & n73624) | (n73458 & n73625) | (n73624 & n73625);
  assign n63306 = n44276 | n44567;
  assign n73627 = n63136 | n63306;
  assign n73628 = n63135 | n63306;
  assign n73629 = (n73458 & n73627) | (n73458 & n73628) | (n73627 & n73628);
  assign n44570 = ~n73626 & n73629;
  assign n44571 = x164 & x215;
  assign n44572 = n44570 & n44571;
  assign n44573 = n44570 | n44571;
  assign n44574 = ~n44572 & n44573;
  assign n44575 = n73576 & n44574;
  assign n44576 = n73576 | n44574;
  assign n44577 = ~n44575 & n44576;
  assign n44578 = x163 & x216;
  assign n44579 = n44577 & n44578;
  assign n44580 = n44577 | n44578;
  assign n44581 = ~n44579 & n44580;
  assign n63237 = n44290 | n44292;
  assign n63308 = n44581 & n63237;
  assign n63309 = n44290 & n44581;
  assign n63310 = (n63072 & n63308) | (n63072 & n63309) | (n63308 & n63309);
  assign n63311 = n44581 | n63237;
  assign n63312 = n44290 | n44581;
  assign n63313 = (n63072 & n63311) | (n63072 & n63312) | (n63311 & n63312);
  assign n44584 = ~n63310 & n63313;
  assign n44585 = x162 & x217;
  assign n44586 = n44584 & n44585;
  assign n44587 = n44584 | n44585;
  assign n44588 = ~n44586 & n44587;
  assign n63314 = n44297 & n44588;
  assign n63315 = (n44588 & n73568) | (n44588 & n63314) | (n73568 & n63314);
  assign n63316 = n44297 | n44588;
  assign n63317 = n73568 | n63316;
  assign n44591 = ~n63315 & n63317;
  assign n44592 = x161 & x218;
  assign n44593 = n44591 & n44592;
  assign n44594 = n44591 | n44592;
  assign n44595 = ~n44593 & n44594;
  assign n63318 = n44304 & n44595;
  assign n63319 = (n44595 & n63150) | (n44595 & n63318) | (n63150 & n63318);
  assign n63320 = n44304 | n44595;
  assign n63321 = n63150 | n63320;
  assign n44598 = ~n63319 & n63321;
  assign n44599 = x160 & x219;
  assign n44600 = n44598 & n44599;
  assign n44601 = n44598 | n44599;
  assign n44602 = ~n44600 & n44601;
  assign n63322 = n44311 & n44602;
  assign n63323 = (n44602 & n63154) | (n44602 & n63322) | (n63154 & n63322);
  assign n63324 = n44311 | n44602;
  assign n63325 = n63154 | n63324;
  assign n44605 = ~n63323 & n63325;
  assign n44606 = x159 & x220;
  assign n44607 = n44605 & n44606;
  assign n44608 = n44605 | n44606;
  assign n44609 = ~n44607 & n44608;
  assign n63326 = n44318 & n44609;
  assign n63327 = (n44609 & n63158) | (n44609 & n63326) | (n63158 & n63326);
  assign n63328 = n44318 | n44609;
  assign n63329 = n63158 | n63328;
  assign n44612 = ~n63327 & n63329;
  assign n44613 = x158 & x221;
  assign n44614 = n44612 & n44613;
  assign n44615 = n44612 | n44613;
  assign n44616 = ~n44614 & n44615;
  assign n63330 = n44325 & n44616;
  assign n63331 = (n44616 & n63162) | (n44616 & n63330) | (n63162 & n63330);
  assign n63332 = n44325 | n44616;
  assign n63333 = n63162 | n63332;
  assign n44619 = ~n63331 & n63333;
  assign n44620 = x157 & x222;
  assign n44621 = n44619 & n44620;
  assign n44622 = n44619 | n44620;
  assign n44623 = ~n44621 & n44622;
  assign n63334 = n44332 & n44623;
  assign n63335 = (n44623 & n63166) | (n44623 & n63334) | (n63166 & n63334);
  assign n63336 = n44332 | n44623;
  assign n63337 = n63166 | n63336;
  assign n44626 = ~n63335 & n63337;
  assign n44627 = x156 & x223;
  assign n44628 = n44626 & n44627;
  assign n44629 = n44626 | n44627;
  assign n44630 = ~n44628 & n44629;
  assign n63338 = n44339 & n44630;
  assign n63339 = (n44630 & n63170) | (n44630 & n63338) | (n63170 & n63338);
  assign n63340 = n44339 | n44630;
  assign n63341 = n63170 | n63340;
  assign n44633 = ~n63339 & n63341;
  assign n44634 = x155 & x224;
  assign n44635 = n44633 & n44634;
  assign n44636 = n44633 | n44634;
  assign n44637 = ~n44635 & n44636;
  assign n63342 = n44346 & n44637;
  assign n63343 = (n44637 & n63174) | (n44637 & n63342) | (n63174 & n63342);
  assign n63344 = n44346 | n44637;
  assign n63345 = n63174 | n63344;
  assign n44640 = ~n63343 & n63345;
  assign n44641 = x154 & x225;
  assign n44642 = n44640 & n44641;
  assign n44643 = n44640 | n44641;
  assign n44644 = ~n44642 & n44643;
  assign n63346 = n44353 & n44644;
  assign n63347 = (n44644 & n63178) | (n44644 & n63346) | (n63178 & n63346);
  assign n63348 = n44353 | n44644;
  assign n63349 = n63178 | n63348;
  assign n44647 = ~n63347 & n63349;
  assign n44648 = x153 & x226;
  assign n44649 = n44647 & n44648;
  assign n44650 = n44647 | n44648;
  assign n44651 = ~n44649 & n44650;
  assign n63350 = n44360 & n44651;
  assign n63351 = (n44651 & n63182) | (n44651 & n63350) | (n63182 & n63350);
  assign n63352 = n44360 | n44651;
  assign n63353 = n63182 | n63352;
  assign n44654 = ~n63351 & n63353;
  assign n44655 = x152 & x227;
  assign n44656 = n44654 & n44655;
  assign n44657 = n44654 | n44655;
  assign n44658 = ~n44656 & n44657;
  assign n63354 = n44367 & n44658;
  assign n63355 = (n44658 & n63186) | (n44658 & n63354) | (n63186 & n63354);
  assign n63356 = n44367 | n44658;
  assign n63357 = n63186 | n63356;
  assign n44661 = ~n63355 & n63357;
  assign n44662 = x151 & x228;
  assign n44663 = n44661 & n44662;
  assign n44664 = n44661 | n44662;
  assign n44665 = ~n44663 & n44664;
  assign n63358 = n44374 & n44665;
  assign n63359 = (n44665 & n63190) | (n44665 & n63358) | (n63190 & n63358);
  assign n63360 = n44374 | n44665;
  assign n63361 = n63190 | n63360;
  assign n44668 = ~n63359 & n63361;
  assign n44669 = x150 & x229;
  assign n44670 = n44668 & n44669;
  assign n44671 = n44668 | n44669;
  assign n44672 = ~n44670 & n44671;
  assign n63362 = n44381 & n44672;
  assign n63363 = (n44672 & n63194) | (n44672 & n63362) | (n63194 & n63362);
  assign n63364 = n44381 | n44672;
  assign n63365 = n63194 | n63364;
  assign n44675 = ~n63363 & n63365;
  assign n44676 = x149 & x230;
  assign n44677 = n44675 & n44676;
  assign n44678 = n44675 | n44676;
  assign n44679 = ~n44677 & n44678;
  assign n63366 = n44388 & n44679;
  assign n63367 = (n44679 & n63198) | (n44679 & n63366) | (n63198 & n63366);
  assign n63368 = n44388 | n44679;
  assign n63369 = n63198 | n63368;
  assign n44682 = ~n63367 & n63369;
  assign n44683 = x148 & x231;
  assign n44684 = n44682 & n44683;
  assign n44685 = n44682 | n44683;
  assign n44686 = ~n44684 & n44685;
  assign n63370 = n44395 & n44686;
  assign n63371 = (n44686 & n63202) | (n44686 & n63370) | (n63202 & n63370);
  assign n63372 = n44395 | n44686;
  assign n63373 = n63202 | n63372;
  assign n44689 = ~n63371 & n63373;
  assign n44690 = x147 & x232;
  assign n44691 = n44689 & n44690;
  assign n44692 = n44689 | n44690;
  assign n44693 = ~n44691 & n44692;
  assign n63374 = n44402 & n44693;
  assign n63375 = (n44693 & n63206) | (n44693 & n63374) | (n63206 & n63374);
  assign n63376 = n44402 | n44693;
  assign n63377 = n63206 | n63376;
  assign n44696 = ~n63375 & n63377;
  assign n44697 = x146 & x233;
  assign n44698 = n44696 & n44697;
  assign n44699 = n44696 | n44697;
  assign n44700 = ~n44698 & n44699;
  assign n63378 = n44409 & n44700;
  assign n63379 = (n44700 & n63210) | (n44700 & n63378) | (n63210 & n63378);
  assign n63380 = n44409 | n44700;
  assign n63381 = n63210 | n63380;
  assign n44703 = ~n63379 & n63381;
  assign n44704 = x145 & x234;
  assign n44705 = n44703 & n44704;
  assign n44706 = n44703 | n44704;
  assign n44707 = ~n44705 & n44706;
  assign n63382 = n44416 & n44707;
  assign n63383 = (n44707 & n63214) | (n44707 & n63382) | (n63214 & n63382);
  assign n63384 = n44416 | n44707;
  assign n63385 = n63214 | n63384;
  assign n44710 = ~n63383 & n63385;
  assign n44711 = x144 & x235;
  assign n44712 = n44710 & n44711;
  assign n44713 = n44710 | n44711;
  assign n44714 = ~n44712 & n44713;
  assign n63386 = n44423 & n44714;
  assign n63387 = (n44714 & n63218) | (n44714 & n63386) | (n63218 & n63386);
  assign n63388 = n44423 | n44714;
  assign n63389 = n63218 | n63388;
  assign n44717 = ~n63387 & n63389;
  assign n44718 = x143 & x236;
  assign n44719 = n44717 & n44718;
  assign n44720 = n44717 | n44718;
  assign n44721 = ~n44719 & n44720;
  assign n63390 = n44430 & n44721;
  assign n63391 = (n44721 & n63222) | (n44721 & n63390) | (n63222 & n63390);
  assign n63392 = n44430 | n44721;
  assign n63393 = n63222 | n63392;
  assign n44724 = ~n63391 & n63393;
  assign n44725 = x142 & x237;
  assign n44726 = n44724 & n44725;
  assign n44727 = n44724 | n44725;
  assign n44728 = ~n44726 & n44727;
  assign n63394 = n44437 & n44728;
  assign n63395 = (n44728 & n63226) | (n44728 & n63394) | (n63226 & n63394);
  assign n63396 = n44437 | n44728;
  assign n63397 = n63226 | n63396;
  assign n44731 = ~n63395 & n63397;
  assign n44732 = x141 & x238;
  assign n44733 = n44731 & n44732;
  assign n44734 = n44731 | n44732;
  assign n44735 = ~n44733 & n44734;
  assign n63398 = n44444 & n44735;
  assign n63399 = (n44735 & n63230) | (n44735 & n63398) | (n63230 & n63398);
  assign n63400 = n44444 | n44735;
  assign n63401 = n63230 | n63400;
  assign n44738 = ~n63399 & n63401;
  assign n44739 = x140 & x239;
  assign n44740 = n44738 & n44739;
  assign n44741 = n44738 | n44739;
  assign n44742 = ~n44740 & n44741;
  assign n63402 = n44451 & n44742;
  assign n63403 = (n44742 & n63234) | (n44742 & n63402) | (n63234 & n63402);
  assign n63404 = n44451 | n44742;
  assign n63405 = n63234 | n63404;
  assign n44745 = ~n63403 & n63405;
  assign n63412 = n44565 | n44567;
  assign n73632 = n44276 | n44565;
  assign n73633 = (n44565 & n44567) | (n44565 & n73632) | (n44567 & n73632);
  assign n73634 = (n63136 & n63412) | (n63136 & n73633) | (n63412 & n73633);
  assign n73635 = (n63135 & n63412) | (n63135 & n73633) | (n63412 & n73633);
  assign n73636 = (n73458 & n73634) | (n73458 & n73635) | (n73634 & n73635);
  assign n63417 = n44544 | n44546;
  assign n73637 = n44255 | n44544;
  assign n73638 = (n44544 & n44546) | (n44544 & n73637) | (n44546 & n73637);
  assign n73639 = (n63126 & n63417) | (n63126 & n73638) | (n63417 & n73638);
  assign n73640 = (n63125 & n63417) | (n63125 & n73638) | (n63417 & n73638);
  assign n73641 = (n73463 & n73639) | (n73463 & n73640) | (n73639 & n73640);
  assign n63251 = (n62950 & n73583) | (n62950 & n63250) | (n73583 & n63250);
  assign n63422 = n44523 | n44525;
  assign n73642 = n44234 | n44523;
  assign n73643 = (n44523 & n44525) | (n44523 & n73642) | (n44525 & n73642);
  assign n73644 = (n63116 & n63422) | (n63116 & n73643) | (n63422 & n73643);
  assign n73645 = (n63115 & n63422) | (n63115 & n73643) | (n63422 & n73643);
  assign n73646 = (n62913 & n73644) | (n62913 & n73645) | (n73644 & n73645);
  assign n63256 = (n62940 & n73585) | (n62940 & n63255) | (n73585 & n63255);
  assign n63427 = n44502 | n44504;
  assign n73647 = n44213 | n44502;
  assign n73648 = (n44502 & n44504) | (n44502 & n73647) | (n44504 & n73647);
  assign n73649 = (n63106 & n63427) | (n63106 & n73648) | (n63427 & n73648);
  assign n73650 = (n63105 & n63427) | (n63105 & n73648) | (n63427 & n73648);
  assign n73651 = (n62918 & n73649) | (n62918 & n73650) | (n73649 & n73650);
  assign n44782 = x175 & x205;
  assign n73652 = n44782 & n63262;
  assign n73653 = n44782 & n73589;
  assign n73654 = (n62930 & n73652) | (n62930 & n73653) | (n73652 & n73653);
  assign n73655 = (n44782 & n73592) | (n44782 & n73654) | (n73592 & n73654);
  assign n73656 = (n44782 & n63269) | (n44782 & n73654) | (n63269 & n73654);
  assign n73657 = (n73533 & n73655) | (n73533 & n73656) | (n73655 & n73656);
  assign n73658 = n44782 | n63262;
  assign n73659 = n44782 | n73589;
  assign n73660 = (n62930 & n73658) | (n62930 & n73659) | (n73658 & n73659);
  assign n73661 = n73592 | n73660;
  assign n73662 = n63269 | n73660;
  assign n73663 = (n73533 & n73661) | (n73533 & n73662) | (n73661 & n73662);
  assign n44785 = ~n73657 & n73663;
  assign n44786 = n73651 & n44785;
  assign n44787 = n73651 | n44785;
  assign n44788 = ~n44786 & n44787;
  assign n44789 = x174 & x206;
  assign n44790 = n44788 & n44789;
  assign n44791 = n44788 | n44789;
  assign n44792 = ~n44790 & n44791;
  assign n63424 = n44509 | n44511;
  assign n63433 = n44792 & n63424;
  assign n63434 = n44509 & n44792;
  assign n63435 = (n63256 & n63433) | (n63256 & n63434) | (n63433 & n63434);
  assign n63436 = n44792 | n63424;
  assign n63437 = n44509 | n44792;
  assign n63438 = (n63256 & n63436) | (n63256 & n63437) | (n63436 & n63437);
  assign n44795 = ~n63435 & n63438;
  assign n44796 = x173 & x207;
  assign n44797 = n44795 & n44796;
  assign n44798 = n44795 | n44796;
  assign n44799 = ~n44797 & n44798;
  assign n63439 = n44516 & n44799;
  assign n63440 = (n44799 & n63280) | (n44799 & n63439) | (n63280 & n63439);
  assign n63441 = n44516 | n44799;
  assign n63442 = n63280 | n63441;
  assign n44802 = ~n63440 & n63442;
  assign n44803 = x172 & x208;
  assign n44804 = n44802 & n44803;
  assign n44805 = n44802 | n44803;
  assign n44806 = ~n44804 & n44805;
  assign n44807 = n73646 & n44806;
  assign n44808 = n73646 | n44806;
  assign n44809 = ~n44807 & n44808;
  assign n44810 = x171 & x209;
  assign n44811 = n44809 & n44810;
  assign n44812 = n44809 | n44810;
  assign n44813 = ~n44811 & n44812;
  assign n63419 = n44530 | n44532;
  assign n63443 = n44813 & n63419;
  assign n63444 = n44530 & n44813;
  assign n63445 = (n63251 & n63443) | (n63251 & n63444) | (n63443 & n63444);
  assign n63446 = n44813 | n63419;
  assign n63447 = n44530 | n44813;
  assign n63448 = (n63251 & n63446) | (n63251 & n63447) | (n63446 & n63447);
  assign n44816 = ~n63445 & n63448;
  assign n44817 = x170 & x210;
  assign n44818 = n44816 & n44817;
  assign n44819 = n44816 | n44817;
  assign n44820 = ~n44818 & n44819;
  assign n63449 = n44537 & n44820;
  assign n63450 = (n44820 & n63290) | (n44820 & n63449) | (n63290 & n63449);
  assign n63451 = n44537 | n44820;
  assign n63452 = n63290 | n63451;
  assign n44823 = ~n63450 & n63452;
  assign n44824 = x169 & x211;
  assign n44825 = n44823 & n44824;
  assign n44826 = n44823 | n44824;
  assign n44827 = ~n44825 & n44826;
  assign n44828 = n73641 & n44827;
  assign n44829 = n73641 | n44827;
  assign n44830 = ~n44828 & n44829;
  assign n44831 = x168 & x212;
  assign n44832 = n44830 & n44831;
  assign n44833 = n44830 | n44831;
  assign n44834 = ~n44832 & n44833;
  assign n63414 = n44551 | n44553;
  assign n63453 = n44834 & n63414;
  assign n63454 = n44551 & n44834;
  assign n63455 = (n73581 & n63453) | (n73581 & n63454) | (n63453 & n63454);
  assign n63456 = n44834 | n63414;
  assign n63457 = n44551 | n44834;
  assign n63458 = (n73581 & n63456) | (n73581 & n63457) | (n63456 & n63457);
  assign n44837 = ~n63455 & n63458;
  assign n44838 = x167 & x213;
  assign n44839 = n44837 & n44838;
  assign n44840 = n44837 | n44838;
  assign n44841 = ~n44839 & n44840;
  assign n63459 = n44558 & n44841;
  assign n73664 = (n44841 & n63299) | (n44841 & n63459) | (n63299 & n63459);
  assign n73665 = (n44841 & n63298) | (n44841 & n63459) | (n63298 & n63459);
  assign n73666 = (n73518 & n73664) | (n73518 & n73665) | (n73664 & n73665);
  assign n63461 = n44558 | n44841;
  assign n73667 = n63299 | n63461;
  assign n73668 = n63298 | n63461;
  assign n73669 = (n73518 & n73667) | (n73518 & n73668) | (n73667 & n73668);
  assign n44844 = ~n73666 & n73669;
  assign n44845 = x166 & x214;
  assign n44846 = n44844 & n44845;
  assign n44847 = n44844 | n44845;
  assign n44848 = ~n44846 & n44847;
  assign n44849 = n73636 & n44848;
  assign n44850 = n73636 | n44848;
  assign n44851 = ~n44849 & n44850;
  assign n44852 = x165 & x215;
  assign n44853 = n44851 & n44852;
  assign n44854 = n44851 | n44852;
  assign n44855 = ~n44853 & n44854;
  assign n63409 = n44572 | n44574;
  assign n63463 = n44855 & n63409;
  assign n63464 = n44572 & n44855;
  assign n63465 = (n73576 & n63463) | (n73576 & n63464) | (n63463 & n63464);
  assign n63466 = n44855 | n63409;
  assign n63467 = n44572 | n44855;
  assign n63468 = (n73576 & n63466) | (n73576 & n63467) | (n63466 & n63467);
  assign n44858 = ~n63465 & n63468;
  assign n44859 = x164 & x216;
  assign n44860 = n44858 & n44859;
  assign n44861 = n44858 | n44859;
  assign n44862 = ~n44860 & n44861;
  assign n63469 = n44579 & n44862;
  assign n73670 = (n44862 & n63309) | (n44862 & n63469) | (n63309 & n63469);
  assign n73671 = (n44862 & n63308) | (n44862 & n63469) | (n63308 & n63469);
  assign n73672 = (n63072 & n73670) | (n63072 & n73671) | (n73670 & n73671);
  assign n63471 = n44579 | n44862;
  assign n73673 = n63309 | n63471;
  assign n73674 = n63308 | n63471;
  assign n73675 = (n63072 & n73673) | (n63072 & n73674) | (n73673 & n73674);
  assign n44865 = ~n73672 & n73675;
  assign n44866 = x163 & x217;
  assign n44867 = n44865 & n44866;
  assign n44868 = n44865 | n44866;
  assign n44869 = ~n44867 & n44868;
  assign n63407 = n44586 | n44588;
  assign n73676 = n44869 & n63407;
  assign n73630 = n44297 | n44586;
  assign n73631 = (n44586 & n44588) | (n44586 & n73630) | (n44588 & n73630);
  assign n73677 = n44869 & n73631;
  assign n73678 = (n73568 & n73676) | (n73568 & n73677) | (n73676 & n73677);
  assign n73679 = n44869 | n63407;
  assign n73680 = n44869 | n73631;
  assign n73681 = (n73568 & n73679) | (n73568 & n73680) | (n73679 & n73680);
  assign n44872 = ~n73678 & n73681;
  assign n44873 = x162 & x218;
  assign n44874 = n44872 & n44873;
  assign n44875 = n44872 | n44873;
  assign n44876 = ~n44874 & n44875;
  assign n63473 = n44593 & n44876;
  assign n73682 = (n44876 & n63318) | (n44876 & n63473) | (n63318 & n63473);
  assign n73683 = (n44595 & n44876) | (n44595 & n63473) | (n44876 & n63473);
  assign n73684 = (n63150 & n73682) | (n63150 & n73683) | (n73682 & n73683);
  assign n63475 = n44593 | n44876;
  assign n73685 = n63318 | n63475;
  assign n73686 = n44595 | n63475;
  assign n73687 = (n63150 & n73685) | (n63150 & n73686) | (n73685 & n73686);
  assign n44879 = ~n73684 & n73687;
  assign n44880 = x161 & x219;
  assign n44881 = n44879 & n44880;
  assign n44882 = n44879 | n44880;
  assign n44883 = ~n44881 & n44882;
  assign n63477 = n44600 & n44883;
  assign n63478 = (n44883 & n63323) | (n44883 & n63477) | (n63323 & n63477);
  assign n63479 = n44600 | n44883;
  assign n63480 = n63323 | n63479;
  assign n44886 = ~n63478 & n63480;
  assign n44887 = x160 & x220;
  assign n44888 = n44886 & n44887;
  assign n44889 = n44886 | n44887;
  assign n44890 = ~n44888 & n44889;
  assign n63481 = n44607 & n44890;
  assign n63482 = (n44890 & n63327) | (n44890 & n63481) | (n63327 & n63481);
  assign n63483 = n44607 | n44890;
  assign n63484 = n63327 | n63483;
  assign n44893 = ~n63482 & n63484;
  assign n44894 = x159 & x221;
  assign n44895 = n44893 & n44894;
  assign n44896 = n44893 | n44894;
  assign n44897 = ~n44895 & n44896;
  assign n63485 = n44614 & n44897;
  assign n63486 = (n44897 & n63331) | (n44897 & n63485) | (n63331 & n63485);
  assign n63487 = n44614 | n44897;
  assign n63488 = n63331 | n63487;
  assign n44900 = ~n63486 & n63488;
  assign n44901 = x158 & x222;
  assign n44902 = n44900 & n44901;
  assign n44903 = n44900 | n44901;
  assign n44904 = ~n44902 & n44903;
  assign n63489 = n44621 & n44904;
  assign n63490 = (n44904 & n63335) | (n44904 & n63489) | (n63335 & n63489);
  assign n63491 = n44621 | n44904;
  assign n63492 = n63335 | n63491;
  assign n44907 = ~n63490 & n63492;
  assign n44908 = x157 & x223;
  assign n44909 = n44907 & n44908;
  assign n44910 = n44907 | n44908;
  assign n44911 = ~n44909 & n44910;
  assign n63493 = n44628 & n44911;
  assign n63494 = (n44911 & n63339) | (n44911 & n63493) | (n63339 & n63493);
  assign n63495 = n44628 | n44911;
  assign n63496 = n63339 | n63495;
  assign n44914 = ~n63494 & n63496;
  assign n44915 = x156 & x224;
  assign n44916 = n44914 & n44915;
  assign n44917 = n44914 | n44915;
  assign n44918 = ~n44916 & n44917;
  assign n63497 = n44635 & n44918;
  assign n63498 = (n44918 & n63343) | (n44918 & n63497) | (n63343 & n63497);
  assign n63499 = n44635 | n44918;
  assign n63500 = n63343 | n63499;
  assign n44921 = ~n63498 & n63500;
  assign n44922 = x155 & x225;
  assign n44923 = n44921 & n44922;
  assign n44924 = n44921 | n44922;
  assign n44925 = ~n44923 & n44924;
  assign n63501 = n44642 & n44925;
  assign n63502 = (n44925 & n63347) | (n44925 & n63501) | (n63347 & n63501);
  assign n63503 = n44642 | n44925;
  assign n63504 = n63347 | n63503;
  assign n44928 = ~n63502 & n63504;
  assign n44929 = x154 & x226;
  assign n44930 = n44928 & n44929;
  assign n44931 = n44928 | n44929;
  assign n44932 = ~n44930 & n44931;
  assign n63505 = n44649 & n44932;
  assign n63506 = (n44932 & n63351) | (n44932 & n63505) | (n63351 & n63505);
  assign n63507 = n44649 | n44932;
  assign n63508 = n63351 | n63507;
  assign n44935 = ~n63506 & n63508;
  assign n44936 = x153 & x227;
  assign n44937 = n44935 & n44936;
  assign n44938 = n44935 | n44936;
  assign n44939 = ~n44937 & n44938;
  assign n63509 = n44656 & n44939;
  assign n63510 = (n44939 & n63355) | (n44939 & n63509) | (n63355 & n63509);
  assign n63511 = n44656 | n44939;
  assign n63512 = n63355 | n63511;
  assign n44942 = ~n63510 & n63512;
  assign n44943 = x152 & x228;
  assign n44944 = n44942 & n44943;
  assign n44945 = n44942 | n44943;
  assign n44946 = ~n44944 & n44945;
  assign n63513 = n44663 & n44946;
  assign n63514 = (n44946 & n63359) | (n44946 & n63513) | (n63359 & n63513);
  assign n63515 = n44663 | n44946;
  assign n63516 = n63359 | n63515;
  assign n44949 = ~n63514 & n63516;
  assign n44950 = x151 & x229;
  assign n44951 = n44949 & n44950;
  assign n44952 = n44949 | n44950;
  assign n44953 = ~n44951 & n44952;
  assign n63517 = n44670 & n44953;
  assign n63518 = (n44953 & n63363) | (n44953 & n63517) | (n63363 & n63517);
  assign n63519 = n44670 | n44953;
  assign n63520 = n63363 | n63519;
  assign n44956 = ~n63518 & n63520;
  assign n44957 = x150 & x230;
  assign n44958 = n44956 & n44957;
  assign n44959 = n44956 | n44957;
  assign n44960 = ~n44958 & n44959;
  assign n63521 = n44677 & n44960;
  assign n63522 = (n44960 & n63367) | (n44960 & n63521) | (n63367 & n63521);
  assign n63523 = n44677 | n44960;
  assign n63524 = n63367 | n63523;
  assign n44963 = ~n63522 & n63524;
  assign n44964 = x149 & x231;
  assign n44965 = n44963 & n44964;
  assign n44966 = n44963 | n44964;
  assign n44967 = ~n44965 & n44966;
  assign n63525 = n44684 & n44967;
  assign n63526 = (n44967 & n63371) | (n44967 & n63525) | (n63371 & n63525);
  assign n63527 = n44684 | n44967;
  assign n63528 = n63371 | n63527;
  assign n44970 = ~n63526 & n63528;
  assign n44971 = x148 & x232;
  assign n44972 = n44970 & n44971;
  assign n44973 = n44970 | n44971;
  assign n44974 = ~n44972 & n44973;
  assign n63529 = n44691 & n44974;
  assign n63530 = (n44974 & n63375) | (n44974 & n63529) | (n63375 & n63529);
  assign n63531 = n44691 | n44974;
  assign n63532 = n63375 | n63531;
  assign n44977 = ~n63530 & n63532;
  assign n44978 = x147 & x233;
  assign n44979 = n44977 & n44978;
  assign n44980 = n44977 | n44978;
  assign n44981 = ~n44979 & n44980;
  assign n63533 = n44698 & n44981;
  assign n63534 = (n44981 & n63379) | (n44981 & n63533) | (n63379 & n63533);
  assign n63535 = n44698 | n44981;
  assign n63536 = n63379 | n63535;
  assign n44984 = ~n63534 & n63536;
  assign n44985 = x146 & x234;
  assign n44986 = n44984 & n44985;
  assign n44987 = n44984 | n44985;
  assign n44988 = ~n44986 & n44987;
  assign n63537 = n44705 & n44988;
  assign n63538 = (n44988 & n63383) | (n44988 & n63537) | (n63383 & n63537);
  assign n63539 = n44705 | n44988;
  assign n63540 = n63383 | n63539;
  assign n44991 = ~n63538 & n63540;
  assign n44992 = x145 & x235;
  assign n44993 = n44991 & n44992;
  assign n44994 = n44991 | n44992;
  assign n44995 = ~n44993 & n44994;
  assign n63541 = n44712 & n44995;
  assign n63542 = (n44995 & n63387) | (n44995 & n63541) | (n63387 & n63541);
  assign n63543 = n44712 | n44995;
  assign n63544 = n63387 | n63543;
  assign n44998 = ~n63542 & n63544;
  assign n44999 = x144 & x236;
  assign n45000 = n44998 & n44999;
  assign n45001 = n44998 | n44999;
  assign n45002 = ~n45000 & n45001;
  assign n63545 = n44719 & n45002;
  assign n63546 = (n45002 & n63391) | (n45002 & n63545) | (n63391 & n63545);
  assign n63547 = n44719 | n45002;
  assign n63548 = n63391 | n63547;
  assign n45005 = ~n63546 & n63548;
  assign n45006 = x143 & x237;
  assign n45007 = n45005 & n45006;
  assign n45008 = n45005 | n45006;
  assign n45009 = ~n45007 & n45008;
  assign n63549 = n44726 & n45009;
  assign n63550 = (n45009 & n63395) | (n45009 & n63549) | (n63395 & n63549);
  assign n63551 = n44726 | n45009;
  assign n63552 = n63395 | n63551;
  assign n45012 = ~n63550 & n63552;
  assign n45013 = x142 & x238;
  assign n45014 = n45012 & n45013;
  assign n45015 = n45012 | n45013;
  assign n45016 = ~n45014 & n45015;
  assign n63553 = n44733 & n45016;
  assign n63554 = (n45016 & n63399) | (n45016 & n63553) | (n63399 & n63553);
  assign n63555 = n44733 | n45016;
  assign n63556 = n63399 | n63555;
  assign n45019 = ~n63554 & n63556;
  assign n45020 = x141 & x239;
  assign n45021 = n45019 & n45020;
  assign n45022 = n45019 | n45020;
  assign n45023 = ~n45021 & n45022;
  assign n63557 = n44740 & n45023;
  assign n63558 = (n45023 & n63403) | (n45023 & n63557) | (n63403 & n63557);
  assign n63559 = n44740 | n45023;
  assign n63560 = n63403 | n63559;
  assign n45026 = ~n63558 & n63560;
  assign n63408 = (n73568 & n73631) | (n73568 & n63407) | (n73631 & n63407);
  assign n63564 = n44860 | n44862;
  assign n73688 = n44579 | n44860;
  assign n73689 = (n44860 & n44862) | (n44860 & n73688) | (n44862 & n73688);
  assign n73690 = (n63309 & n63564) | (n63309 & n73689) | (n63564 & n73689);
  assign n73691 = (n63308 & n63564) | (n63308 & n73689) | (n63564 & n73689);
  assign n73692 = (n63072 & n73690) | (n63072 & n73691) | (n73690 & n73691);
  assign n63569 = n44839 | n44841;
  assign n73693 = n44558 | n44839;
  assign n73694 = (n44839 & n44841) | (n44839 & n73693) | (n44841 & n73693);
  assign n73695 = (n63299 & n63569) | (n63299 & n73694) | (n63569 & n73694);
  assign n73696 = (n63298 & n63569) | (n63298 & n73694) | (n63569 & n73694);
  assign n73697 = (n73518 & n73695) | (n73518 & n73696) | (n73695 & n73696);
  assign n45062 = x175 & x206;
  assign n73702 = n45062 & n73657;
  assign n73703 = (n44785 & n45062) | (n44785 & n73702) | (n45062 & n73702);
  assign n63584 = n45062 & n73657;
  assign n63585 = (n73651 & n73703) | (n73651 & n63584) | (n73703 & n63584);
  assign n73704 = n45062 | n73657;
  assign n73705 = n44785 | n73704;
  assign n63587 = n45062 | n73657;
  assign n63588 = (n73651 & n73705) | (n73651 & n63587) | (n73705 & n63587);
  assign n45065 = ~n63585 & n63588;
  assign n63589 = n44790 & n45065;
  assign n73706 = (n45065 & n63434) | (n45065 & n63589) | (n63434 & n63589);
  assign n73707 = (n45065 & n63433) | (n45065 & n63589) | (n63433 & n63589);
  assign n73708 = (n63256 & n73706) | (n63256 & n73707) | (n73706 & n73707);
  assign n63591 = n44790 | n45065;
  assign n73709 = n63434 | n63591;
  assign n73710 = n63433 | n63591;
  assign n73711 = (n63256 & n73709) | (n63256 & n73710) | (n73709 & n73710);
  assign n45068 = ~n73708 & n73711;
  assign n45069 = x174 & x207;
  assign n45070 = n45068 & n45069;
  assign n45071 = n45068 | n45069;
  assign n45072 = ~n45070 & n45071;
  assign n63579 = n44797 | n44799;
  assign n73712 = n45072 & n63579;
  assign n73700 = n44516 | n44797;
  assign n73701 = (n44797 & n44799) | (n44797 & n73700) | (n44799 & n73700);
  assign n73713 = n45072 & n73701;
  assign n73714 = (n63280 & n73712) | (n63280 & n73713) | (n73712 & n73713);
  assign n73715 = n45072 | n63579;
  assign n73716 = n45072 | n73701;
  assign n73717 = (n63280 & n73715) | (n63280 & n73716) | (n73715 & n73716);
  assign n45075 = ~n73714 & n73717;
  assign n45076 = x173 & x208;
  assign n45077 = n45075 & n45076;
  assign n45078 = n45075 | n45076;
  assign n45079 = ~n45077 & n45078;
  assign n63576 = n44804 | n44806;
  assign n63593 = n45079 & n63576;
  assign n63594 = n44804 & n45079;
  assign n63595 = (n73646 & n63593) | (n73646 & n63594) | (n63593 & n63594);
  assign n63596 = n45079 | n63576;
  assign n63597 = n44804 | n45079;
  assign n63598 = (n73646 & n63596) | (n73646 & n63597) | (n63596 & n63597);
  assign n45082 = ~n63595 & n63598;
  assign n45083 = x172 & x209;
  assign n45084 = n45082 & n45083;
  assign n45085 = n45082 | n45083;
  assign n45086 = ~n45084 & n45085;
  assign n63599 = n44811 & n45086;
  assign n73718 = (n45086 & n63444) | (n45086 & n63599) | (n63444 & n63599);
  assign n73719 = (n45086 & n63443) | (n45086 & n63599) | (n63443 & n63599);
  assign n73720 = (n63251 & n73718) | (n63251 & n73719) | (n73718 & n73719);
  assign n63601 = n44811 | n45086;
  assign n73721 = n63444 | n63601;
  assign n73722 = n63443 | n63601;
  assign n73723 = (n63251 & n73721) | (n63251 & n73722) | (n73721 & n73722);
  assign n45089 = ~n73720 & n73723;
  assign n45090 = x171 & x210;
  assign n45091 = n45089 & n45090;
  assign n45092 = n45089 | n45090;
  assign n45093 = ~n45091 & n45092;
  assign n63574 = n44818 | n44820;
  assign n73724 = n45093 & n63574;
  assign n73698 = n44537 | n44818;
  assign n73699 = (n44818 & n44820) | (n44818 & n73698) | (n44820 & n73698);
  assign n73725 = n45093 & n73699;
  assign n73726 = (n63290 & n73724) | (n63290 & n73725) | (n73724 & n73725);
  assign n73727 = n45093 | n63574;
  assign n73728 = n45093 | n73699;
  assign n73729 = (n63290 & n73727) | (n63290 & n73728) | (n73727 & n73728);
  assign n45096 = ~n73726 & n73729;
  assign n45097 = x170 & x211;
  assign n45098 = n45096 & n45097;
  assign n45099 = n45096 | n45097;
  assign n45100 = ~n45098 & n45099;
  assign n63571 = n44825 | n44827;
  assign n63603 = n45100 & n63571;
  assign n63604 = n44825 & n45100;
  assign n63605 = (n73641 & n63603) | (n73641 & n63604) | (n63603 & n63604);
  assign n63606 = n45100 | n63571;
  assign n63607 = n44825 | n45100;
  assign n63608 = (n73641 & n63606) | (n73641 & n63607) | (n63606 & n63607);
  assign n45103 = ~n63605 & n63608;
  assign n45104 = x169 & x212;
  assign n45105 = n45103 & n45104;
  assign n45106 = n45103 | n45104;
  assign n45107 = ~n45105 & n45106;
  assign n63609 = n44832 & n45107;
  assign n73730 = (n45107 & n63454) | (n45107 & n63609) | (n63454 & n63609);
  assign n73731 = (n45107 & n63453) | (n45107 & n63609) | (n63453 & n63609);
  assign n73732 = (n73581 & n73730) | (n73581 & n73731) | (n73730 & n73731);
  assign n63611 = n44832 | n45107;
  assign n73733 = n63454 | n63611;
  assign n73734 = n63453 | n63611;
  assign n73735 = (n73581 & n73733) | (n73581 & n73734) | (n73733 & n73734);
  assign n45110 = ~n73732 & n73735;
  assign n45111 = x168 & x213;
  assign n45112 = n45110 & n45111;
  assign n45113 = n45110 | n45111;
  assign n45114 = ~n45112 & n45113;
  assign n45115 = n73697 & n45114;
  assign n45116 = n73697 | n45114;
  assign n45117 = ~n45115 & n45116;
  assign n45118 = x167 & x214;
  assign n45119 = n45117 & n45118;
  assign n45120 = n45117 | n45118;
  assign n45121 = ~n45119 & n45120;
  assign n63566 = n44846 | n44848;
  assign n63613 = n45121 & n63566;
  assign n63614 = n44846 & n45121;
  assign n63615 = (n73636 & n63613) | (n73636 & n63614) | (n63613 & n63614);
  assign n63616 = n45121 | n63566;
  assign n63617 = n44846 | n45121;
  assign n63618 = (n73636 & n63616) | (n73636 & n63617) | (n63616 & n63617);
  assign n45124 = ~n63615 & n63618;
  assign n45125 = x166 & x215;
  assign n45126 = n45124 & n45125;
  assign n45127 = n45124 | n45125;
  assign n45128 = ~n45126 & n45127;
  assign n63619 = n44853 & n45128;
  assign n73736 = (n45128 & n63464) | (n45128 & n63619) | (n63464 & n63619);
  assign n73737 = (n45128 & n63463) | (n45128 & n63619) | (n63463 & n63619);
  assign n73738 = (n73576 & n73736) | (n73576 & n73737) | (n73736 & n73737);
  assign n63621 = n44853 | n45128;
  assign n73739 = n63464 | n63621;
  assign n73740 = n63463 | n63621;
  assign n73741 = (n73576 & n73739) | (n73576 & n73740) | (n73739 & n73740);
  assign n45131 = ~n73738 & n73741;
  assign n45132 = x165 & x216;
  assign n45133 = n45131 & n45132;
  assign n45134 = n45131 | n45132;
  assign n45135 = ~n45133 & n45134;
  assign n45136 = n73692 & n45135;
  assign n45137 = n73692 | n45135;
  assign n45138 = ~n45136 & n45137;
  assign n45139 = x164 & x217;
  assign n45140 = n45138 & n45139;
  assign n45141 = n45138 | n45139;
  assign n45142 = ~n45140 & n45141;
  assign n63561 = n44867 | n44869;
  assign n63623 = n45142 & n63561;
  assign n63624 = n44867 & n45142;
  assign n63625 = (n63408 & n63623) | (n63408 & n63624) | (n63623 & n63624);
  assign n63626 = n45142 | n63561;
  assign n63627 = n44867 | n45142;
  assign n63628 = (n63408 & n63626) | (n63408 & n63627) | (n63626 & n63627);
  assign n45145 = ~n63625 & n63628;
  assign n45146 = x163 & x218;
  assign n45147 = n45145 & n45146;
  assign n45148 = n45145 | n45146;
  assign n45149 = ~n45147 & n45148;
  assign n63629 = n44874 & n45149;
  assign n63630 = (n45149 & n73684) | (n45149 & n63629) | (n73684 & n63629);
  assign n63631 = n44874 | n45149;
  assign n63632 = n73684 | n63631;
  assign n45152 = ~n63630 & n63632;
  assign n45153 = x162 & x219;
  assign n45154 = n45152 & n45153;
  assign n45155 = n45152 | n45153;
  assign n45156 = ~n45154 & n45155;
  assign n63633 = n44881 & n45156;
  assign n63634 = (n45156 & n63478) | (n45156 & n63633) | (n63478 & n63633);
  assign n63635 = n44881 | n45156;
  assign n63636 = n63478 | n63635;
  assign n45159 = ~n63634 & n63636;
  assign n45160 = x161 & x220;
  assign n45161 = n45159 & n45160;
  assign n45162 = n45159 | n45160;
  assign n45163 = ~n45161 & n45162;
  assign n63637 = n44888 & n45163;
  assign n63638 = (n45163 & n63482) | (n45163 & n63637) | (n63482 & n63637);
  assign n63639 = n44888 | n45163;
  assign n63640 = n63482 | n63639;
  assign n45166 = ~n63638 & n63640;
  assign n45167 = x160 & x221;
  assign n45168 = n45166 & n45167;
  assign n45169 = n45166 | n45167;
  assign n45170 = ~n45168 & n45169;
  assign n63641 = n44895 & n45170;
  assign n63642 = (n45170 & n63486) | (n45170 & n63641) | (n63486 & n63641);
  assign n63643 = n44895 | n45170;
  assign n63644 = n63486 | n63643;
  assign n45173 = ~n63642 & n63644;
  assign n45174 = x159 & x222;
  assign n45175 = n45173 & n45174;
  assign n45176 = n45173 | n45174;
  assign n45177 = ~n45175 & n45176;
  assign n63645 = n44902 & n45177;
  assign n63646 = (n45177 & n63490) | (n45177 & n63645) | (n63490 & n63645);
  assign n63647 = n44902 | n45177;
  assign n63648 = n63490 | n63647;
  assign n45180 = ~n63646 & n63648;
  assign n45181 = x158 & x223;
  assign n45182 = n45180 & n45181;
  assign n45183 = n45180 | n45181;
  assign n45184 = ~n45182 & n45183;
  assign n63649 = n44909 & n45184;
  assign n63650 = (n45184 & n63494) | (n45184 & n63649) | (n63494 & n63649);
  assign n63651 = n44909 | n45184;
  assign n63652 = n63494 | n63651;
  assign n45187 = ~n63650 & n63652;
  assign n45188 = x157 & x224;
  assign n45189 = n45187 & n45188;
  assign n45190 = n45187 | n45188;
  assign n45191 = ~n45189 & n45190;
  assign n63653 = n44916 & n45191;
  assign n63654 = (n45191 & n63498) | (n45191 & n63653) | (n63498 & n63653);
  assign n63655 = n44916 | n45191;
  assign n63656 = n63498 | n63655;
  assign n45194 = ~n63654 & n63656;
  assign n45195 = x156 & x225;
  assign n45196 = n45194 & n45195;
  assign n45197 = n45194 | n45195;
  assign n45198 = ~n45196 & n45197;
  assign n63657 = n44923 & n45198;
  assign n63658 = (n45198 & n63502) | (n45198 & n63657) | (n63502 & n63657);
  assign n63659 = n44923 | n45198;
  assign n63660 = n63502 | n63659;
  assign n45201 = ~n63658 & n63660;
  assign n45202 = x155 & x226;
  assign n45203 = n45201 & n45202;
  assign n45204 = n45201 | n45202;
  assign n45205 = ~n45203 & n45204;
  assign n63661 = n44930 & n45205;
  assign n63662 = (n45205 & n63506) | (n45205 & n63661) | (n63506 & n63661);
  assign n63663 = n44930 | n45205;
  assign n63664 = n63506 | n63663;
  assign n45208 = ~n63662 & n63664;
  assign n45209 = x154 & x227;
  assign n45210 = n45208 & n45209;
  assign n45211 = n45208 | n45209;
  assign n45212 = ~n45210 & n45211;
  assign n63665 = n44937 & n45212;
  assign n63666 = (n45212 & n63510) | (n45212 & n63665) | (n63510 & n63665);
  assign n63667 = n44937 | n45212;
  assign n63668 = n63510 | n63667;
  assign n45215 = ~n63666 & n63668;
  assign n45216 = x153 & x228;
  assign n45217 = n45215 & n45216;
  assign n45218 = n45215 | n45216;
  assign n45219 = ~n45217 & n45218;
  assign n63669 = n44944 & n45219;
  assign n63670 = (n45219 & n63514) | (n45219 & n63669) | (n63514 & n63669);
  assign n63671 = n44944 | n45219;
  assign n63672 = n63514 | n63671;
  assign n45222 = ~n63670 & n63672;
  assign n45223 = x152 & x229;
  assign n45224 = n45222 & n45223;
  assign n45225 = n45222 | n45223;
  assign n45226 = ~n45224 & n45225;
  assign n63673 = n44951 & n45226;
  assign n63674 = (n45226 & n63518) | (n45226 & n63673) | (n63518 & n63673);
  assign n63675 = n44951 | n45226;
  assign n63676 = n63518 | n63675;
  assign n45229 = ~n63674 & n63676;
  assign n45230 = x151 & x230;
  assign n45231 = n45229 & n45230;
  assign n45232 = n45229 | n45230;
  assign n45233 = ~n45231 & n45232;
  assign n63677 = n44958 & n45233;
  assign n63678 = (n45233 & n63522) | (n45233 & n63677) | (n63522 & n63677);
  assign n63679 = n44958 | n45233;
  assign n63680 = n63522 | n63679;
  assign n45236 = ~n63678 & n63680;
  assign n45237 = x150 & x231;
  assign n45238 = n45236 & n45237;
  assign n45239 = n45236 | n45237;
  assign n45240 = ~n45238 & n45239;
  assign n63681 = n44965 & n45240;
  assign n63682 = (n45240 & n63526) | (n45240 & n63681) | (n63526 & n63681);
  assign n63683 = n44965 | n45240;
  assign n63684 = n63526 | n63683;
  assign n45243 = ~n63682 & n63684;
  assign n45244 = x149 & x232;
  assign n45245 = n45243 & n45244;
  assign n45246 = n45243 | n45244;
  assign n45247 = ~n45245 & n45246;
  assign n63685 = n44972 & n45247;
  assign n63686 = (n45247 & n63530) | (n45247 & n63685) | (n63530 & n63685);
  assign n63687 = n44972 | n45247;
  assign n63688 = n63530 | n63687;
  assign n45250 = ~n63686 & n63688;
  assign n45251 = x148 & x233;
  assign n45252 = n45250 & n45251;
  assign n45253 = n45250 | n45251;
  assign n45254 = ~n45252 & n45253;
  assign n63689 = n44979 & n45254;
  assign n63690 = (n45254 & n63534) | (n45254 & n63689) | (n63534 & n63689);
  assign n63691 = n44979 | n45254;
  assign n63692 = n63534 | n63691;
  assign n45257 = ~n63690 & n63692;
  assign n45258 = x147 & x234;
  assign n45259 = n45257 & n45258;
  assign n45260 = n45257 | n45258;
  assign n45261 = ~n45259 & n45260;
  assign n63693 = n44986 & n45261;
  assign n63694 = (n45261 & n63538) | (n45261 & n63693) | (n63538 & n63693);
  assign n63695 = n44986 | n45261;
  assign n63696 = n63538 | n63695;
  assign n45264 = ~n63694 & n63696;
  assign n45265 = x146 & x235;
  assign n45266 = n45264 & n45265;
  assign n45267 = n45264 | n45265;
  assign n45268 = ~n45266 & n45267;
  assign n63697 = n44993 & n45268;
  assign n63698 = (n45268 & n63542) | (n45268 & n63697) | (n63542 & n63697);
  assign n63699 = n44993 | n45268;
  assign n63700 = n63542 | n63699;
  assign n45271 = ~n63698 & n63700;
  assign n45272 = x145 & x236;
  assign n45273 = n45271 & n45272;
  assign n45274 = n45271 | n45272;
  assign n45275 = ~n45273 & n45274;
  assign n63701 = n45000 & n45275;
  assign n63702 = (n45275 & n63546) | (n45275 & n63701) | (n63546 & n63701);
  assign n63703 = n45000 | n45275;
  assign n63704 = n63546 | n63703;
  assign n45278 = ~n63702 & n63704;
  assign n45279 = x144 & x237;
  assign n45280 = n45278 & n45279;
  assign n45281 = n45278 | n45279;
  assign n45282 = ~n45280 & n45281;
  assign n63705 = n45007 & n45282;
  assign n63706 = (n45282 & n63550) | (n45282 & n63705) | (n63550 & n63705);
  assign n63707 = n45007 | n45282;
  assign n63708 = n63550 | n63707;
  assign n45285 = ~n63706 & n63708;
  assign n45286 = x143 & x238;
  assign n45287 = n45285 & n45286;
  assign n45288 = n45285 | n45286;
  assign n45289 = ~n45287 & n45288;
  assign n63709 = n45014 & n45289;
  assign n63710 = (n45289 & n63554) | (n45289 & n63709) | (n63554 & n63709);
  assign n63711 = n45014 | n45289;
  assign n63712 = n63554 | n63711;
  assign n45292 = ~n63710 & n63712;
  assign n45293 = x142 & x239;
  assign n45294 = n45292 & n45293;
  assign n45295 = n45292 | n45293;
  assign n45296 = ~n45294 & n45295;
  assign n63713 = n45021 & n45296;
  assign n63714 = (n45296 & n63558) | (n45296 & n63713) | (n63558 & n63713);
  assign n63715 = n45021 | n45296;
  assign n63716 = n63558 | n63715;
  assign n45299 = ~n63714 & n63716;
  assign n63723 = n45126 | n45128;
  assign n73744 = n44853 | n45126;
  assign n73745 = (n45126 & n45128) | (n45126 & n73744) | (n45128 & n73744);
  assign n73746 = (n63464 & n63723) | (n63464 & n73745) | (n63723 & n73745);
  assign n73747 = (n63463 & n63723) | (n63463 & n73745) | (n63723 & n73745);
  assign n73748 = (n73576 & n73746) | (n73576 & n73747) | (n73746 & n73747);
  assign n63728 = n45105 | n45107;
  assign n73749 = n44832 | n45105;
  assign n73750 = (n45105 & n45107) | (n45105 & n73749) | (n45107 & n73749);
  assign n73751 = (n63454 & n63728) | (n63454 & n73750) | (n63728 & n73750);
  assign n73752 = (n63453 & n63728) | (n63453 & n73750) | (n63728 & n73750);
  assign n73753 = (n73581 & n73751) | (n73581 & n73752) | (n73751 & n73752);
  assign n63575 = (n63290 & n73699) | (n63290 & n63574) | (n73699 & n63574);
  assign n63733 = n45084 | n45086;
  assign n73754 = n44811 | n45084;
  assign n73755 = (n45084 & n45086) | (n45084 & n73754) | (n45086 & n73754);
  assign n73756 = (n63444 & n63733) | (n63444 & n73755) | (n63733 & n73755);
  assign n73757 = (n63443 & n63733) | (n63443 & n73755) | (n63733 & n73755);
  assign n73758 = (n63251 & n73756) | (n63251 & n73757) | (n73756 & n73757);
  assign n45334 = x175 & x207;
  assign n63738 = n45065 | n63585;
  assign n73759 = (n44790 & n63585) | (n44790 & n63738) | (n63585 & n63738);
  assign n63740 = n45334 & n73759;
  assign n73760 = n45334 & n63585;
  assign n73761 = (n45065 & n45334) | (n45065 & n73760) | (n45334 & n73760);
  assign n73762 = (n63434 & n63740) | (n63434 & n73761) | (n63740 & n73761);
  assign n73763 = (n63433 & n63740) | (n63433 & n73761) | (n63740 & n73761);
  assign n73764 = (n63256 & n73762) | (n63256 & n73763) | (n73762 & n73763);
  assign n63743 = n45334 | n73759;
  assign n73765 = n45334 | n63585;
  assign n73766 = n45065 | n73765;
  assign n73767 = (n63434 & n63743) | (n63434 & n73766) | (n63743 & n73766);
  assign n73768 = (n63433 & n63743) | (n63433 & n73766) | (n63743 & n73766);
  assign n73769 = (n63256 & n73767) | (n63256 & n73768) | (n73767 & n73768);
  assign n45337 = ~n73764 & n73769;
  assign n63747 = n45070 & n45337;
  assign n73770 = (n45072 & n45337) | (n45072 & n63747) | (n45337 & n63747);
  assign n73771 = (n63579 & n63747) | (n63579 & n73770) | (n63747 & n73770);
  assign n73772 = (n63747 & n73701) | (n63747 & n73770) | (n73701 & n73770);
  assign n73773 = (n63280 & n73771) | (n63280 & n73772) | (n73771 & n73772);
  assign n63750 = n45070 | n45337;
  assign n73774 = n45072 | n63750;
  assign n73775 = (n63579 & n63750) | (n63579 & n73774) | (n63750 & n73774);
  assign n73776 = (n63750 & n73701) | (n63750 & n73774) | (n73701 & n73774);
  assign n73777 = (n63280 & n73775) | (n63280 & n73776) | (n73775 & n73776);
  assign n45340 = ~n73773 & n73777;
  assign n45341 = x174 & x208;
  assign n45342 = n45340 & n45341;
  assign n45343 = n45340 | n45341;
  assign n45344 = ~n45342 & n45343;
  assign n63752 = n45077 & n45344;
  assign n63753 = (n45344 & n63595) | (n45344 & n63752) | (n63595 & n63752);
  assign n63754 = n45077 | n45344;
  assign n63755 = n63595 | n63754;
  assign n45347 = ~n63753 & n63755;
  assign n45348 = x173 & x209;
  assign n45349 = n45347 & n45348;
  assign n45350 = n45347 | n45348;
  assign n45351 = ~n45349 & n45350;
  assign n45352 = n73758 & n45351;
  assign n45353 = n73758 | n45351;
  assign n45354 = ~n45352 & n45353;
  assign n45355 = x172 & x210;
  assign n45356 = n45354 & n45355;
  assign n45357 = n45354 | n45355;
  assign n45358 = ~n45356 & n45357;
  assign n63730 = n45091 | n45093;
  assign n63756 = n45358 & n63730;
  assign n63757 = n45091 & n45358;
  assign n63758 = (n63575 & n63756) | (n63575 & n63757) | (n63756 & n63757);
  assign n63759 = n45358 | n63730;
  assign n63760 = n45091 | n45358;
  assign n63761 = (n63575 & n63759) | (n63575 & n63760) | (n63759 & n63760);
  assign n45361 = ~n63758 & n63761;
  assign n45362 = x171 & x211;
  assign n45363 = n45361 & n45362;
  assign n45364 = n45361 | n45362;
  assign n45365 = ~n45363 & n45364;
  assign n63762 = n45098 & n45365;
  assign n63763 = (n45365 & n63605) | (n45365 & n63762) | (n63605 & n63762);
  assign n63764 = n45098 | n45365;
  assign n63765 = n63605 | n63764;
  assign n45368 = ~n63763 & n63765;
  assign n45369 = x170 & x212;
  assign n45370 = n45368 & n45369;
  assign n45371 = n45368 | n45369;
  assign n45372 = ~n45370 & n45371;
  assign n45373 = n73753 & n45372;
  assign n45374 = n73753 | n45372;
  assign n45375 = ~n45373 & n45374;
  assign n45376 = x169 & x213;
  assign n45377 = n45375 & n45376;
  assign n45378 = n45375 | n45376;
  assign n45379 = ~n45377 & n45378;
  assign n63725 = n45112 | n45114;
  assign n63766 = n45379 & n63725;
  assign n63767 = n45112 & n45379;
  assign n63768 = (n73697 & n63766) | (n73697 & n63767) | (n63766 & n63767);
  assign n63769 = n45379 | n63725;
  assign n63770 = n45112 | n45379;
  assign n63771 = (n73697 & n63769) | (n73697 & n63770) | (n63769 & n63770);
  assign n45382 = ~n63768 & n63771;
  assign n45383 = x168 & x214;
  assign n45384 = n45382 & n45383;
  assign n45385 = n45382 | n45383;
  assign n45386 = ~n45384 & n45385;
  assign n63772 = n45119 & n45386;
  assign n73778 = (n45386 & n63614) | (n45386 & n63772) | (n63614 & n63772);
  assign n73779 = (n45386 & n63613) | (n45386 & n63772) | (n63613 & n63772);
  assign n73780 = (n73636 & n73778) | (n73636 & n73779) | (n73778 & n73779);
  assign n63774 = n45119 | n45386;
  assign n73781 = n63614 | n63774;
  assign n73782 = n63613 | n63774;
  assign n73783 = (n73636 & n73781) | (n73636 & n73782) | (n73781 & n73782);
  assign n45389 = ~n73780 & n73783;
  assign n45390 = x167 & x215;
  assign n45391 = n45389 & n45390;
  assign n45392 = n45389 | n45390;
  assign n45393 = ~n45391 & n45392;
  assign n45394 = n73748 & n45393;
  assign n45395 = n73748 | n45393;
  assign n45396 = ~n45394 & n45395;
  assign n45397 = x166 & x216;
  assign n45398 = n45396 & n45397;
  assign n45399 = n45396 | n45397;
  assign n45400 = ~n45398 & n45399;
  assign n63720 = n45133 | n45135;
  assign n63776 = n45400 & n63720;
  assign n63777 = n45133 & n45400;
  assign n63778 = (n73692 & n63776) | (n73692 & n63777) | (n63776 & n63777);
  assign n63779 = n45400 | n63720;
  assign n63780 = n45133 | n45400;
  assign n63781 = (n73692 & n63779) | (n73692 & n63780) | (n63779 & n63780);
  assign n45403 = ~n63778 & n63781;
  assign n45404 = x165 & x217;
  assign n45405 = n45403 & n45404;
  assign n45406 = n45403 | n45404;
  assign n45407 = ~n45405 & n45406;
  assign n63782 = n45140 & n45407;
  assign n73784 = (n45407 & n63624) | (n45407 & n63782) | (n63624 & n63782);
  assign n73785 = (n45407 & n63623) | (n45407 & n63782) | (n63623 & n63782);
  assign n73786 = (n63408 & n73784) | (n63408 & n73785) | (n73784 & n73785);
  assign n63784 = n45140 | n45407;
  assign n73787 = n63624 | n63784;
  assign n73788 = n63623 | n63784;
  assign n73789 = (n63408 & n73787) | (n63408 & n73788) | (n73787 & n73788);
  assign n45410 = ~n73786 & n73789;
  assign n45411 = x164 & x218;
  assign n45412 = n45410 & n45411;
  assign n45413 = n45410 | n45411;
  assign n45414 = ~n45412 & n45413;
  assign n63718 = n45147 | n45149;
  assign n73790 = n45414 & n63718;
  assign n73742 = n44874 | n45147;
  assign n73743 = (n45147 & n45149) | (n45147 & n73742) | (n45149 & n73742);
  assign n73791 = n45414 & n73743;
  assign n73792 = (n73684 & n73790) | (n73684 & n73791) | (n73790 & n73791);
  assign n73793 = n45414 | n63718;
  assign n73794 = n45414 | n73743;
  assign n73795 = (n73684 & n73793) | (n73684 & n73794) | (n73793 & n73794);
  assign n45417 = ~n73792 & n73795;
  assign n45418 = x163 & x219;
  assign n45419 = n45417 & n45418;
  assign n45420 = n45417 | n45418;
  assign n45421 = ~n45419 & n45420;
  assign n63786 = n45154 & n45421;
  assign n73796 = (n45421 & n63633) | (n45421 & n63786) | (n63633 & n63786);
  assign n73797 = (n45156 & n45421) | (n45156 & n63786) | (n45421 & n63786);
  assign n73798 = (n63478 & n73796) | (n63478 & n73797) | (n73796 & n73797);
  assign n63788 = n45154 | n45421;
  assign n73799 = n63633 | n63788;
  assign n73800 = n45156 | n63788;
  assign n73801 = (n63478 & n73799) | (n63478 & n73800) | (n73799 & n73800);
  assign n45424 = ~n73798 & n73801;
  assign n45425 = x162 & x220;
  assign n45426 = n45424 & n45425;
  assign n45427 = n45424 | n45425;
  assign n45428 = ~n45426 & n45427;
  assign n63790 = n45161 & n45428;
  assign n63791 = (n45428 & n63638) | (n45428 & n63790) | (n63638 & n63790);
  assign n63792 = n45161 | n45428;
  assign n63793 = n63638 | n63792;
  assign n45431 = ~n63791 & n63793;
  assign n45432 = x161 & x221;
  assign n45433 = n45431 & n45432;
  assign n45434 = n45431 | n45432;
  assign n45435 = ~n45433 & n45434;
  assign n63794 = n45168 & n45435;
  assign n63795 = (n45435 & n63642) | (n45435 & n63794) | (n63642 & n63794);
  assign n63796 = n45168 | n45435;
  assign n63797 = n63642 | n63796;
  assign n45438 = ~n63795 & n63797;
  assign n45439 = x160 & x222;
  assign n45440 = n45438 & n45439;
  assign n45441 = n45438 | n45439;
  assign n45442 = ~n45440 & n45441;
  assign n63798 = n45175 & n45442;
  assign n63799 = (n45442 & n63646) | (n45442 & n63798) | (n63646 & n63798);
  assign n63800 = n45175 | n45442;
  assign n63801 = n63646 | n63800;
  assign n45445 = ~n63799 & n63801;
  assign n45446 = x159 & x223;
  assign n45447 = n45445 & n45446;
  assign n45448 = n45445 | n45446;
  assign n45449 = ~n45447 & n45448;
  assign n63802 = n45182 & n45449;
  assign n63803 = (n45449 & n63650) | (n45449 & n63802) | (n63650 & n63802);
  assign n63804 = n45182 | n45449;
  assign n63805 = n63650 | n63804;
  assign n45452 = ~n63803 & n63805;
  assign n45453 = x158 & x224;
  assign n45454 = n45452 & n45453;
  assign n45455 = n45452 | n45453;
  assign n45456 = ~n45454 & n45455;
  assign n63806 = n45189 & n45456;
  assign n63807 = (n45456 & n63654) | (n45456 & n63806) | (n63654 & n63806);
  assign n63808 = n45189 | n45456;
  assign n63809 = n63654 | n63808;
  assign n45459 = ~n63807 & n63809;
  assign n45460 = x157 & x225;
  assign n45461 = n45459 & n45460;
  assign n45462 = n45459 | n45460;
  assign n45463 = ~n45461 & n45462;
  assign n63810 = n45196 & n45463;
  assign n63811 = (n45463 & n63658) | (n45463 & n63810) | (n63658 & n63810);
  assign n63812 = n45196 | n45463;
  assign n63813 = n63658 | n63812;
  assign n45466 = ~n63811 & n63813;
  assign n45467 = x156 & x226;
  assign n45468 = n45466 & n45467;
  assign n45469 = n45466 | n45467;
  assign n45470 = ~n45468 & n45469;
  assign n63814 = n45203 & n45470;
  assign n63815 = (n45470 & n63662) | (n45470 & n63814) | (n63662 & n63814);
  assign n63816 = n45203 | n45470;
  assign n63817 = n63662 | n63816;
  assign n45473 = ~n63815 & n63817;
  assign n45474 = x155 & x227;
  assign n45475 = n45473 & n45474;
  assign n45476 = n45473 | n45474;
  assign n45477 = ~n45475 & n45476;
  assign n63818 = n45210 & n45477;
  assign n63819 = (n45477 & n63666) | (n45477 & n63818) | (n63666 & n63818);
  assign n63820 = n45210 | n45477;
  assign n63821 = n63666 | n63820;
  assign n45480 = ~n63819 & n63821;
  assign n45481 = x154 & x228;
  assign n45482 = n45480 & n45481;
  assign n45483 = n45480 | n45481;
  assign n45484 = ~n45482 & n45483;
  assign n63822 = n45217 & n45484;
  assign n63823 = (n45484 & n63670) | (n45484 & n63822) | (n63670 & n63822);
  assign n63824 = n45217 | n45484;
  assign n63825 = n63670 | n63824;
  assign n45487 = ~n63823 & n63825;
  assign n45488 = x153 & x229;
  assign n45489 = n45487 & n45488;
  assign n45490 = n45487 | n45488;
  assign n45491 = ~n45489 & n45490;
  assign n63826 = n45224 & n45491;
  assign n63827 = (n45491 & n63674) | (n45491 & n63826) | (n63674 & n63826);
  assign n63828 = n45224 | n45491;
  assign n63829 = n63674 | n63828;
  assign n45494 = ~n63827 & n63829;
  assign n45495 = x152 & x230;
  assign n45496 = n45494 & n45495;
  assign n45497 = n45494 | n45495;
  assign n45498 = ~n45496 & n45497;
  assign n63830 = n45231 & n45498;
  assign n63831 = (n45498 & n63678) | (n45498 & n63830) | (n63678 & n63830);
  assign n63832 = n45231 | n45498;
  assign n63833 = n63678 | n63832;
  assign n45501 = ~n63831 & n63833;
  assign n45502 = x151 & x231;
  assign n45503 = n45501 & n45502;
  assign n45504 = n45501 | n45502;
  assign n45505 = ~n45503 & n45504;
  assign n63834 = n45238 & n45505;
  assign n63835 = (n45505 & n63682) | (n45505 & n63834) | (n63682 & n63834);
  assign n63836 = n45238 | n45505;
  assign n63837 = n63682 | n63836;
  assign n45508 = ~n63835 & n63837;
  assign n45509 = x150 & x232;
  assign n45510 = n45508 & n45509;
  assign n45511 = n45508 | n45509;
  assign n45512 = ~n45510 & n45511;
  assign n63838 = n45245 & n45512;
  assign n63839 = (n45512 & n63686) | (n45512 & n63838) | (n63686 & n63838);
  assign n63840 = n45245 | n45512;
  assign n63841 = n63686 | n63840;
  assign n45515 = ~n63839 & n63841;
  assign n45516 = x149 & x233;
  assign n45517 = n45515 & n45516;
  assign n45518 = n45515 | n45516;
  assign n45519 = ~n45517 & n45518;
  assign n63842 = n45252 & n45519;
  assign n63843 = (n45519 & n63690) | (n45519 & n63842) | (n63690 & n63842);
  assign n63844 = n45252 | n45519;
  assign n63845 = n63690 | n63844;
  assign n45522 = ~n63843 & n63845;
  assign n45523 = x148 & x234;
  assign n45524 = n45522 & n45523;
  assign n45525 = n45522 | n45523;
  assign n45526 = ~n45524 & n45525;
  assign n63846 = n45259 & n45526;
  assign n63847 = (n45526 & n63694) | (n45526 & n63846) | (n63694 & n63846);
  assign n63848 = n45259 | n45526;
  assign n63849 = n63694 | n63848;
  assign n45529 = ~n63847 & n63849;
  assign n45530 = x147 & x235;
  assign n45531 = n45529 & n45530;
  assign n45532 = n45529 | n45530;
  assign n45533 = ~n45531 & n45532;
  assign n63850 = n45266 & n45533;
  assign n63851 = (n45533 & n63698) | (n45533 & n63850) | (n63698 & n63850);
  assign n63852 = n45266 | n45533;
  assign n63853 = n63698 | n63852;
  assign n45536 = ~n63851 & n63853;
  assign n45537 = x146 & x236;
  assign n45538 = n45536 & n45537;
  assign n45539 = n45536 | n45537;
  assign n45540 = ~n45538 & n45539;
  assign n63854 = n45273 & n45540;
  assign n63855 = (n45540 & n63702) | (n45540 & n63854) | (n63702 & n63854);
  assign n63856 = n45273 | n45540;
  assign n63857 = n63702 | n63856;
  assign n45543 = ~n63855 & n63857;
  assign n45544 = x145 & x237;
  assign n45545 = n45543 & n45544;
  assign n45546 = n45543 | n45544;
  assign n45547 = ~n45545 & n45546;
  assign n63858 = n45280 & n45547;
  assign n63859 = (n45547 & n63706) | (n45547 & n63858) | (n63706 & n63858);
  assign n63860 = n45280 | n45547;
  assign n63861 = n63706 | n63860;
  assign n45550 = ~n63859 & n63861;
  assign n45551 = x144 & x238;
  assign n45552 = n45550 & n45551;
  assign n45553 = n45550 | n45551;
  assign n45554 = ~n45552 & n45553;
  assign n63862 = n45287 & n45554;
  assign n63863 = (n45554 & n63710) | (n45554 & n63862) | (n63710 & n63862);
  assign n63864 = n45287 | n45554;
  assign n63865 = n63710 | n63864;
  assign n45557 = ~n63863 & n63865;
  assign n45558 = x143 & x239;
  assign n45559 = n45557 & n45558;
  assign n45560 = n45557 | n45558;
  assign n45561 = ~n45559 & n45560;
  assign n63866 = n45294 & n45561;
  assign n63867 = (n45561 & n63714) | (n45561 & n63866) | (n63714 & n63866);
  assign n63868 = n45294 | n45561;
  assign n63869 = n63714 | n63868;
  assign n45564 = ~n63867 & n63869;
  assign n63719 = (n73684 & n73743) | (n73684 & n63718) | (n73743 & n63718);
  assign n63873 = n45405 | n45407;
  assign n73802 = n45140 | n45405;
  assign n73803 = (n45405 & n45407) | (n45405 & n73802) | (n45407 & n73802);
  assign n73804 = (n63624 & n63873) | (n63624 & n73803) | (n63873 & n73803);
  assign n73805 = (n63623 & n63873) | (n63623 & n73803) | (n63873 & n73803);
  assign n73806 = (n63408 & n73804) | (n63408 & n73805) | (n73804 & n73805);
  assign n63878 = n45384 | n45386;
  assign n73807 = n45119 | n45384;
  assign n73808 = (n45384 & n45386) | (n45384 & n73807) | (n45386 & n73807);
  assign n73809 = (n63614 & n63878) | (n63614 & n73808) | (n63878 & n73808);
  assign n73810 = (n63613 & n63878) | (n63613 & n73808) | (n63878 & n73808);
  assign n73811 = (n73636 & n73809) | (n73636 & n73810) | (n73809 & n73810);
  assign n45598 = x175 & x208;
  assign n63890 = n45598 & n73764;
  assign n63891 = (n45598 & n73773) | (n45598 & n63890) | (n73773 & n63890);
  assign n63892 = n45598 | n73764;
  assign n63893 = n73773 | n63892;
  assign n45601 = ~n63891 & n63893;
  assign n63888 = n45342 | n45344;
  assign n73816 = n45601 & n63888;
  assign n73814 = n45077 | n45342;
  assign n73815 = (n45342 & n45344) | (n45342 & n73814) | (n45344 & n73814);
  assign n73817 = n45601 & n73815;
  assign n73818 = (n63595 & n73816) | (n63595 & n73817) | (n73816 & n73817);
  assign n73819 = n45601 | n63888;
  assign n73820 = n45601 | n73815;
  assign n73821 = (n63595 & n73819) | (n63595 & n73820) | (n73819 & n73820);
  assign n45604 = ~n73818 & n73821;
  assign n45605 = x174 & x209;
  assign n45606 = n45604 & n45605;
  assign n45607 = n45604 | n45605;
  assign n45608 = ~n45606 & n45607;
  assign n63885 = n45349 | n45351;
  assign n63894 = n45608 & n63885;
  assign n63895 = n45349 & n45608;
  assign n63896 = (n73758 & n63894) | (n73758 & n63895) | (n63894 & n63895);
  assign n63897 = n45608 | n63885;
  assign n63898 = n45349 | n45608;
  assign n63899 = (n73758 & n63897) | (n73758 & n63898) | (n63897 & n63898);
  assign n45611 = ~n63896 & n63899;
  assign n45612 = x173 & x210;
  assign n45613 = n45611 & n45612;
  assign n45614 = n45611 | n45612;
  assign n45615 = ~n45613 & n45614;
  assign n63900 = n45356 & n45615;
  assign n73822 = (n45615 & n63757) | (n45615 & n63900) | (n63757 & n63900);
  assign n73823 = (n45615 & n63756) | (n45615 & n63900) | (n63756 & n63900);
  assign n73824 = (n63575 & n73822) | (n63575 & n73823) | (n73822 & n73823);
  assign n63902 = n45356 | n45615;
  assign n73825 = n63757 | n63902;
  assign n73826 = n63756 | n63902;
  assign n73827 = (n63575 & n73825) | (n63575 & n73826) | (n73825 & n73826);
  assign n45618 = ~n73824 & n73827;
  assign n45619 = x172 & x211;
  assign n45620 = n45618 & n45619;
  assign n45621 = n45618 | n45619;
  assign n45622 = ~n45620 & n45621;
  assign n63883 = n45363 | n45365;
  assign n73828 = n45622 & n63883;
  assign n73812 = n45098 | n45363;
  assign n73813 = (n45363 & n45365) | (n45363 & n73812) | (n45365 & n73812);
  assign n73829 = n45622 & n73813;
  assign n73830 = (n63605 & n73828) | (n63605 & n73829) | (n73828 & n73829);
  assign n73831 = n45622 | n63883;
  assign n73832 = n45622 | n73813;
  assign n73833 = (n63605 & n73831) | (n63605 & n73832) | (n73831 & n73832);
  assign n45625 = ~n73830 & n73833;
  assign n45626 = x171 & x212;
  assign n45627 = n45625 & n45626;
  assign n45628 = n45625 | n45626;
  assign n45629 = ~n45627 & n45628;
  assign n63880 = n45370 | n45372;
  assign n63904 = n45629 & n63880;
  assign n63905 = n45370 & n45629;
  assign n63906 = (n73753 & n63904) | (n73753 & n63905) | (n63904 & n63905);
  assign n63907 = n45629 | n63880;
  assign n63908 = n45370 | n45629;
  assign n63909 = (n73753 & n63907) | (n73753 & n63908) | (n63907 & n63908);
  assign n45632 = ~n63906 & n63909;
  assign n45633 = x170 & x213;
  assign n45634 = n45632 & n45633;
  assign n45635 = n45632 | n45633;
  assign n45636 = ~n45634 & n45635;
  assign n63910 = n45377 & n45636;
  assign n73834 = (n45636 & n63767) | (n45636 & n63910) | (n63767 & n63910);
  assign n73835 = (n45636 & n63766) | (n45636 & n63910) | (n63766 & n63910);
  assign n73836 = (n73697 & n73834) | (n73697 & n73835) | (n73834 & n73835);
  assign n63912 = n45377 | n45636;
  assign n73837 = n63767 | n63912;
  assign n73838 = n63766 | n63912;
  assign n73839 = (n73697 & n73837) | (n73697 & n73838) | (n73837 & n73838);
  assign n45639 = ~n73836 & n73839;
  assign n45640 = x169 & x214;
  assign n45641 = n45639 & n45640;
  assign n45642 = n45639 | n45640;
  assign n45643 = ~n45641 & n45642;
  assign n45644 = n73811 & n45643;
  assign n45645 = n73811 | n45643;
  assign n45646 = ~n45644 & n45645;
  assign n45647 = x168 & x215;
  assign n45648 = n45646 & n45647;
  assign n45649 = n45646 | n45647;
  assign n45650 = ~n45648 & n45649;
  assign n63875 = n45391 | n45393;
  assign n63914 = n45650 & n63875;
  assign n63915 = n45391 & n45650;
  assign n63916 = (n73748 & n63914) | (n73748 & n63915) | (n63914 & n63915);
  assign n63917 = n45650 | n63875;
  assign n63918 = n45391 | n45650;
  assign n63919 = (n73748 & n63917) | (n73748 & n63918) | (n63917 & n63918);
  assign n45653 = ~n63916 & n63919;
  assign n45654 = x167 & x216;
  assign n45655 = n45653 & n45654;
  assign n45656 = n45653 | n45654;
  assign n45657 = ~n45655 & n45656;
  assign n63920 = n45398 & n45657;
  assign n73840 = (n45657 & n63777) | (n45657 & n63920) | (n63777 & n63920);
  assign n73841 = (n45657 & n63776) | (n45657 & n63920) | (n63776 & n63920);
  assign n73842 = (n73692 & n73840) | (n73692 & n73841) | (n73840 & n73841);
  assign n63922 = n45398 | n45657;
  assign n73843 = n63777 | n63922;
  assign n73844 = n63776 | n63922;
  assign n73845 = (n73692 & n73843) | (n73692 & n73844) | (n73843 & n73844);
  assign n45660 = ~n73842 & n73845;
  assign n45661 = x166 & x217;
  assign n45662 = n45660 & n45661;
  assign n45663 = n45660 | n45661;
  assign n45664 = ~n45662 & n45663;
  assign n45665 = n73806 & n45664;
  assign n45666 = n73806 | n45664;
  assign n45667 = ~n45665 & n45666;
  assign n45668 = x165 & x218;
  assign n45669 = n45667 & n45668;
  assign n45670 = n45667 | n45668;
  assign n45671 = ~n45669 & n45670;
  assign n63870 = n45412 | n45414;
  assign n63924 = n45671 & n63870;
  assign n63925 = n45412 & n45671;
  assign n63926 = (n63719 & n63924) | (n63719 & n63925) | (n63924 & n63925);
  assign n63927 = n45671 | n63870;
  assign n63928 = n45412 | n45671;
  assign n63929 = (n63719 & n63927) | (n63719 & n63928) | (n63927 & n63928);
  assign n45674 = ~n63926 & n63929;
  assign n45675 = x164 & x219;
  assign n45676 = n45674 & n45675;
  assign n45677 = n45674 | n45675;
  assign n45678 = ~n45676 & n45677;
  assign n63930 = n45419 & n45678;
  assign n63931 = (n45678 & n73798) | (n45678 & n63930) | (n73798 & n63930);
  assign n63932 = n45419 | n45678;
  assign n63933 = n73798 | n63932;
  assign n45681 = ~n63931 & n63933;
  assign n45682 = x163 & x220;
  assign n45683 = n45681 & n45682;
  assign n45684 = n45681 | n45682;
  assign n45685 = ~n45683 & n45684;
  assign n63934 = n45426 & n45685;
  assign n63935 = (n45685 & n63791) | (n45685 & n63934) | (n63791 & n63934);
  assign n63936 = n45426 | n45685;
  assign n63937 = n63791 | n63936;
  assign n45688 = ~n63935 & n63937;
  assign n45689 = x162 & x221;
  assign n45690 = n45688 & n45689;
  assign n45691 = n45688 | n45689;
  assign n45692 = ~n45690 & n45691;
  assign n63938 = n45433 & n45692;
  assign n63939 = (n45692 & n63795) | (n45692 & n63938) | (n63795 & n63938);
  assign n63940 = n45433 | n45692;
  assign n63941 = n63795 | n63940;
  assign n45695 = ~n63939 & n63941;
  assign n45696 = x161 & x222;
  assign n45697 = n45695 & n45696;
  assign n45698 = n45695 | n45696;
  assign n45699 = ~n45697 & n45698;
  assign n63942 = n45440 & n45699;
  assign n63943 = (n45699 & n63799) | (n45699 & n63942) | (n63799 & n63942);
  assign n63944 = n45440 | n45699;
  assign n63945 = n63799 | n63944;
  assign n45702 = ~n63943 & n63945;
  assign n45703 = x160 & x223;
  assign n45704 = n45702 & n45703;
  assign n45705 = n45702 | n45703;
  assign n45706 = ~n45704 & n45705;
  assign n63946 = n45447 & n45706;
  assign n63947 = (n45706 & n63803) | (n45706 & n63946) | (n63803 & n63946);
  assign n63948 = n45447 | n45706;
  assign n63949 = n63803 | n63948;
  assign n45709 = ~n63947 & n63949;
  assign n45710 = x159 & x224;
  assign n45711 = n45709 & n45710;
  assign n45712 = n45709 | n45710;
  assign n45713 = ~n45711 & n45712;
  assign n63950 = n45454 & n45713;
  assign n63951 = (n45713 & n63807) | (n45713 & n63950) | (n63807 & n63950);
  assign n63952 = n45454 | n45713;
  assign n63953 = n63807 | n63952;
  assign n45716 = ~n63951 & n63953;
  assign n45717 = x158 & x225;
  assign n45718 = n45716 & n45717;
  assign n45719 = n45716 | n45717;
  assign n45720 = ~n45718 & n45719;
  assign n63954 = n45461 & n45720;
  assign n63955 = (n45720 & n63811) | (n45720 & n63954) | (n63811 & n63954);
  assign n63956 = n45461 | n45720;
  assign n63957 = n63811 | n63956;
  assign n45723 = ~n63955 & n63957;
  assign n45724 = x157 & x226;
  assign n45725 = n45723 & n45724;
  assign n45726 = n45723 | n45724;
  assign n45727 = ~n45725 & n45726;
  assign n63958 = n45468 & n45727;
  assign n63959 = (n45727 & n63815) | (n45727 & n63958) | (n63815 & n63958);
  assign n63960 = n45468 | n45727;
  assign n63961 = n63815 | n63960;
  assign n45730 = ~n63959 & n63961;
  assign n45731 = x156 & x227;
  assign n45732 = n45730 & n45731;
  assign n45733 = n45730 | n45731;
  assign n45734 = ~n45732 & n45733;
  assign n63962 = n45475 & n45734;
  assign n63963 = (n45734 & n63819) | (n45734 & n63962) | (n63819 & n63962);
  assign n63964 = n45475 | n45734;
  assign n63965 = n63819 | n63964;
  assign n45737 = ~n63963 & n63965;
  assign n45738 = x155 & x228;
  assign n45739 = n45737 & n45738;
  assign n45740 = n45737 | n45738;
  assign n45741 = ~n45739 & n45740;
  assign n63966 = n45482 & n45741;
  assign n63967 = (n45741 & n63823) | (n45741 & n63966) | (n63823 & n63966);
  assign n63968 = n45482 | n45741;
  assign n63969 = n63823 | n63968;
  assign n45744 = ~n63967 & n63969;
  assign n45745 = x154 & x229;
  assign n45746 = n45744 & n45745;
  assign n45747 = n45744 | n45745;
  assign n45748 = ~n45746 & n45747;
  assign n63970 = n45489 & n45748;
  assign n63971 = (n45748 & n63827) | (n45748 & n63970) | (n63827 & n63970);
  assign n63972 = n45489 | n45748;
  assign n63973 = n63827 | n63972;
  assign n45751 = ~n63971 & n63973;
  assign n45752 = x153 & x230;
  assign n45753 = n45751 & n45752;
  assign n45754 = n45751 | n45752;
  assign n45755 = ~n45753 & n45754;
  assign n63974 = n45496 & n45755;
  assign n63975 = (n45755 & n63831) | (n45755 & n63974) | (n63831 & n63974);
  assign n63976 = n45496 | n45755;
  assign n63977 = n63831 | n63976;
  assign n45758 = ~n63975 & n63977;
  assign n45759 = x152 & x231;
  assign n45760 = n45758 & n45759;
  assign n45761 = n45758 | n45759;
  assign n45762 = ~n45760 & n45761;
  assign n63978 = n45503 & n45762;
  assign n63979 = (n45762 & n63835) | (n45762 & n63978) | (n63835 & n63978);
  assign n63980 = n45503 | n45762;
  assign n63981 = n63835 | n63980;
  assign n45765 = ~n63979 & n63981;
  assign n45766 = x151 & x232;
  assign n45767 = n45765 & n45766;
  assign n45768 = n45765 | n45766;
  assign n45769 = ~n45767 & n45768;
  assign n63982 = n45510 & n45769;
  assign n63983 = (n45769 & n63839) | (n45769 & n63982) | (n63839 & n63982);
  assign n63984 = n45510 | n45769;
  assign n63985 = n63839 | n63984;
  assign n45772 = ~n63983 & n63985;
  assign n45773 = x150 & x233;
  assign n45774 = n45772 & n45773;
  assign n45775 = n45772 | n45773;
  assign n45776 = ~n45774 & n45775;
  assign n63986 = n45517 & n45776;
  assign n63987 = (n45776 & n63843) | (n45776 & n63986) | (n63843 & n63986);
  assign n63988 = n45517 | n45776;
  assign n63989 = n63843 | n63988;
  assign n45779 = ~n63987 & n63989;
  assign n45780 = x149 & x234;
  assign n45781 = n45779 & n45780;
  assign n45782 = n45779 | n45780;
  assign n45783 = ~n45781 & n45782;
  assign n63990 = n45524 & n45783;
  assign n63991 = (n45783 & n63847) | (n45783 & n63990) | (n63847 & n63990);
  assign n63992 = n45524 | n45783;
  assign n63993 = n63847 | n63992;
  assign n45786 = ~n63991 & n63993;
  assign n45787 = x148 & x235;
  assign n45788 = n45786 & n45787;
  assign n45789 = n45786 | n45787;
  assign n45790 = ~n45788 & n45789;
  assign n63994 = n45531 & n45790;
  assign n63995 = (n45790 & n63851) | (n45790 & n63994) | (n63851 & n63994);
  assign n63996 = n45531 | n45790;
  assign n63997 = n63851 | n63996;
  assign n45793 = ~n63995 & n63997;
  assign n45794 = x147 & x236;
  assign n45795 = n45793 & n45794;
  assign n45796 = n45793 | n45794;
  assign n45797 = ~n45795 & n45796;
  assign n63998 = n45538 & n45797;
  assign n63999 = (n45797 & n63855) | (n45797 & n63998) | (n63855 & n63998);
  assign n64000 = n45538 | n45797;
  assign n64001 = n63855 | n64000;
  assign n45800 = ~n63999 & n64001;
  assign n45801 = x146 & x237;
  assign n45802 = n45800 & n45801;
  assign n45803 = n45800 | n45801;
  assign n45804 = ~n45802 & n45803;
  assign n64002 = n45545 & n45804;
  assign n64003 = (n45804 & n63859) | (n45804 & n64002) | (n63859 & n64002);
  assign n64004 = n45545 | n45804;
  assign n64005 = n63859 | n64004;
  assign n45807 = ~n64003 & n64005;
  assign n45808 = x145 & x238;
  assign n45809 = n45807 & n45808;
  assign n45810 = n45807 | n45808;
  assign n45811 = ~n45809 & n45810;
  assign n64006 = n45552 & n45811;
  assign n64007 = (n45811 & n63863) | (n45811 & n64006) | (n63863 & n64006);
  assign n64008 = n45552 | n45811;
  assign n64009 = n63863 | n64008;
  assign n45814 = ~n64007 & n64009;
  assign n45815 = x144 & x239;
  assign n45816 = n45814 & n45815;
  assign n45817 = n45814 | n45815;
  assign n45818 = ~n45816 & n45817;
  assign n64010 = n45559 & n45818;
  assign n64011 = (n45818 & n63867) | (n45818 & n64010) | (n63867 & n64010);
  assign n64012 = n45559 | n45818;
  assign n64013 = n63867 | n64012;
  assign n45821 = ~n64011 & n64013;
  assign n64020 = n45655 | n45657;
  assign n73848 = n45398 | n45655;
  assign n73849 = (n45655 & n45657) | (n45655 & n73848) | (n45657 & n73848);
  assign n73850 = (n63777 & n64020) | (n63777 & n73849) | (n64020 & n73849);
  assign n73851 = (n63776 & n64020) | (n63776 & n73849) | (n64020 & n73849);
  assign n73852 = (n73692 & n73850) | (n73692 & n73851) | (n73850 & n73851);
  assign n64025 = n45634 | n45636;
  assign n73853 = n45377 | n45634;
  assign n73854 = (n45634 & n45636) | (n45634 & n73853) | (n45636 & n73853);
  assign n73855 = (n63767 & n64025) | (n63767 & n73854) | (n64025 & n73854);
  assign n73856 = (n63766 & n64025) | (n63766 & n73854) | (n64025 & n73854);
  assign n73857 = (n73697 & n73855) | (n73697 & n73856) | (n73855 & n73856);
  assign n63884 = (n63605 & n73813) | (n63605 & n63883) | (n73813 & n63883);
  assign n64030 = n45613 | n45615;
  assign n73858 = n45356 | n45613;
  assign n73859 = (n45613 & n45615) | (n45613 & n73858) | (n45615 & n73858);
  assign n73860 = (n63757 & n64030) | (n63757 & n73859) | (n64030 & n73859);
  assign n73861 = (n63756 & n64030) | (n63756 & n73859) | (n64030 & n73859);
  assign n73862 = (n63575 & n73860) | (n63575 & n73861) | (n73860 & n73861);
  assign n45854 = x175 & x209;
  assign n73864 = n45854 & n63890;
  assign n73865 = n45598 & n45854;
  assign n73866 = (n73773 & n73864) | (n73773 & n73865) | (n73864 & n73865);
  assign n73863 = (n45601 & n45854) | (n45601 & n73866) | (n45854 & n73866);
  assign n73867 = (n63888 & n73863) | (n63888 & n73866) | (n73863 & n73866);
  assign n73868 = (n73815 & n73863) | (n73815 & n73866) | (n73863 & n73866);
  assign n73869 = (n63595 & n73867) | (n63595 & n73868) | (n73867 & n73868);
  assign n73871 = n45854 | n63890;
  assign n73872 = n45598 | n45854;
  assign n73873 = (n73773 & n73871) | (n73773 & n73872) | (n73871 & n73872);
  assign n73870 = n45601 | n73873;
  assign n73874 = (n63888 & n73870) | (n63888 & n73873) | (n73870 & n73873);
  assign n73875 = (n73815 & n73870) | (n73815 & n73873) | (n73870 & n73873);
  assign n73876 = (n63595 & n73874) | (n63595 & n73875) | (n73874 & n73875);
  assign n45857 = ~n73869 & n73876;
  assign n64040 = n45606 & n45857;
  assign n64041 = (n45857 & n63896) | (n45857 & n64040) | (n63896 & n64040);
  assign n64042 = n45606 | n45857;
  assign n64043 = n63896 | n64042;
  assign n45860 = ~n64041 & n64043;
  assign n45861 = x174 & x210;
  assign n45862 = n45860 & n45861;
  assign n45863 = n45860 | n45861;
  assign n45864 = ~n45862 & n45863;
  assign n45865 = n73862 & n45864;
  assign n45866 = n73862 | n45864;
  assign n45867 = ~n45865 & n45866;
  assign n45868 = x173 & x211;
  assign n45869 = n45867 & n45868;
  assign n45870 = n45867 | n45868;
  assign n45871 = ~n45869 & n45870;
  assign n64027 = n45620 | n45622;
  assign n64044 = n45871 & n64027;
  assign n64045 = n45620 & n45871;
  assign n64046 = (n63884 & n64044) | (n63884 & n64045) | (n64044 & n64045);
  assign n64047 = n45871 | n64027;
  assign n64048 = n45620 | n45871;
  assign n64049 = (n63884 & n64047) | (n63884 & n64048) | (n64047 & n64048);
  assign n45874 = ~n64046 & n64049;
  assign n45875 = x172 & x212;
  assign n45876 = n45874 & n45875;
  assign n45877 = n45874 | n45875;
  assign n45878 = ~n45876 & n45877;
  assign n64050 = n45627 & n45878;
  assign n64051 = (n45878 & n63906) | (n45878 & n64050) | (n63906 & n64050);
  assign n64052 = n45627 | n45878;
  assign n64053 = n63906 | n64052;
  assign n45881 = ~n64051 & n64053;
  assign n45882 = x171 & x213;
  assign n45883 = n45881 & n45882;
  assign n45884 = n45881 | n45882;
  assign n45885 = ~n45883 & n45884;
  assign n45886 = n73857 & n45885;
  assign n45887 = n73857 | n45885;
  assign n45888 = ~n45886 & n45887;
  assign n45889 = x170 & x214;
  assign n45890 = n45888 & n45889;
  assign n45891 = n45888 | n45889;
  assign n45892 = ~n45890 & n45891;
  assign n64022 = n45641 | n45643;
  assign n64054 = n45892 & n64022;
  assign n64055 = n45641 & n45892;
  assign n64056 = (n73811 & n64054) | (n73811 & n64055) | (n64054 & n64055);
  assign n64057 = n45892 | n64022;
  assign n64058 = n45641 | n45892;
  assign n64059 = (n73811 & n64057) | (n73811 & n64058) | (n64057 & n64058);
  assign n45895 = ~n64056 & n64059;
  assign n45896 = x169 & x215;
  assign n45897 = n45895 & n45896;
  assign n45898 = n45895 | n45896;
  assign n45899 = ~n45897 & n45898;
  assign n64060 = n45648 & n45899;
  assign n73877 = (n45899 & n63915) | (n45899 & n64060) | (n63915 & n64060);
  assign n73878 = (n45899 & n63914) | (n45899 & n64060) | (n63914 & n64060);
  assign n73879 = (n73748 & n73877) | (n73748 & n73878) | (n73877 & n73878);
  assign n64062 = n45648 | n45899;
  assign n73880 = n63915 | n64062;
  assign n73881 = n63914 | n64062;
  assign n73882 = (n73748 & n73880) | (n73748 & n73881) | (n73880 & n73881);
  assign n45902 = ~n73879 & n73882;
  assign n45903 = x168 & x216;
  assign n45904 = n45902 & n45903;
  assign n45905 = n45902 | n45903;
  assign n45906 = ~n45904 & n45905;
  assign n45907 = n73852 & n45906;
  assign n45908 = n73852 | n45906;
  assign n45909 = ~n45907 & n45908;
  assign n45910 = x167 & x217;
  assign n45911 = n45909 & n45910;
  assign n45912 = n45909 | n45910;
  assign n45913 = ~n45911 & n45912;
  assign n64017 = n45662 | n45664;
  assign n64064 = n45913 & n64017;
  assign n64065 = n45662 & n45913;
  assign n64066 = (n73806 & n64064) | (n73806 & n64065) | (n64064 & n64065);
  assign n64067 = n45913 | n64017;
  assign n64068 = n45662 | n45913;
  assign n64069 = (n73806 & n64067) | (n73806 & n64068) | (n64067 & n64068);
  assign n45916 = ~n64066 & n64069;
  assign n45917 = x166 & x218;
  assign n45918 = n45916 & n45917;
  assign n45919 = n45916 | n45917;
  assign n45920 = ~n45918 & n45919;
  assign n64070 = n45669 & n45920;
  assign n73883 = (n45920 & n63925) | (n45920 & n64070) | (n63925 & n64070);
  assign n73884 = (n45920 & n63924) | (n45920 & n64070) | (n63924 & n64070);
  assign n73885 = (n63719 & n73883) | (n63719 & n73884) | (n73883 & n73884);
  assign n64072 = n45669 | n45920;
  assign n73886 = n63925 | n64072;
  assign n73887 = n63924 | n64072;
  assign n73888 = (n63719 & n73886) | (n63719 & n73887) | (n73886 & n73887);
  assign n45923 = ~n73885 & n73888;
  assign n45924 = x165 & x219;
  assign n45925 = n45923 & n45924;
  assign n45926 = n45923 | n45924;
  assign n45927 = ~n45925 & n45926;
  assign n64015 = n45676 | n45678;
  assign n73889 = n45927 & n64015;
  assign n73846 = n45419 | n45676;
  assign n73847 = (n45676 & n45678) | (n45676 & n73846) | (n45678 & n73846);
  assign n73890 = n45927 & n73847;
  assign n73891 = (n73798 & n73889) | (n73798 & n73890) | (n73889 & n73890);
  assign n73892 = n45927 | n64015;
  assign n73893 = n45927 | n73847;
  assign n73894 = (n73798 & n73892) | (n73798 & n73893) | (n73892 & n73893);
  assign n45930 = ~n73891 & n73894;
  assign n45931 = x164 & x220;
  assign n45932 = n45930 & n45931;
  assign n45933 = n45930 | n45931;
  assign n45934 = ~n45932 & n45933;
  assign n64074 = n45683 & n45934;
  assign n73895 = (n45934 & n63934) | (n45934 & n64074) | (n63934 & n64074);
  assign n73896 = (n45685 & n45934) | (n45685 & n64074) | (n45934 & n64074);
  assign n73897 = (n63791 & n73895) | (n63791 & n73896) | (n73895 & n73896);
  assign n64076 = n45683 | n45934;
  assign n73898 = n63934 | n64076;
  assign n73899 = n45685 | n64076;
  assign n73900 = (n63791 & n73898) | (n63791 & n73899) | (n73898 & n73899);
  assign n45937 = ~n73897 & n73900;
  assign n45938 = x163 & x221;
  assign n45939 = n45937 & n45938;
  assign n45940 = n45937 | n45938;
  assign n45941 = ~n45939 & n45940;
  assign n64078 = n45690 & n45941;
  assign n64079 = (n45941 & n63939) | (n45941 & n64078) | (n63939 & n64078);
  assign n64080 = n45690 | n45941;
  assign n64081 = n63939 | n64080;
  assign n45944 = ~n64079 & n64081;
  assign n45945 = x162 & x222;
  assign n45946 = n45944 & n45945;
  assign n45947 = n45944 | n45945;
  assign n45948 = ~n45946 & n45947;
  assign n64082 = n45697 & n45948;
  assign n64083 = (n45948 & n63943) | (n45948 & n64082) | (n63943 & n64082);
  assign n64084 = n45697 | n45948;
  assign n64085 = n63943 | n64084;
  assign n45951 = ~n64083 & n64085;
  assign n45952 = x161 & x223;
  assign n45953 = n45951 & n45952;
  assign n45954 = n45951 | n45952;
  assign n45955 = ~n45953 & n45954;
  assign n64086 = n45704 & n45955;
  assign n64087 = (n45955 & n63947) | (n45955 & n64086) | (n63947 & n64086);
  assign n64088 = n45704 | n45955;
  assign n64089 = n63947 | n64088;
  assign n45958 = ~n64087 & n64089;
  assign n45959 = x160 & x224;
  assign n45960 = n45958 & n45959;
  assign n45961 = n45958 | n45959;
  assign n45962 = ~n45960 & n45961;
  assign n64090 = n45711 & n45962;
  assign n64091 = (n45962 & n63951) | (n45962 & n64090) | (n63951 & n64090);
  assign n64092 = n45711 | n45962;
  assign n64093 = n63951 | n64092;
  assign n45965 = ~n64091 & n64093;
  assign n45966 = x159 & x225;
  assign n45967 = n45965 & n45966;
  assign n45968 = n45965 | n45966;
  assign n45969 = ~n45967 & n45968;
  assign n64094 = n45718 & n45969;
  assign n64095 = (n45969 & n63955) | (n45969 & n64094) | (n63955 & n64094);
  assign n64096 = n45718 | n45969;
  assign n64097 = n63955 | n64096;
  assign n45972 = ~n64095 & n64097;
  assign n45973 = x158 & x226;
  assign n45974 = n45972 & n45973;
  assign n45975 = n45972 | n45973;
  assign n45976 = ~n45974 & n45975;
  assign n64098 = n45725 & n45976;
  assign n64099 = (n45976 & n63959) | (n45976 & n64098) | (n63959 & n64098);
  assign n64100 = n45725 | n45976;
  assign n64101 = n63959 | n64100;
  assign n45979 = ~n64099 & n64101;
  assign n45980 = x157 & x227;
  assign n45981 = n45979 & n45980;
  assign n45982 = n45979 | n45980;
  assign n45983 = ~n45981 & n45982;
  assign n64102 = n45732 & n45983;
  assign n64103 = (n45983 & n63963) | (n45983 & n64102) | (n63963 & n64102);
  assign n64104 = n45732 | n45983;
  assign n64105 = n63963 | n64104;
  assign n45986 = ~n64103 & n64105;
  assign n45987 = x156 & x228;
  assign n45988 = n45986 & n45987;
  assign n45989 = n45986 | n45987;
  assign n45990 = ~n45988 & n45989;
  assign n64106 = n45739 & n45990;
  assign n64107 = (n45990 & n63967) | (n45990 & n64106) | (n63967 & n64106);
  assign n64108 = n45739 | n45990;
  assign n64109 = n63967 | n64108;
  assign n45993 = ~n64107 & n64109;
  assign n45994 = x155 & x229;
  assign n45995 = n45993 & n45994;
  assign n45996 = n45993 | n45994;
  assign n45997 = ~n45995 & n45996;
  assign n64110 = n45746 & n45997;
  assign n64111 = (n45997 & n63971) | (n45997 & n64110) | (n63971 & n64110);
  assign n64112 = n45746 | n45997;
  assign n64113 = n63971 | n64112;
  assign n46000 = ~n64111 & n64113;
  assign n46001 = x154 & x230;
  assign n46002 = n46000 & n46001;
  assign n46003 = n46000 | n46001;
  assign n46004 = ~n46002 & n46003;
  assign n64114 = n45753 & n46004;
  assign n64115 = (n46004 & n63975) | (n46004 & n64114) | (n63975 & n64114);
  assign n64116 = n45753 | n46004;
  assign n64117 = n63975 | n64116;
  assign n46007 = ~n64115 & n64117;
  assign n46008 = x153 & x231;
  assign n46009 = n46007 & n46008;
  assign n46010 = n46007 | n46008;
  assign n46011 = ~n46009 & n46010;
  assign n64118 = n45760 & n46011;
  assign n64119 = (n46011 & n63979) | (n46011 & n64118) | (n63979 & n64118);
  assign n64120 = n45760 | n46011;
  assign n64121 = n63979 | n64120;
  assign n46014 = ~n64119 & n64121;
  assign n46015 = x152 & x232;
  assign n46016 = n46014 & n46015;
  assign n46017 = n46014 | n46015;
  assign n46018 = ~n46016 & n46017;
  assign n64122 = n45767 & n46018;
  assign n64123 = (n46018 & n63983) | (n46018 & n64122) | (n63983 & n64122);
  assign n64124 = n45767 | n46018;
  assign n64125 = n63983 | n64124;
  assign n46021 = ~n64123 & n64125;
  assign n46022 = x151 & x233;
  assign n46023 = n46021 & n46022;
  assign n46024 = n46021 | n46022;
  assign n46025 = ~n46023 & n46024;
  assign n64126 = n45774 & n46025;
  assign n64127 = (n46025 & n63987) | (n46025 & n64126) | (n63987 & n64126);
  assign n64128 = n45774 | n46025;
  assign n64129 = n63987 | n64128;
  assign n46028 = ~n64127 & n64129;
  assign n46029 = x150 & x234;
  assign n46030 = n46028 & n46029;
  assign n46031 = n46028 | n46029;
  assign n46032 = ~n46030 & n46031;
  assign n64130 = n45781 & n46032;
  assign n64131 = (n46032 & n63991) | (n46032 & n64130) | (n63991 & n64130);
  assign n64132 = n45781 | n46032;
  assign n64133 = n63991 | n64132;
  assign n46035 = ~n64131 & n64133;
  assign n46036 = x149 & x235;
  assign n46037 = n46035 & n46036;
  assign n46038 = n46035 | n46036;
  assign n46039 = ~n46037 & n46038;
  assign n64134 = n45788 & n46039;
  assign n64135 = (n46039 & n63995) | (n46039 & n64134) | (n63995 & n64134);
  assign n64136 = n45788 | n46039;
  assign n64137 = n63995 | n64136;
  assign n46042 = ~n64135 & n64137;
  assign n46043 = x148 & x236;
  assign n46044 = n46042 & n46043;
  assign n46045 = n46042 | n46043;
  assign n46046 = ~n46044 & n46045;
  assign n64138 = n45795 & n46046;
  assign n64139 = (n46046 & n63999) | (n46046 & n64138) | (n63999 & n64138);
  assign n64140 = n45795 | n46046;
  assign n64141 = n63999 | n64140;
  assign n46049 = ~n64139 & n64141;
  assign n46050 = x147 & x237;
  assign n46051 = n46049 & n46050;
  assign n46052 = n46049 | n46050;
  assign n46053 = ~n46051 & n46052;
  assign n64142 = n45802 & n46053;
  assign n64143 = (n46053 & n64003) | (n46053 & n64142) | (n64003 & n64142);
  assign n64144 = n45802 | n46053;
  assign n64145 = n64003 | n64144;
  assign n46056 = ~n64143 & n64145;
  assign n46057 = x146 & x238;
  assign n46058 = n46056 & n46057;
  assign n46059 = n46056 | n46057;
  assign n46060 = ~n46058 & n46059;
  assign n64146 = n45809 & n46060;
  assign n64147 = (n46060 & n64007) | (n46060 & n64146) | (n64007 & n64146);
  assign n64148 = n45809 | n46060;
  assign n64149 = n64007 | n64148;
  assign n46063 = ~n64147 & n64149;
  assign n46064 = x145 & x239;
  assign n46065 = n46063 & n46064;
  assign n46066 = n46063 | n46064;
  assign n46067 = ~n46065 & n46066;
  assign n64150 = n45816 & n46067;
  assign n64151 = (n46067 & n64011) | (n46067 & n64150) | (n64011 & n64150);
  assign n64152 = n45816 | n46067;
  assign n64153 = n64011 | n64152;
  assign n46070 = ~n64151 & n64153;
  assign n64016 = (n73798 & n73847) | (n73798 & n64015) | (n73847 & n64015);
  assign n64157 = n45918 | n45920;
  assign n73901 = n45669 | n45918;
  assign n73902 = (n45918 & n45920) | (n45918 & n73901) | (n45920 & n73901);
  assign n73903 = (n63925 & n64157) | (n63925 & n73902) | (n64157 & n73902);
  assign n73904 = (n63924 & n64157) | (n63924 & n73902) | (n64157 & n73902);
  assign n73905 = (n63719 & n73903) | (n63719 & n73904) | (n73903 & n73904);
  assign n64162 = n45897 | n45899;
  assign n73906 = n45648 | n45897;
  assign n73907 = (n45897 & n45899) | (n45897 & n73906) | (n45899 & n73906);
  assign n73908 = (n63915 & n64162) | (n63915 & n73907) | (n64162 & n73907);
  assign n73909 = (n63914 & n64162) | (n63914 & n73907) | (n64162 & n73907);
  assign n73910 = (n73748 & n73908) | (n73748 & n73909) | (n73908 & n73909);
  assign n46102 = x175 & x210;
  assign n73913 = n45857 | n73869;
  assign n73914 = (n45606 & n73869) | (n45606 & n73913) | (n73869 & n73913);
  assign n64174 = n46102 & n73914;
  assign n73915 = n46102 & n73869;
  assign n73916 = (n45857 & n46102) | (n45857 & n73915) | (n46102 & n73915);
  assign n64176 = (n63896 & n64174) | (n63896 & n73916) | (n64174 & n73916);
  assign n64177 = n46102 | n73914;
  assign n73917 = n46102 | n73869;
  assign n73918 = n45857 | n73917;
  assign n64179 = (n63896 & n64177) | (n63896 & n73918) | (n64177 & n73918);
  assign n46105 = ~n64176 & n64179;
  assign n64181 = n45862 & n46105;
  assign n73919 = (n45864 & n46105) | (n45864 & n64181) | (n46105 & n64181);
  assign n64182 = (n73862 & n73919) | (n73862 & n64181) | (n73919 & n64181);
  assign n64184 = n45862 | n46105;
  assign n73920 = n45864 | n64184;
  assign n64185 = (n73862 & n73920) | (n73862 & n64184) | (n73920 & n64184);
  assign n46108 = ~n64182 & n64185;
  assign n46109 = x174 & x211;
  assign n46110 = n46108 & n46109;
  assign n46111 = n46108 | n46109;
  assign n46112 = ~n46110 & n46111;
  assign n64186 = n45869 & n46112;
  assign n73921 = (n46112 & n64045) | (n46112 & n64186) | (n64045 & n64186);
  assign n73922 = (n46112 & n64044) | (n46112 & n64186) | (n64044 & n64186);
  assign n73923 = (n63884 & n73921) | (n63884 & n73922) | (n73921 & n73922);
  assign n64188 = n45869 | n46112;
  assign n73924 = n64045 | n64188;
  assign n73925 = n64044 | n64188;
  assign n73926 = (n63884 & n73924) | (n63884 & n73925) | (n73924 & n73925);
  assign n46115 = ~n73923 & n73926;
  assign n46116 = x173 & x212;
  assign n46117 = n46115 & n46116;
  assign n46118 = n46115 | n46116;
  assign n46119 = ~n46117 & n46118;
  assign n64167 = n45876 | n45878;
  assign n73927 = n46119 & n64167;
  assign n73911 = n45627 | n45876;
  assign n73912 = (n45876 & n45878) | (n45876 & n73911) | (n45878 & n73911);
  assign n73928 = n46119 & n73912;
  assign n73929 = (n63906 & n73927) | (n63906 & n73928) | (n73927 & n73928);
  assign n73930 = n46119 | n64167;
  assign n73931 = n46119 | n73912;
  assign n73932 = (n63906 & n73930) | (n63906 & n73931) | (n73930 & n73931);
  assign n46122 = ~n73929 & n73932;
  assign n46123 = x172 & x213;
  assign n46124 = n46122 & n46123;
  assign n46125 = n46122 | n46123;
  assign n46126 = ~n46124 & n46125;
  assign n64164 = n45883 | n45885;
  assign n64190 = n46126 & n64164;
  assign n64191 = n45883 & n46126;
  assign n64192 = (n73857 & n64190) | (n73857 & n64191) | (n64190 & n64191);
  assign n64193 = n46126 | n64164;
  assign n64194 = n45883 | n46126;
  assign n64195 = (n73857 & n64193) | (n73857 & n64194) | (n64193 & n64194);
  assign n46129 = ~n64192 & n64195;
  assign n46130 = x171 & x214;
  assign n46131 = n46129 & n46130;
  assign n46132 = n46129 | n46130;
  assign n46133 = ~n46131 & n46132;
  assign n64196 = n45890 & n46133;
  assign n73933 = (n46133 & n64055) | (n46133 & n64196) | (n64055 & n64196);
  assign n73934 = (n46133 & n64054) | (n46133 & n64196) | (n64054 & n64196);
  assign n73935 = (n73811 & n73933) | (n73811 & n73934) | (n73933 & n73934);
  assign n64198 = n45890 | n46133;
  assign n73936 = n64055 | n64198;
  assign n73937 = n64054 | n64198;
  assign n73938 = (n73811 & n73936) | (n73811 & n73937) | (n73936 & n73937);
  assign n46136 = ~n73935 & n73938;
  assign n46137 = x170 & x215;
  assign n46138 = n46136 & n46137;
  assign n46139 = n46136 | n46137;
  assign n46140 = ~n46138 & n46139;
  assign n46141 = n73910 & n46140;
  assign n46142 = n73910 | n46140;
  assign n46143 = ~n46141 & n46142;
  assign n46144 = x169 & x216;
  assign n46145 = n46143 & n46144;
  assign n46146 = n46143 | n46144;
  assign n46147 = ~n46145 & n46146;
  assign n64159 = n45904 | n45906;
  assign n64200 = n46147 & n64159;
  assign n64201 = n45904 & n46147;
  assign n64202 = (n73852 & n64200) | (n73852 & n64201) | (n64200 & n64201);
  assign n64203 = n46147 | n64159;
  assign n64204 = n45904 | n46147;
  assign n64205 = (n73852 & n64203) | (n73852 & n64204) | (n64203 & n64204);
  assign n46150 = ~n64202 & n64205;
  assign n46151 = x168 & x217;
  assign n46152 = n46150 & n46151;
  assign n46153 = n46150 | n46151;
  assign n46154 = ~n46152 & n46153;
  assign n64206 = n45911 & n46154;
  assign n73939 = (n46154 & n64065) | (n46154 & n64206) | (n64065 & n64206);
  assign n73940 = (n46154 & n64064) | (n46154 & n64206) | (n64064 & n64206);
  assign n73941 = (n73806 & n73939) | (n73806 & n73940) | (n73939 & n73940);
  assign n64208 = n45911 | n46154;
  assign n73942 = n64065 | n64208;
  assign n73943 = n64064 | n64208;
  assign n73944 = (n73806 & n73942) | (n73806 & n73943) | (n73942 & n73943);
  assign n46157 = ~n73941 & n73944;
  assign n46158 = x167 & x218;
  assign n46159 = n46157 & n46158;
  assign n46160 = n46157 | n46158;
  assign n46161 = ~n46159 & n46160;
  assign n46162 = n73905 & n46161;
  assign n46163 = n73905 | n46161;
  assign n46164 = ~n46162 & n46163;
  assign n46165 = x166 & x219;
  assign n46166 = n46164 & n46165;
  assign n46167 = n46164 | n46165;
  assign n46168 = ~n46166 & n46167;
  assign n64154 = n45925 | n45927;
  assign n64210 = n46168 & n64154;
  assign n64211 = n45925 & n46168;
  assign n64212 = (n64016 & n64210) | (n64016 & n64211) | (n64210 & n64211);
  assign n64213 = n46168 | n64154;
  assign n64214 = n45925 | n46168;
  assign n64215 = (n64016 & n64213) | (n64016 & n64214) | (n64213 & n64214);
  assign n46171 = ~n64212 & n64215;
  assign n46172 = x165 & x220;
  assign n46173 = n46171 & n46172;
  assign n46174 = n46171 | n46172;
  assign n46175 = ~n46173 & n46174;
  assign n64216 = n45932 & n46175;
  assign n64217 = (n46175 & n73897) | (n46175 & n64216) | (n73897 & n64216);
  assign n64218 = n45932 | n46175;
  assign n64219 = n73897 | n64218;
  assign n46178 = ~n64217 & n64219;
  assign n46179 = x164 & x221;
  assign n46180 = n46178 & n46179;
  assign n46181 = n46178 | n46179;
  assign n46182 = ~n46180 & n46181;
  assign n64220 = n45939 & n46182;
  assign n64221 = (n46182 & n64079) | (n46182 & n64220) | (n64079 & n64220);
  assign n64222 = n45939 | n46182;
  assign n64223 = n64079 | n64222;
  assign n46185 = ~n64221 & n64223;
  assign n46186 = x163 & x222;
  assign n46187 = n46185 & n46186;
  assign n46188 = n46185 | n46186;
  assign n46189 = ~n46187 & n46188;
  assign n64224 = n45946 & n46189;
  assign n64225 = (n46189 & n64083) | (n46189 & n64224) | (n64083 & n64224);
  assign n64226 = n45946 | n46189;
  assign n64227 = n64083 | n64226;
  assign n46192 = ~n64225 & n64227;
  assign n46193 = x162 & x223;
  assign n46194 = n46192 & n46193;
  assign n46195 = n46192 | n46193;
  assign n46196 = ~n46194 & n46195;
  assign n64228 = n45953 & n46196;
  assign n64229 = (n46196 & n64087) | (n46196 & n64228) | (n64087 & n64228);
  assign n64230 = n45953 | n46196;
  assign n64231 = n64087 | n64230;
  assign n46199 = ~n64229 & n64231;
  assign n46200 = x161 & x224;
  assign n46201 = n46199 & n46200;
  assign n46202 = n46199 | n46200;
  assign n46203 = ~n46201 & n46202;
  assign n64232 = n45960 & n46203;
  assign n64233 = (n46203 & n64091) | (n46203 & n64232) | (n64091 & n64232);
  assign n64234 = n45960 | n46203;
  assign n64235 = n64091 | n64234;
  assign n46206 = ~n64233 & n64235;
  assign n46207 = x160 & x225;
  assign n46208 = n46206 & n46207;
  assign n46209 = n46206 | n46207;
  assign n46210 = ~n46208 & n46209;
  assign n64236 = n45967 & n46210;
  assign n64237 = (n46210 & n64095) | (n46210 & n64236) | (n64095 & n64236);
  assign n64238 = n45967 | n46210;
  assign n64239 = n64095 | n64238;
  assign n46213 = ~n64237 & n64239;
  assign n46214 = x159 & x226;
  assign n46215 = n46213 & n46214;
  assign n46216 = n46213 | n46214;
  assign n46217 = ~n46215 & n46216;
  assign n64240 = n45974 & n46217;
  assign n64241 = (n46217 & n64099) | (n46217 & n64240) | (n64099 & n64240);
  assign n64242 = n45974 | n46217;
  assign n64243 = n64099 | n64242;
  assign n46220 = ~n64241 & n64243;
  assign n46221 = x158 & x227;
  assign n46222 = n46220 & n46221;
  assign n46223 = n46220 | n46221;
  assign n46224 = ~n46222 & n46223;
  assign n64244 = n45981 & n46224;
  assign n64245 = (n46224 & n64103) | (n46224 & n64244) | (n64103 & n64244);
  assign n64246 = n45981 | n46224;
  assign n64247 = n64103 | n64246;
  assign n46227 = ~n64245 & n64247;
  assign n46228 = x157 & x228;
  assign n46229 = n46227 & n46228;
  assign n46230 = n46227 | n46228;
  assign n46231 = ~n46229 & n46230;
  assign n64248 = n45988 & n46231;
  assign n64249 = (n46231 & n64107) | (n46231 & n64248) | (n64107 & n64248);
  assign n64250 = n45988 | n46231;
  assign n64251 = n64107 | n64250;
  assign n46234 = ~n64249 & n64251;
  assign n46235 = x156 & x229;
  assign n46236 = n46234 & n46235;
  assign n46237 = n46234 | n46235;
  assign n46238 = ~n46236 & n46237;
  assign n64252 = n45995 & n46238;
  assign n64253 = (n46238 & n64111) | (n46238 & n64252) | (n64111 & n64252);
  assign n64254 = n45995 | n46238;
  assign n64255 = n64111 | n64254;
  assign n46241 = ~n64253 & n64255;
  assign n46242 = x155 & x230;
  assign n46243 = n46241 & n46242;
  assign n46244 = n46241 | n46242;
  assign n46245 = ~n46243 & n46244;
  assign n64256 = n46002 & n46245;
  assign n64257 = (n46245 & n64115) | (n46245 & n64256) | (n64115 & n64256);
  assign n64258 = n46002 | n46245;
  assign n64259 = n64115 | n64258;
  assign n46248 = ~n64257 & n64259;
  assign n46249 = x154 & x231;
  assign n46250 = n46248 & n46249;
  assign n46251 = n46248 | n46249;
  assign n46252 = ~n46250 & n46251;
  assign n64260 = n46009 & n46252;
  assign n64261 = (n46252 & n64119) | (n46252 & n64260) | (n64119 & n64260);
  assign n64262 = n46009 | n46252;
  assign n64263 = n64119 | n64262;
  assign n46255 = ~n64261 & n64263;
  assign n46256 = x153 & x232;
  assign n46257 = n46255 & n46256;
  assign n46258 = n46255 | n46256;
  assign n46259 = ~n46257 & n46258;
  assign n64264 = n46016 & n46259;
  assign n64265 = (n46259 & n64123) | (n46259 & n64264) | (n64123 & n64264);
  assign n64266 = n46016 | n46259;
  assign n64267 = n64123 | n64266;
  assign n46262 = ~n64265 & n64267;
  assign n46263 = x152 & x233;
  assign n46264 = n46262 & n46263;
  assign n46265 = n46262 | n46263;
  assign n46266 = ~n46264 & n46265;
  assign n64268 = n46023 & n46266;
  assign n64269 = (n46266 & n64127) | (n46266 & n64268) | (n64127 & n64268);
  assign n64270 = n46023 | n46266;
  assign n64271 = n64127 | n64270;
  assign n46269 = ~n64269 & n64271;
  assign n46270 = x151 & x234;
  assign n46271 = n46269 & n46270;
  assign n46272 = n46269 | n46270;
  assign n46273 = ~n46271 & n46272;
  assign n64272 = n46030 & n46273;
  assign n64273 = (n46273 & n64131) | (n46273 & n64272) | (n64131 & n64272);
  assign n64274 = n46030 | n46273;
  assign n64275 = n64131 | n64274;
  assign n46276 = ~n64273 & n64275;
  assign n46277 = x150 & x235;
  assign n46278 = n46276 & n46277;
  assign n46279 = n46276 | n46277;
  assign n46280 = ~n46278 & n46279;
  assign n64276 = n46037 & n46280;
  assign n64277 = (n46280 & n64135) | (n46280 & n64276) | (n64135 & n64276);
  assign n64278 = n46037 | n46280;
  assign n64279 = n64135 | n64278;
  assign n46283 = ~n64277 & n64279;
  assign n46284 = x149 & x236;
  assign n46285 = n46283 & n46284;
  assign n46286 = n46283 | n46284;
  assign n46287 = ~n46285 & n46286;
  assign n64280 = n46044 & n46287;
  assign n64281 = (n46287 & n64139) | (n46287 & n64280) | (n64139 & n64280);
  assign n64282 = n46044 | n46287;
  assign n64283 = n64139 | n64282;
  assign n46290 = ~n64281 & n64283;
  assign n46291 = x148 & x237;
  assign n46292 = n46290 & n46291;
  assign n46293 = n46290 | n46291;
  assign n46294 = ~n46292 & n46293;
  assign n64284 = n46051 & n46294;
  assign n64285 = (n46294 & n64143) | (n46294 & n64284) | (n64143 & n64284);
  assign n64286 = n46051 | n46294;
  assign n64287 = n64143 | n64286;
  assign n46297 = ~n64285 & n64287;
  assign n46298 = x147 & x238;
  assign n46299 = n46297 & n46298;
  assign n46300 = n46297 | n46298;
  assign n46301 = ~n46299 & n46300;
  assign n64288 = n46058 & n46301;
  assign n64289 = (n46301 & n64147) | (n46301 & n64288) | (n64147 & n64288);
  assign n64290 = n46058 | n46301;
  assign n64291 = n64147 | n64290;
  assign n46304 = ~n64289 & n64291;
  assign n46305 = x146 & x239;
  assign n46306 = n46304 & n46305;
  assign n46307 = n46304 | n46305;
  assign n46308 = ~n46306 & n46307;
  assign n64292 = n46065 & n46308;
  assign n64293 = (n46308 & n64151) | (n46308 & n64292) | (n64151 & n64292);
  assign n64294 = n46065 | n46308;
  assign n64295 = n64151 | n64294;
  assign n46311 = ~n64293 & n64295;
  assign n64302 = n46152 | n46154;
  assign n73947 = n45911 | n46152;
  assign n73948 = (n46152 & n46154) | (n46152 & n73947) | (n46154 & n73947);
  assign n73949 = (n64065 & n64302) | (n64065 & n73948) | (n64302 & n73948);
  assign n73950 = (n64064 & n64302) | (n64064 & n73948) | (n64302 & n73948);
  assign n73951 = (n73806 & n73949) | (n73806 & n73950) | (n73949 & n73950);
  assign n64307 = n46131 | n46133;
  assign n73952 = n45890 | n46131;
  assign n73953 = (n46131 & n46133) | (n46131 & n73952) | (n46133 & n73952);
  assign n73954 = (n64055 & n64307) | (n64055 & n73953) | (n64307 & n73953);
  assign n73955 = (n64054 & n64307) | (n64054 & n73953) | (n64307 & n73953);
  assign n73956 = (n73811 & n73954) | (n73811 & n73955) | (n73954 & n73955);
  assign n64168 = (n63906 & n73912) | (n63906 & n64167) | (n73912 & n64167);
  assign n64312 = n46110 | n46112;
  assign n73957 = n45869 | n46110;
  assign n73958 = (n46110 & n46112) | (n46110 & n73957) | (n46112 & n73957);
  assign n73959 = (n64045 & n64312) | (n64045 & n73958) | (n64312 & n73958);
  assign n73960 = (n64044 & n64312) | (n64044 & n73958) | (n64312 & n73958);
  assign n73961 = (n63884 & n73959) | (n63884 & n73960) | (n73959 & n73960);
  assign n46342 = x175 & x211;
  assign n73962 = n46342 & n64174;
  assign n73963 = n46342 & n73916;
  assign n73964 = (n63896 & n73962) | (n63896 & n73963) | (n73962 & n73963);
  assign n73965 = (n46342 & n73919) | (n46342 & n73964) | (n73919 & n73964);
  assign n73966 = (n46342 & n64181) | (n46342 & n73964) | (n64181 & n73964);
  assign n73967 = (n73862 & n73965) | (n73862 & n73966) | (n73965 & n73966);
  assign n73968 = n46342 | n64174;
  assign n73969 = n46342 | n73916;
  assign n73970 = (n63896 & n73968) | (n63896 & n73969) | (n73968 & n73969);
  assign n73971 = n73919 | n73970;
  assign n73972 = n64181 | n73970;
  assign n73973 = (n73862 & n73971) | (n73862 & n73972) | (n73971 & n73972);
  assign n46345 = ~n73967 & n73973;
  assign n46346 = n73961 & n46345;
  assign n46347 = n73961 | n46345;
  assign n46348 = ~n46346 & n46347;
  assign n46349 = x174 & x212;
  assign n46350 = n46348 & n46349;
  assign n46351 = n46348 | n46349;
  assign n46352 = ~n46350 & n46351;
  assign n64309 = n46117 | n46119;
  assign n64318 = n46352 & n64309;
  assign n64319 = n46117 & n46352;
  assign n64320 = (n64168 & n64318) | (n64168 & n64319) | (n64318 & n64319);
  assign n64321 = n46352 | n64309;
  assign n64322 = n46117 | n46352;
  assign n64323 = (n64168 & n64321) | (n64168 & n64322) | (n64321 & n64322);
  assign n46355 = ~n64320 & n64323;
  assign n46356 = x173 & x213;
  assign n46357 = n46355 & n46356;
  assign n46358 = n46355 | n46356;
  assign n46359 = ~n46357 & n46358;
  assign n64324 = n46124 & n46359;
  assign n64325 = (n46359 & n64192) | (n46359 & n64324) | (n64192 & n64324);
  assign n64326 = n46124 | n46359;
  assign n64327 = n64192 | n64326;
  assign n46362 = ~n64325 & n64327;
  assign n46363 = x172 & x214;
  assign n46364 = n46362 & n46363;
  assign n46365 = n46362 | n46363;
  assign n46366 = ~n46364 & n46365;
  assign n46367 = n73956 & n46366;
  assign n46368 = n73956 | n46366;
  assign n46369 = ~n46367 & n46368;
  assign n46370 = x171 & x215;
  assign n46371 = n46369 & n46370;
  assign n46372 = n46369 | n46370;
  assign n46373 = ~n46371 & n46372;
  assign n64304 = n46138 | n46140;
  assign n64328 = n46373 & n64304;
  assign n64329 = n46138 & n46373;
  assign n64330 = (n73910 & n64328) | (n73910 & n64329) | (n64328 & n64329);
  assign n64331 = n46373 | n64304;
  assign n64332 = n46138 | n46373;
  assign n64333 = (n73910 & n64331) | (n73910 & n64332) | (n64331 & n64332);
  assign n46376 = ~n64330 & n64333;
  assign n46377 = x170 & x216;
  assign n46378 = n46376 & n46377;
  assign n46379 = n46376 | n46377;
  assign n46380 = ~n46378 & n46379;
  assign n64334 = n46145 & n46380;
  assign n73974 = (n46380 & n64201) | (n46380 & n64334) | (n64201 & n64334);
  assign n73975 = (n46380 & n64200) | (n46380 & n64334) | (n64200 & n64334);
  assign n73976 = (n73852 & n73974) | (n73852 & n73975) | (n73974 & n73975);
  assign n64336 = n46145 | n46380;
  assign n73977 = n64201 | n64336;
  assign n73978 = n64200 | n64336;
  assign n73979 = (n73852 & n73977) | (n73852 & n73978) | (n73977 & n73978);
  assign n46383 = ~n73976 & n73979;
  assign n46384 = x169 & x217;
  assign n46385 = n46383 & n46384;
  assign n46386 = n46383 | n46384;
  assign n46387 = ~n46385 & n46386;
  assign n46388 = n73951 & n46387;
  assign n46389 = n73951 | n46387;
  assign n46390 = ~n46388 & n46389;
  assign n46391 = x168 & x218;
  assign n46392 = n46390 & n46391;
  assign n46393 = n46390 | n46391;
  assign n46394 = ~n46392 & n46393;
  assign n64299 = n46159 | n46161;
  assign n64338 = n46394 & n64299;
  assign n64339 = n46159 & n46394;
  assign n64340 = (n73905 & n64338) | (n73905 & n64339) | (n64338 & n64339);
  assign n64341 = n46394 | n64299;
  assign n64342 = n46159 | n46394;
  assign n64343 = (n73905 & n64341) | (n73905 & n64342) | (n64341 & n64342);
  assign n46397 = ~n64340 & n64343;
  assign n46398 = x167 & x219;
  assign n46399 = n46397 & n46398;
  assign n46400 = n46397 | n46398;
  assign n46401 = ~n46399 & n46400;
  assign n64344 = n46166 & n46401;
  assign n73980 = (n46401 & n64211) | (n46401 & n64344) | (n64211 & n64344);
  assign n73981 = (n46401 & n64210) | (n46401 & n64344) | (n64210 & n64344);
  assign n73982 = (n64016 & n73980) | (n64016 & n73981) | (n73980 & n73981);
  assign n64346 = n46166 | n46401;
  assign n73983 = n64211 | n64346;
  assign n73984 = n64210 | n64346;
  assign n73985 = (n64016 & n73983) | (n64016 & n73984) | (n73983 & n73984);
  assign n46404 = ~n73982 & n73985;
  assign n46405 = x166 & x220;
  assign n46406 = n46404 & n46405;
  assign n46407 = n46404 | n46405;
  assign n46408 = ~n46406 & n46407;
  assign n64297 = n46173 | n46175;
  assign n73986 = n46408 & n64297;
  assign n73945 = n45932 | n46173;
  assign n73946 = (n46173 & n46175) | (n46173 & n73945) | (n46175 & n73945);
  assign n73987 = n46408 & n73946;
  assign n73988 = (n73897 & n73986) | (n73897 & n73987) | (n73986 & n73987);
  assign n73989 = n46408 | n64297;
  assign n73990 = n46408 | n73946;
  assign n73991 = (n73897 & n73989) | (n73897 & n73990) | (n73989 & n73990);
  assign n46411 = ~n73988 & n73991;
  assign n46412 = x165 & x221;
  assign n46413 = n46411 & n46412;
  assign n46414 = n46411 | n46412;
  assign n46415 = ~n46413 & n46414;
  assign n64348 = n46180 & n46415;
  assign n73992 = (n46415 & n64220) | (n46415 & n64348) | (n64220 & n64348);
  assign n73993 = (n46182 & n46415) | (n46182 & n64348) | (n46415 & n64348);
  assign n73994 = (n64079 & n73992) | (n64079 & n73993) | (n73992 & n73993);
  assign n64350 = n46180 | n46415;
  assign n73995 = n64220 | n64350;
  assign n73996 = n46182 | n64350;
  assign n73997 = (n64079 & n73995) | (n64079 & n73996) | (n73995 & n73996);
  assign n46418 = ~n73994 & n73997;
  assign n46419 = x164 & x222;
  assign n46420 = n46418 & n46419;
  assign n46421 = n46418 | n46419;
  assign n46422 = ~n46420 & n46421;
  assign n64352 = n46187 & n46422;
  assign n64353 = (n46422 & n64225) | (n46422 & n64352) | (n64225 & n64352);
  assign n64354 = n46187 | n46422;
  assign n64355 = n64225 | n64354;
  assign n46425 = ~n64353 & n64355;
  assign n46426 = x163 & x223;
  assign n46427 = n46425 & n46426;
  assign n46428 = n46425 | n46426;
  assign n46429 = ~n46427 & n46428;
  assign n64356 = n46194 & n46429;
  assign n64357 = (n46429 & n64229) | (n46429 & n64356) | (n64229 & n64356);
  assign n64358 = n46194 | n46429;
  assign n64359 = n64229 | n64358;
  assign n46432 = ~n64357 & n64359;
  assign n46433 = x162 & x224;
  assign n46434 = n46432 & n46433;
  assign n46435 = n46432 | n46433;
  assign n46436 = ~n46434 & n46435;
  assign n64360 = n46201 & n46436;
  assign n64361 = (n46436 & n64233) | (n46436 & n64360) | (n64233 & n64360);
  assign n64362 = n46201 | n46436;
  assign n64363 = n64233 | n64362;
  assign n46439 = ~n64361 & n64363;
  assign n46440 = x161 & x225;
  assign n46441 = n46439 & n46440;
  assign n46442 = n46439 | n46440;
  assign n46443 = ~n46441 & n46442;
  assign n64364 = n46208 & n46443;
  assign n64365 = (n46443 & n64237) | (n46443 & n64364) | (n64237 & n64364);
  assign n64366 = n46208 | n46443;
  assign n64367 = n64237 | n64366;
  assign n46446 = ~n64365 & n64367;
  assign n46447 = x160 & x226;
  assign n46448 = n46446 & n46447;
  assign n46449 = n46446 | n46447;
  assign n46450 = ~n46448 & n46449;
  assign n64368 = n46215 & n46450;
  assign n64369 = (n46450 & n64241) | (n46450 & n64368) | (n64241 & n64368);
  assign n64370 = n46215 | n46450;
  assign n64371 = n64241 | n64370;
  assign n46453 = ~n64369 & n64371;
  assign n46454 = x159 & x227;
  assign n46455 = n46453 & n46454;
  assign n46456 = n46453 | n46454;
  assign n46457 = ~n46455 & n46456;
  assign n64372 = n46222 & n46457;
  assign n64373 = (n46457 & n64245) | (n46457 & n64372) | (n64245 & n64372);
  assign n64374 = n46222 | n46457;
  assign n64375 = n64245 | n64374;
  assign n46460 = ~n64373 & n64375;
  assign n46461 = x158 & x228;
  assign n46462 = n46460 & n46461;
  assign n46463 = n46460 | n46461;
  assign n46464 = ~n46462 & n46463;
  assign n64376 = n46229 & n46464;
  assign n64377 = (n46464 & n64249) | (n46464 & n64376) | (n64249 & n64376);
  assign n64378 = n46229 | n46464;
  assign n64379 = n64249 | n64378;
  assign n46467 = ~n64377 & n64379;
  assign n46468 = x157 & x229;
  assign n46469 = n46467 & n46468;
  assign n46470 = n46467 | n46468;
  assign n46471 = ~n46469 & n46470;
  assign n64380 = n46236 & n46471;
  assign n64381 = (n46471 & n64253) | (n46471 & n64380) | (n64253 & n64380);
  assign n64382 = n46236 | n46471;
  assign n64383 = n64253 | n64382;
  assign n46474 = ~n64381 & n64383;
  assign n46475 = x156 & x230;
  assign n46476 = n46474 & n46475;
  assign n46477 = n46474 | n46475;
  assign n46478 = ~n46476 & n46477;
  assign n64384 = n46243 & n46478;
  assign n64385 = (n46478 & n64257) | (n46478 & n64384) | (n64257 & n64384);
  assign n64386 = n46243 | n46478;
  assign n64387 = n64257 | n64386;
  assign n46481 = ~n64385 & n64387;
  assign n46482 = x155 & x231;
  assign n46483 = n46481 & n46482;
  assign n46484 = n46481 | n46482;
  assign n46485 = ~n46483 & n46484;
  assign n64388 = n46250 & n46485;
  assign n64389 = (n46485 & n64261) | (n46485 & n64388) | (n64261 & n64388);
  assign n64390 = n46250 | n46485;
  assign n64391 = n64261 | n64390;
  assign n46488 = ~n64389 & n64391;
  assign n46489 = x154 & x232;
  assign n46490 = n46488 & n46489;
  assign n46491 = n46488 | n46489;
  assign n46492 = ~n46490 & n46491;
  assign n64392 = n46257 & n46492;
  assign n64393 = (n46492 & n64265) | (n46492 & n64392) | (n64265 & n64392);
  assign n64394 = n46257 | n46492;
  assign n64395 = n64265 | n64394;
  assign n46495 = ~n64393 & n64395;
  assign n46496 = x153 & x233;
  assign n46497 = n46495 & n46496;
  assign n46498 = n46495 | n46496;
  assign n46499 = ~n46497 & n46498;
  assign n64396 = n46264 & n46499;
  assign n64397 = (n46499 & n64269) | (n46499 & n64396) | (n64269 & n64396);
  assign n64398 = n46264 | n46499;
  assign n64399 = n64269 | n64398;
  assign n46502 = ~n64397 & n64399;
  assign n46503 = x152 & x234;
  assign n46504 = n46502 & n46503;
  assign n46505 = n46502 | n46503;
  assign n46506 = ~n46504 & n46505;
  assign n64400 = n46271 & n46506;
  assign n64401 = (n46506 & n64273) | (n46506 & n64400) | (n64273 & n64400);
  assign n64402 = n46271 | n46506;
  assign n64403 = n64273 | n64402;
  assign n46509 = ~n64401 & n64403;
  assign n46510 = x151 & x235;
  assign n46511 = n46509 & n46510;
  assign n46512 = n46509 | n46510;
  assign n46513 = ~n46511 & n46512;
  assign n64404 = n46278 & n46513;
  assign n64405 = (n46513 & n64277) | (n46513 & n64404) | (n64277 & n64404);
  assign n64406 = n46278 | n46513;
  assign n64407 = n64277 | n64406;
  assign n46516 = ~n64405 & n64407;
  assign n46517 = x150 & x236;
  assign n46518 = n46516 & n46517;
  assign n46519 = n46516 | n46517;
  assign n46520 = ~n46518 & n46519;
  assign n64408 = n46285 & n46520;
  assign n64409 = (n46520 & n64281) | (n46520 & n64408) | (n64281 & n64408);
  assign n64410 = n46285 | n46520;
  assign n64411 = n64281 | n64410;
  assign n46523 = ~n64409 & n64411;
  assign n46524 = x149 & x237;
  assign n46525 = n46523 & n46524;
  assign n46526 = n46523 | n46524;
  assign n46527 = ~n46525 & n46526;
  assign n64412 = n46292 & n46527;
  assign n64413 = (n46527 & n64285) | (n46527 & n64412) | (n64285 & n64412);
  assign n64414 = n46292 | n46527;
  assign n64415 = n64285 | n64414;
  assign n46530 = ~n64413 & n64415;
  assign n46531 = x148 & x238;
  assign n46532 = n46530 & n46531;
  assign n46533 = n46530 | n46531;
  assign n46534 = ~n46532 & n46533;
  assign n64416 = n46299 & n46534;
  assign n64417 = (n46534 & n64289) | (n46534 & n64416) | (n64289 & n64416);
  assign n64418 = n46299 | n46534;
  assign n64419 = n64289 | n64418;
  assign n46537 = ~n64417 & n64419;
  assign n46538 = x147 & x239;
  assign n46539 = n46537 & n46538;
  assign n46540 = n46537 | n46538;
  assign n46541 = ~n46539 & n46540;
  assign n64420 = n46306 & n46541;
  assign n64421 = (n46541 & n64293) | (n46541 & n64420) | (n64293 & n64420);
  assign n64422 = n46306 | n46541;
  assign n64423 = n64293 | n64422;
  assign n46544 = ~n64421 & n64423;
  assign n64298 = (n73897 & n73946) | (n73897 & n64297) | (n73946 & n64297);
  assign n64427 = n46399 | n46401;
  assign n73998 = n46166 | n46399;
  assign n73999 = (n46399 & n46401) | (n46399 & n73998) | (n46401 & n73998);
  assign n74000 = (n64211 & n64427) | (n64211 & n73999) | (n64427 & n73999);
  assign n74001 = (n64210 & n64427) | (n64210 & n73999) | (n64427 & n73999);
  assign n74002 = (n64016 & n74000) | (n64016 & n74001) | (n74000 & n74001);
  assign n64432 = n46378 | n46380;
  assign n74003 = n46145 | n46378;
  assign n74004 = (n46378 & n46380) | (n46378 & n74003) | (n46380 & n74003);
  assign n74005 = (n64201 & n64432) | (n64201 & n74004) | (n64432 & n74004);
  assign n74006 = (n64200 & n64432) | (n64200 & n74004) | (n64432 & n74004);
  assign n74007 = (n73852 & n74005) | (n73852 & n74006) | (n74005 & n74006);
  assign n46574 = x175 & x212;
  assign n74010 = n46574 & n73967;
  assign n74011 = (n46345 & n46574) | (n46345 & n74010) | (n46574 & n74010);
  assign n64442 = n46574 & n73967;
  assign n64443 = (n73961 & n74011) | (n73961 & n64442) | (n74011 & n64442);
  assign n74012 = n46574 | n73967;
  assign n74013 = n46345 | n74012;
  assign n64445 = n46574 | n73967;
  assign n64446 = (n73961 & n74013) | (n73961 & n64445) | (n74013 & n64445);
  assign n46577 = ~n64443 & n64446;
  assign n64447 = n46350 & n46577;
  assign n74014 = (n46577 & n64319) | (n46577 & n64447) | (n64319 & n64447);
  assign n74015 = (n46577 & n64318) | (n46577 & n64447) | (n64318 & n64447);
  assign n74016 = (n64168 & n74014) | (n64168 & n74015) | (n74014 & n74015);
  assign n64449 = n46350 | n46577;
  assign n74017 = n64319 | n64449;
  assign n74018 = n64318 | n64449;
  assign n74019 = (n64168 & n74017) | (n64168 & n74018) | (n74017 & n74018);
  assign n46580 = ~n74016 & n74019;
  assign n46581 = x174 & x213;
  assign n46582 = n46580 & n46581;
  assign n46583 = n46580 | n46581;
  assign n46584 = ~n46582 & n46583;
  assign n64437 = n46357 | n46359;
  assign n74020 = n46584 & n64437;
  assign n74008 = n46124 | n46357;
  assign n74009 = (n46357 & n46359) | (n46357 & n74008) | (n46359 & n74008);
  assign n74021 = n46584 & n74009;
  assign n74022 = (n64192 & n74020) | (n64192 & n74021) | (n74020 & n74021);
  assign n74023 = n46584 | n64437;
  assign n74024 = n46584 | n74009;
  assign n74025 = (n64192 & n74023) | (n64192 & n74024) | (n74023 & n74024);
  assign n46587 = ~n74022 & n74025;
  assign n46588 = x173 & x214;
  assign n46589 = n46587 & n46588;
  assign n46590 = n46587 | n46588;
  assign n46591 = ~n46589 & n46590;
  assign n64434 = n46364 | n46366;
  assign n64451 = n46591 & n64434;
  assign n64452 = n46364 & n46591;
  assign n64453 = (n73956 & n64451) | (n73956 & n64452) | (n64451 & n64452);
  assign n64454 = n46591 | n64434;
  assign n64455 = n46364 | n46591;
  assign n64456 = (n73956 & n64454) | (n73956 & n64455) | (n64454 & n64455);
  assign n46594 = ~n64453 & n64456;
  assign n46595 = x172 & x215;
  assign n46596 = n46594 & n46595;
  assign n46597 = n46594 | n46595;
  assign n46598 = ~n46596 & n46597;
  assign n64457 = n46371 & n46598;
  assign n74026 = (n46598 & n64329) | (n46598 & n64457) | (n64329 & n64457);
  assign n74027 = (n46598 & n64328) | (n46598 & n64457) | (n64328 & n64457);
  assign n74028 = (n73910 & n74026) | (n73910 & n74027) | (n74026 & n74027);
  assign n64459 = n46371 | n46598;
  assign n74029 = n64329 | n64459;
  assign n74030 = n64328 | n64459;
  assign n74031 = (n73910 & n74029) | (n73910 & n74030) | (n74029 & n74030);
  assign n46601 = ~n74028 & n74031;
  assign n46602 = x171 & x216;
  assign n46603 = n46601 & n46602;
  assign n46604 = n46601 | n46602;
  assign n46605 = ~n46603 & n46604;
  assign n46606 = n74007 & n46605;
  assign n46607 = n74007 | n46605;
  assign n46608 = ~n46606 & n46607;
  assign n46609 = x170 & x217;
  assign n46610 = n46608 & n46609;
  assign n46611 = n46608 | n46609;
  assign n46612 = ~n46610 & n46611;
  assign n64429 = n46385 | n46387;
  assign n64461 = n46612 & n64429;
  assign n64462 = n46385 & n46612;
  assign n64463 = (n73951 & n64461) | (n73951 & n64462) | (n64461 & n64462);
  assign n64464 = n46612 | n64429;
  assign n64465 = n46385 | n46612;
  assign n64466 = (n73951 & n64464) | (n73951 & n64465) | (n64464 & n64465);
  assign n46615 = ~n64463 & n64466;
  assign n46616 = x169 & x218;
  assign n46617 = n46615 & n46616;
  assign n46618 = n46615 | n46616;
  assign n46619 = ~n46617 & n46618;
  assign n64467 = n46392 & n46619;
  assign n74032 = (n46619 & n64339) | (n46619 & n64467) | (n64339 & n64467);
  assign n74033 = (n46619 & n64338) | (n46619 & n64467) | (n64338 & n64467);
  assign n74034 = (n73905 & n74032) | (n73905 & n74033) | (n74032 & n74033);
  assign n64469 = n46392 | n46619;
  assign n74035 = n64339 | n64469;
  assign n74036 = n64338 | n64469;
  assign n74037 = (n73905 & n74035) | (n73905 & n74036) | (n74035 & n74036);
  assign n46622 = ~n74034 & n74037;
  assign n46623 = x168 & x219;
  assign n46624 = n46622 & n46623;
  assign n46625 = n46622 | n46623;
  assign n46626 = ~n46624 & n46625;
  assign n46627 = n74002 & n46626;
  assign n46628 = n74002 | n46626;
  assign n46629 = ~n46627 & n46628;
  assign n46630 = x167 & x220;
  assign n46631 = n46629 & n46630;
  assign n46632 = n46629 | n46630;
  assign n46633 = ~n46631 & n46632;
  assign n64424 = n46406 | n46408;
  assign n64471 = n46633 & n64424;
  assign n64472 = n46406 & n46633;
  assign n64473 = (n64298 & n64471) | (n64298 & n64472) | (n64471 & n64472);
  assign n64474 = n46633 | n64424;
  assign n64475 = n46406 | n46633;
  assign n64476 = (n64298 & n64474) | (n64298 & n64475) | (n64474 & n64475);
  assign n46636 = ~n64473 & n64476;
  assign n46637 = x166 & x221;
  assign n46638 = n46636 & n46637;
  assign n46639 = n46636 | n46637;
  assign n46640 = ~n46638 & n46639;
  assign n64477 = n46413 & n46640;
  assign n64478 = (n46640 & n73994) | (n46640 & n64477) | (n73994 & n64477);
  assign n64479 = n46413 | n46640;
  assign n64480 = n73994 | n64479;
  assign n46643 = ~n64478 & n64480;
  assign n46644 = x165 & x222;
  assign n46645 = n46643 & n46644;
  assign n46646 = n46643 | n46644;
  assign n46647 = ~n46645 & n46646;
  assign n64481 = n46420 & n46647;
  assign n64482 = (n46647 & n64353) | (n46647 & n64481) | (n64353 & n64481);
  assign n64483 = n46420 | n46647;
  assign n64484 = n64353 | n64483;
  assign n46650 = ~n64482 & n64484;
  assign n46651 = x164 & x223;
  assign n46652 = n46650 & n46651;
  assign n46653 = n46650 | n46651;
  assign n46654 = ~n46652 & n46653;
  assign n64485 = n46427 & n46654;
  assign n64486 = (n46654 & n64357) | (n46654 & n64485) | (n64357 & n64485);
  assign n64487 = n46427 | n46654;
  assign n64488 = n64357 | n64487;
  assign n46657 = ~n64486 & n64488;
  assign n46658 = x163 & x224;
  assign n46659 = n46657 & n46658;
  assign n46660 = n46657 | n46658;
  assign n46661 = ~n46659 & n46660;
  assign n64489 = n46434 & n46661;
  assign n64490 = (n46661 & n64361) | (n46661 & n64489) | (n64361 & n64489);
  assign n64491 = n46434 | n46661;
  assign n64492 = n64361 | n64491;
  assign n46664 = ~n64490 & n64492;
  assign n46665 = x162 & x225;
  assign n46666 = n46664 & n46665;
  assign n46667 = n46664 | n46665;
  assign n46668 = ~n46666 & n46667;
  assign n64493 = n46441 & n46668;
  assign n64494 = (n46668 & n64365) | (n46668 & n64493) | (n64365 & n64493);
  assign n64495 = n46441 | n46668;
  assign n64496 = n64365 | n64495;
  assign n46671 = ~n64494 & n64496;
  assign n46672 = x161 & x226;
  assign n46673 = n46671 & n46672;
  assign n46674 = n46671 | n46672;
  assign n46675 = ~n46673 & n46674;
  assign n64497 = n46448 & n46675;
  assign n64498 = (n46675 & n64369) | (n46675 & n64497) | (n64369 & n64497);
  assign n64499 = n46448 | n46675;
  assign n64500 = n64369 | n64499;
  assign n46678 = ~n64498 & n64500;
  assign n46679 = x160 & x227;
  assign n46680 = n46678 & n46679;
  assign n46681 = n46678 | n46679;
  assign n46682 = ~n46680 & n46681;
  assign n64501 = n46455 & n46682;
  assign n64502 = (n46682 & n64373) | (n46682 & n64501) | (n64373 & n64501);
  assign n64503 = n46455 | n46682;
  assign n64504 = n64373 | n64503;
  assign n46685 = ~n64502 & n64504;
  assign n46686 = x159 & x228;
  assign n46687 = n46685 & n46686;
  assign n46688 = n46685 | n46686;
  assign n46689 = ~n46687 & n46688;
  assign n64505 = n46462 & n46689;
  assign n64506 = (n46689 & n64377) | (n46689 & n64505) | (n64377 & n64505);
  assign n64507 = n46462 | n46689;
  assign n64508 = n64377 | n64507;
  assign n46692 = ~n64506 & n64508;
  assign n46693 = x158 & x229;
  assign n46694 = n46692 & n46693;
  assign n46695 = n46692 | n46693;
  assign n46696 = ~n46694 & n46695;
  assign n64509 = n46469 & n46696;
  assign n64510 = (n46696 & n64381) | (n46696 & n64509) | (n64381 & n64509);
  assign n64511 = n46469 | n46696;
  assign n64512 = n64381 | n64511;
  assign n46699 = ~n64510 & n64512;
  assign n46700 = x157 & x230;
  assign n46701 = n46699 & n46700;
  assign n46702 = n46699 | n46700;
  assign n46703 = ~n46701 & n46702;
  assign n64513 = n46476 & n46703;
  assign n64514 = (n46703 & n64385) | (n46703 & n64513) | (n64385 & n64513);
  assign n64515 = n46476 | n46703;
  assign n64516 = n64385 | n64515;
  assign n46706 = ~n64514 & n64516;
  assign n46707 = x156 & x231;
  assign n46708 = n46706 & n46707;
  assign n46709 = n46706 | n46707;
  assign n46710 = ~n46708 & n46709;
  assign n64517 = n46483 & n46710;
  assign n64518 = (n46710 & n64389) | (n46710 & n64517) | (n64389 & n64517);
  assign n64519 = n46483 | n46710;
  assign n64520 = n64389 | n64519;
  assign n46713 = ~n64518 & n64520;
  assign n46714 = x155 & x232;
  assign n46715 = n46713 & n46714;
  assign n46716 = n46713 | n46714;
  assign n46717 = ~n46715 & n46716;
  assign n64521 = n46490 & n46717;
  assign n64522 = (n46717 & n64393) | (n46717 & n64521) | (n64393 & n64521);
  assign n64523 = n46490 | n46717;
  assign n64524 = n64393 | n64523;
  assign n46720 = ~n64522 & n64524;
  assign n46721 = x154 & x233;
  assign n46722 = n46720 & n46721;
  assign n46723 = n46720 | n46721;
  assign n46724 = ~n46722 & n46723;
  assign n64525 = n46497 & n46724;
  assign n64526 = (n46724 & n64397) | (n46724 & n64525) | (n64397 & n64525);
  assign n64527 = n46497 | n46724;
  assign n64528 = n64397 | n64527;
  assign n46727 = ~n64526 & n64528;
  assign n46728 = x153 & x234;
  assign n46729 = n46727 & n46728;
  assign n46730 = n46727 | n46728;
  assign n46731 = ~n46729 & n46730;
  assign n64529 = n46504 & n46731;
  assign n64530 = (n46731 & n64401) | (n46731 & n64529) | (n64401 & n64529);
  assign n64531 = n46504 | n46731;
  assign n64532 = n64401 | n64531;
  assign n46734 = ~n64530 & n64532;
  assign n46735 = x152 & x235;
  assign n46736 = n46734 & n46735;
  assign n46737 = n46734 | n46735;
  assign n46738 = ~n46736 & n46737;
  assign n64533 = n46511 & n46738;
  assign n64534 = (n46738 & n64405) | (n46738 & n64533) | (n64405 & n64533);
  assign n64535 = n46511 | n46738;
  assign n64536 = n64405 | n64535;
  assign n46741 = ~n64534 & n64536;
  assign n46742 = x151 & x236;
  assign n46743 = n46741 & n46742;
  assign n46744 = n46741 | n46742;
  assign n46745 = ~n46743 & n46744;
  assign n64537 = n46518 & n46745;
  assign n64538 = (n46745 & n64409) | (n46745 & n64537) | (n64409 & n64537);
  assign n64539 = n46518 | n46745;
  assign n64540 = n64409 | n64539;
  assign n46748 = ~n64538 & n64540;
  assign n46749 = x150 & x237;
  assign n46750 = n46748 & n46749;
  assign n46751 = n46748 | n46749;
  assign n46752 = ~n46750 & n46751;
  assign n64541 = n46525 & n46752;
  assign n64542 = (n46752 & n64413) | (n46752 & n64541) | (n64413 & n64541);
  assign n64543 = n46525 | n46752;
  assign n64544 = n64413 | n64543;
  assign n46755 = ~n64542 & n64544;
  assign n46756 = x149 & x238;
  assign n46757 = n46755 & n46756;
  assign n46758 = n46755 | n46756;
  assign n46759 = ~n46757 & n46758;
  assign n64545 = n46532 & n46759;
  assign n64546 = (n46759 & n64417) | (n46759 & n64545) | (n64417 & n64545);
  assign n64547 = n46532 | n46759;
  assign n64548 = n64417 | n64547;
  assign n46762 = ~n64546 & n64548;
  assign n46763 = x148 & x239;
  assign n46764 = n46762 & n46763;
  assign n46765 = n46762 | n46763;
  assign n46766 = ~n46764 & n46765;
  assign n64549 = n46539 & n46766;
  assign n64550 = (n46766 & n64421) | (n46766 & n64549) | (n64421 & n64549);
  assign n64551 = n46539 | n46766;
  assign n64552 = n64421 | n64551;
  assign n46769 = ~n64550 & n64552;
  assign n64559 = n46617 | n46619;
  assign n74040 = n46392 | n46617;
  assign n74041 = (n46617 & n46619) | (n46617 & n74040) | (n46619 & n74040);
  assign n74042 = (n64339 & n64559) | (n64339 & n74041) | (n64559 & n74041);
  assign n74043 = (n64338 & n64559) | (n64338 & n74041) | (n64559 & n74041);
  assign n74044 = (n73905 & n74042) | (n73905 & n74043) | (n74042 & n74043);
  assign n64564 = n46596 | n46598;
  assign n74045 = n46371 | n46596;
  assign n74046 = (n46596 & n46598) | (n46596 & n74045) | (n46598 & n74045);
  assign n74047 = (n64329 & n64564) | (n64329 & n74046) | (n64564 & n74046);
  assign n74048 = (n64328 & n64564) | (n64328 & n74046) | (n64564 & n74046);
  assign n74049 = (n73910 & n74047) | (n73910 & n74048) | (n74047 & n74048);
  assign n46798 = x175 & x213;
  assign n64569 = n46577 | n64443;
  assign n74050 = (n46350 & n64443) | (n46350 & n64569) | (n64443 & n64569);
  assign n64571 = n46798 & n74050;
  assign n74051 = n46798 & n64443;
  assign n74052 = (n46577 & n46798) | (n46577 & n74051) | (n46798 & n74051);
  assign n74053 = (n64319 & n64571) | (n64319 & n74052) | (n64571 & n74052);
  assign n74054 = (n64318 & n64571) | (n64318 & n74052) | (n64571 & n74052);
  assign n74055 = (n64168 & n74053) | (n64168 & n74054) | (n74053 & n74054);
  assign n64574 = n46798 | n74050;
  assign n74056 = n46798 | n64443;
  assign n74057 = n46577 | n74056;
  assign n74058 = (n64319 & n64574) | (n64319 & n74057) | (n64574 & n74057);
  assign n74059 = (n64318 & n64574) | (n64318 & n74057) | (n64574 & n74057);
  assign n74060 = (n64168 & n74058) | (n64168 & n74059) | (n74058 & n74059);
  assign n46801 = ~n74055 & n74060;
  assign n64578 = n46582 & n46801;
  assign n74061 = (n46584 & n46801) | (n46584 & n64578) | (n46801 & n64578);
  assign n74062 = (n64437 & n64578) | (n64437 & n74061) | (n64578 & n74061);
  assign n74063 = (n64578 & n74009) | (n64578 & n74061) | (n74009 & n74061);
  assign n74064 = (n64192 & n74062) | (n64192 & n74063) | (n74062 & n74063);
  assign n64581 = n46582 | n46801;
  assign n74065 = n46584 | n64581;
  assign n74066 = (n64437 & n64581) | (n64437 & n74065) | (n64581 & n74065);
  assign n74067 = (n64581 & n74009) | (n64581 & n74065) | (n74009 & n74065);
  assign n74068 = (n64192 & n74066) | (n64192 & n74067) | (n74066 & n74067);
  assign n46804 = ~n74064 & n74068;
  assign n46805 = x174 & x214;
  assign n46806 = n46804 & n46805;
  assign n46807 = n46804 | n46805;
  assign n46808 = ~n46806 & n46807;
  assign n64583 = n46589 & n46808;
  assign n64584 = (n46808 & n64453) | (n46808 & n64583) | (n64453 & n64583);
  assign n64585 = n46589 | n46808;
  assign n64586 = n64453 | n64585;
  assign n46811 = ~n64584 & n64586;
  assign n46812 = x173 & x215;
  assign n46813 = n46811 & n46812;
  assign n46814 = n46811 | n46812;
  assign n46815 = ~n46813 & n46814;
  assign n46816 = n74049 & n46815;
  assign n46817 = n74049 | n46815;
  assign n46818 = ~n46816 & n46817;
  assign n46819 = x172 & x216;
  assign n46820 = n46818 & n46819;
  assign n46821 = n46818 | n46819;
  assign n46822 = ~n46820 & n46821;
  assign n64561 = n46603 | n46605;
  assign n64587 = n46822 & n64561;
  assign n64588 = n46603 & n46822;
  assign n64589 = (n74007 & n64587) | (n74007 & n64588) | (n64587 & n64588);
  assign n64590 = n46822 | n64561;
  assign n64591 = n46603 | n46822;
  assign n64592 = (n74007 & n64590) | (n74007 & n64591) | (n64590 & n64591);
  assign n46825 = ~n64589 & n64592;
  assign n46826 = x171 & x217;
  assign n46827 = n46825 & n46826;
  assign n46828 = n46825 | n46826;
  assign n46829 = ~n46827 & n46828;
  assign n64593 = n46610 & n46829;
  assign n74069 = (n46829 & n64462) | (n46829 & n64593) | (n64462 & n64593);
  assign n74070 = (n46829 & n64461) | (n46829 & n64593) | (n64461 & n64593);
  assign n74071 = (n73951 & n74069) | (n73951 & n74070) | (n74069 & n74070);
  assign n64595 = n46610 | n46829;
  assign n74072 = n64462 | n64595;
  assign n74073 = n64461 | n64595;
  assign n74074 = (n73951 & n74072) | (n73951 & n74073) | (n74072 & n74073);
  assign n46832 = ~n74071 & n74074;
  assign n46833 = x170 & x218;
  assign n46834 = n46832 & n46833;
  assign n46835 = n46832 | n46833;
  assign n46836 = ~n46834 & n46835;
  assign n46837 = n74044 & n46836;
  assign n46838 = n74044 | n46836;
  assign n46839 = ~n46837 & n46838;
  assign n46840 = x169 & x219;
  assign n46841 = n46839 & n46840;
  assign n46842 = n46839 | n46840;
  assign n46843 = ~n46841 & n46842;
  assign n64556 = n46624 | n46626;
  assign n64597 = n46843 & n64556;
  assign n64598 = n46624 & n46843;
  assign n64599 = (n74002 & n64597) | (n74002 & n64598) | (n64597 & n64598);
  assign n64600 = n46843 | n64556;
  assign n64601 = n46624 | n46843;
  assign n64602 = (n74002 & n64600) | (n74002 & n64601) | (n64600 & n64601);
  assign n46846 = ~n64599 & n64602;
  assign n46847 = x168 & x220;
  assign n46848 = n46846 & n46847;
  assign n46849 = n46846 | n46847;
  assign n46850 = ~n46848 & n46849;
  assign n64603 = n46631 & n46850;
  assign n74075 = (n46850 & n64472) | (n46850 & n64603) | (n64472 & n64603);
  assign n74076 = (n46850 & n64471) | (n46850 & n64603) | (n64471 & n64603);
  assign n74077 = (n64298 & n74075) | (n64298 & n74076) | (n74075 & n74076);
  assign n64605 = n46631 | n46850;
  assign n74078 = n64472 | n64605;
  assign n74079 = n64471 | n64605;
  assign n74080 = (n64298 & n74078) | (n64298 & n74079) | (n74078 & n74079);
  assign n46853 = ~n74077 & n74080;
  assign n46854 = x167 & x221;
  assign n46855 = n46853 & n46854;
  assign n46856 = n46853 | n46854;
  assign n46857 = ~n46855 & n46856;
  assign n64554 = n46638 | n46640;
  assign n74081 = n46857 & n64554;
  assign n74038 = n46413 | n46638;
  assign n74039 = (n46638 & n46640) | (n46638 & n74038) | (n46640 & n74038);
  assign n74082 = n46857 & n74039;
  assign n74083 = (n73994 & n74081) | (n73994 & n74082) | (n74081 & n74082);
  assign n74084 = n46857 | n64554;
  assign n74085 = n46857 | n74039;
  assign n74086 = (n73994 & n74084) | (n73994 & n74085) | (n74084 & n74085);
  assign n46860 = ~n74083 & n74086;
  assign n46861 = x166 & x222;
  assign n46862 = n46860 & n46861;
  assign n46863 = n46860 | n46861;
  assign n46864 = ~n46862 & n46863;
  assign n64607 = n46645 & n46864;
  assign n74087 = (n46864 & n64481) | (n46864 & n64607) | (n64481 & n64607);
  assign n74088 = (n46647 & n46864) | (n46647 & n64607) | (n46864 & n64607);
  assign n74089 = (n64353 & n74087) | (n64353 & n74088) | (n74087 & n74088);
  assign n64609 = n46645 | n46864;
  assign n74090 = n64481 | n64609;
  assign n74091 = n46647 | n64609;
  assign n74092 = (n64353 & n74090) | (n64353 & n74091) | (n74090 & n74091);
  assign n46867 = ~n74089 & n74092;
  assign n46868 = x165 & x223;
  assign n46869 = n46867 & n46868;
  assign n46870 = n46867 | n46868;
  assign n46871 = ~n46869 & n46870;
  assign n64611 = n46652 & n46871;
  assign n64612 = (n46871 & n64486) | (n46871 & n64611) | (n64486 & n64611);
  assign n64613 = n46652 | n46871;
  assign n64614 = n64486 | n64613;
  assign n46874 = ~n64612 & n64614;
  assign n46875 = x164 & x224;
  assign n46876 = n46874 & n46875;
  assign n46877 = n46874 | n46875;
  assign n46878 = ~n46876 & n46877;
  assign n64615 = n46659 & n46878;
  assign n64616 = (n46878 & n64490) | (n46878 & n64615) | (n64490 & n64615);
  assign n64617 = n46659 | n46878;
  assign n64618 = n64490 | n64617;
  assign n46881 = ~n64616 & n64618;
  assign n46882 = x163 & x225;
  assign n46883 = n46881 & n46882;
  assign n46884 = n46881 | n46882;
  assign n46885 = ~n46883 & n46884;
  assign n64619 = n46666 & n46885;
  assign n64620 = (n46885 & n64494) | (n46885 & n64619) | (n64494 & n64619);
  assign n64621 = n46666 | n46885;
  assign n64622 = n64494 | n64621;
  assign n46888 = ~n64620 & n64622;
  assign n46889 = x162 & x226;
  assign n46890 = n46888 & n46889;
  assign n46891 = n46888 | n46889;
  assign n46892 = ~n46890 & n46891;
  assign n64623 = n46673 & n46892;
  assign n64624 = (n46892 & n64498) | (n46892 & n64623) | (n64498 & n64623);
  assign n64625 = n46673 | n46892;
  assign n64626 = n64498 | n64625;
  assign n46895 = ~n64624 & n64626;
  assign n46896 = x161 & x227;
  assign n46897 = n46895 & n46896;
  assign n46898 = n46895 | n46896;
  assign n46899 = ~n46897 & n46898;
  assign n64627 = n46680 & n46899;
  assign n64628 = (n46899 & n64502) | (n46899 & n64627) | (n64502 & n64627);
  assign n64629 = n46680 | n46899;
  assign n64630 = n64502 | n64629;
  assign n46902 = ~n64628 & n64630;
  assign n46903 = x160 & x228;
  assign n46904 = n46902 & n46903;
  assign n46905 = n46902 | n46903;
  assign n46906 = ~n46904 & n46905;
  assign n64631 = n46687 & n46906;
  assign n64632 = (n46906 & n64506) | (n46906 & n64631) | (n64506 & n64631);
  assign n64633 = n46687 | n46906;
  assign n64634 = n64506 | n64633;
  assign n46909 = ~n64632 & n64634;
  assign n46910 = x159 & x229;
  assign n46911 = n46909 & n46910;
  assign n46912 = n46909 | n46910;
  assign n46913 = ~n46911 & n46912;
  assign n64635 = n46694 & n46913;
  assign n64636 = (n46913 & n64510) | (n46913 & n64635) | (n64510 & n64635);
  assign n64637 = n46694 | n46913;
  assign n64638 = n64510 | n64637;
  assign n46916 = ~n64636 & n64638;
  assign n46917 = x158 & x230;
  assign n46918 = n46916 & n46917;
  assign n46919 = n46916 | n46917;
  assign n46920 = ~n46918 & n46919;
  assign n64639 = n46701 & n46920;
  assign n64640 = (n46920 & n64514) | (n46920 & n64639) | (n64514 & n64639);
  assign n64641 = n46701 | n46920;
  assign n64642 = n64514 | n64641;
  assign n46923 = ~n64640 & n64642;
  assign n46924 = x157 & x231;
  assign n46925 = n46923 & n46924;
  assign n46926 = n46923 | n46924;
  assign n46927 = ~n46925 & n46926;
  assign n64643 = n46708 & n46927;
  assign n64644 = (n46927 & n64518) | (n46927 & n64643) | (n64518 & n64643);
  assign n64645 = n46708 | n46927;
  assign n64646 = n64518 | n64645;
  assign n46930 = ~n64644 & n64646;
  assign n46931 = x156 & x232;
  assign n46932 = n46930 & n46931;
  assign n46933 = n46930 | n46931;
  assign n46934 = ~n46932 & n46933;
  assign n64647 = n46715 & n46934;
  assign n64648 = (n46934 & n64522) | (n46934 & n64647) | (n64522 & n64647);
  assign n64649 = n46715 | n46934;
  assign n64650 = n64522 | n64649;
  assign n46937 = ~n64648 & n64650;
  assign n46938 = x155 & x233;
  assign n46939 = n46937 & n46938;
  assign n46940 = n46937 | n46938;
  assign n46941 = ~n46939 & n46940;
  assign n64651 = n46722 & n46941;
  assign n64652 = (n46941 & n64526) | (n46941 & n64651) | (n64526 & n64651);
  assign n64653 = n46722 | n46941;
  assign n64654 = n64526 | n64653;
  assign n46944 = ~n64652 & n64654;
  assign n46945 = x154 & x234;
  assign n46946 = n46944 & n46945;
  assign n46947 = n46944 | n46945;
  assign n46948 = ~n46946 & n46947;
  assign n64655 = n46729 & n46948;
  assign n64656 = (n46948 & n64530) | (n46948 & n64655) | (n64530 & n64655);
  assign n64657 = n46729 | n46948;
  assign n64658 = n64530 | n64657;
  assign n46951 = ~n64656 & n64658;
  assign n46952 = x153 & x235;
  assign n46953 = n46951 & n46952;
  assign n46954 = n46951 | n46952;
  assign n46955 = ~n46953 & n46954;
  assign n64659 = n46736 & n46955;
  assign n64660 = (n46955 & n64534) | (n46955 & n64659) | (n64534 & n64659);
  assign n64661 = n46736 | n46955;
  assign n64662 = n64534 | n64661;
  assign n46958 = ~n64660 & n64662;
  assign n46959 = x152 & x236;
  assign n46960 = n46958 & n46959;
  assign n46961 = n46958 | n46959;
  assign n46962 = ~n46960 & n46961;
  assign n64663 = n46743 & n46962;
  assign n64664 = (n46962 & n64538) | (n46962 & n64663) | (n64538 & n64663);
  assign n64665 = n46743 | n46962;
  assign n64666 = n64538 | n64665;
  assign n46965 = ~n64664 & n64666;
  assign n46966 = x151 & x237;
  assign n46967 = n46965 & n46966;
  assign n46968 = n46965 | n46966;
  assign n46969 = ~n46967 & n46968;
  assign n64667 = n46750 & n46969;
  assign n64668 = (n46969 & n64542) | (n46969 & n64667) | (n64542 & n64667);
  assign n64669 = n46750 | n46969;
  assign n64670 = n64542 | n64669;
  assign n46972 = ~n64668 & n64670;
  assign n46973 = x150 & x238;
  assign n46974 = n46972 & n46973;
  assign n46975 = n46972 | n46973;
  assign n46976 = ~n46974 & n46975;
  assign n64671 = n46757 & n46976;
  assign n64672 = (n46976 & n64546) | (n46976 & n64671) | (n64546 & n64671);
  assign n64673 = n46757 | n46976;
  assign n64674 = n64546 | n64673;
  assign n46979 = ~n64672 & n64674;
  assign n46980 = x149 & x239;
  assign n46981 = n46979 & n46980;
  assign n46982 = n46979 | n46980;
  assign n46983 = ~n46981 & n46982;
  assign n64675 = n46764 & n46983;
  assign n64676 = (n46983 & n64550) | (n46983 & n64675) | (n64550 & n64675);
  assign n64677 = n46764 | n46983;
  assign n64678 = n64550 | n64677;
  assign n46986 = ~n64676 & n64678;
  assign n64555 = (n73994 & n74039) | (n73994 & n64554) | (n74039 & n64554);
  assign n64682 = n46848 | n46850;
  assign n74093 = n46631 | n46848;
  assign n74094 = (n46848 & n46850) | (n46848 & n74093) | (n46850 & n74093);
  assign n74095 = (n64472 & n64682) | (n64472 & n74094) | (n64682 & n74094);
  assign n74096 = (n64471 & n64682) | (n64471 & n74094) | (n64682 & n74094);
  assign n74097 = (n64298 & n74095) | (n64298 & n74096) | (n74095 & n74096);
  assign n64687 = n46827 | n46829;
  assign n74098 = n46610 | n46827;
  assign n74099 = (n46827 & n46829) | (n46827 & n74098) | (n46829 & n74098);
  assign n74100 = (n64462 & n64687) | (n64462 & n74099) | (n64687 & n74099);
  assign n74101 = (n64461 & n64687) | (n64461 & n74099) | (n64687 & n74099);
  assign n74102 = (n73951 & n74100) | (n73951 & n74101) | (n74100 & n74101);
  assign n47014 = x175 & x214;
  assign n64694 = n47014 & n74055;
  assign n64695 = (n47014 & n74064) | (n47014 & n64694) | (n74064 & n64694);
  assign n64696 = n47014 | n74055;
  assign n64697 = n74064 | n64696;
  assign n47017 = ~n64695 & n64697;
  assign n64692 = n46806 | n46808;
  assign n74105 = n47017 & n64692;
  assign n74103 = n46589 | n46806;
  assign n74104 = (n46806 & n46808) | (n46806 & n74103) | (n46808 & n74103);
  assign n74106 = n47017 & n74104;
  assign n74107 = (n64453 & n74105) | (n64453 & n74106) | (n74105 & n74106);
  assign n74108 = n47017 | n64692;
  assign n74109 = n47017 | n74104;
  assign n74110 = (n64453 & n74108) | (n64453 & n74109) | (n74108 & n74109);
  assign n47020 = ~n74107 & n74110;
  assign n47021 = x174 & x215;
  assign n47022 = n47020 & n47021;
  assign n47023 = n47020 | n47021;
  assign n47024 = ~n47022 & n47023;
  assign n64689 = n46813 | n46815;
  assign n64698 = n47024 & n64689;
  assign n64699 = n46813 & n47024;
  assign n64700 = (n74049 & n64698) | (n74049 & n64699) | (n64698 & n64699);
  assign n64701 = n47024 | n64689;
  assign n64702 = n46813 | n47024;
  assign n64703 = (n74049 & n64701) | (n74049 & n64702) | (n64701 & n64702);
  assign n47027 = ~n64700 & n64703;
  assign n47028 = x173 & x216;
  assign n47029 = n47027 & n47028;
  assign n47030 = n47027 | n47028;
  assign n47031 = ~n47029 & n47030;
  assign n64704 = n46820 & n47031;
  assign n74111 = (n47031 & n64588) | (n47031 & n64704) | (n64588 & n64704);
  assign n74112 = (n47031 & n64587) | (n47031 & n64704) | (n64587 & n64704);
  assign n74113 = (n74007 & n74111) | (n74007 & n74112) | (n74111 & n74112);
  assign n64706 = n46820 | n47031;
  assign n74114 = n64588 | n64706;
  assign n74115 = n64587 | n64706;
  assign n74116 = (n74007 & n74114) | (n74007 & n74115) | (n74114 & n74115);
  assign n47034 = ~n74113 & n74116;
  assign n47035 = x172 & x217;
  assign n47036 = n47034 & n47035;
  assign n47037 = n47034 | n47035;
  assign n47038 = ~n47036 & n47037;
  assign n47039 = n74102 & n47038;
  assign n47040 = n74102 | n47038;
  assign n47041 = ~n47039 & n47040;
  assign n47042 = x171 & x218;
  assign n47043 = n47041 & n47042;
  assign n47044 = n47041 | n47042;
  assign n47045 = ~n47043 & n47044;
  assign n64684 = n46834 | n46836;
  assign n64708 = n47045 & n64684;
  assign n64709 = n46834 & n47045;
  assign n64710 = (n74044 & n64708) | (n74044 & n64709) | (n64708 & n64709);
  assign n64711 = n47045 | n64684;
  assign n64712 = n46834 | n47045;
  assign n64713 = (n74044 & n64711) | (n74044 & n64712) | (n64711 & n64712);
  assign n47048 = ~n64710 & n64713;
  assign n47049 = x170 & x219;
  assign n47050 = n47048 & n47049;
  assign n47051 = n47048 | n47049;
  assign n47052 = ~n47050 & n47051;
  assign n64714 = n46841 & n47052;
  assign n74117 = (n47052 & n64598) | (n47052 & n64714) | (n64598 & n64714);
  assign n74118 = (n47052 & n64597) | (n47052 & n64714) | (n64597 & n64714);
  assign n74119 = (n74002 & n74117) | (n74002 & n74118) | (n74117 & n74118);
  assign n64716 = n46841 | n47052;
  assign n74120 = n64598 | n64716;
  assign n74121 = n64597 | n64716;
  assign n74122 = (n74002 & n74120) | (n74002 & n74121) | (n74120 & n74121);
  assign n47055 = ~n74119 & n74122;
  assign n47056 = x169 & x220;
  assign n47057 = n47055 & n47056;
  assign n47058 = n47055 | n47056;
  assign n47059 = ~n47057 & n47058;
  assign n47060 = n74097 & n47059;
  assign n47061 = n74097 | n47059;
  assign n47062 = ~n47060 & n47061;
  assign n47063 = x168 & x221;
  assign n47064 = n47062 & n47063;
  assign n47065 = n47062 | n47063;
  assign n47066 = ~n47064 & n47065;
  assign n64679 = n46855 | n46857;
  assign n64718 = n47066 & n64679;
  assign n64719 = n46855 & n47066;
  assign n64720 = (n64555 & n64718) | (n64555 & n64719) | (n64718 & n64719);
  assign n64721 = n47066 | n64679;
  assign n64722 = n46855 | n47066;
  assign n64723 = (n64555 & n64721) | (n64555 & n64722) | (n64721 & n64722);
  assign n47069 = ~n64720 & n64723;
  assign n47070 = x167 & x222;
  assign n47071 = n47069 & n47070;
  assign n47072 = n47069 | n47070;
  assign n47073 = ~n47071 & n47072;
  assign n64724 = n46862 & n47073;
  assign n64725 = (n47073 & n74089) | (n47073 & n64724) | (n74089 & n64724);
  assign n64726 = n46862 | n47073;
  assign n64727 = n74089 | n64726;
  assign n47076 = ~n64725 & n64727;
  assign n47077 = x166 & x223;
  assign n47078 = n47076 & n47077;
  assign n47079 = n47076 | n47077;
  assign n47080 = ~n47078 & n47079;
  assign n64728 = n46869 & n47080;
  assign n64729 = (n47080 & n64612) | (n47080 & n64728) | (n64612 & n64728);
  assign n64730 = n46869 | n47080;
  assign n64731 = n64612 | n64730;
  assign n47083 = ~n64729 & n64731;
  assign n47084 = x165 & x224;
  assign n47085 = n47083 & n47084;
  assign n47086 = n47083 | n47084;
  assign n47087 = ~n47085 & n47086;
  assign n64732 = n46876 & n47087;
  assign n64733 = (n47087 & n64616) | (n47087 & n64732) | (n64616 & n64732);
  assign n64734 = n46876 | n47087;
  assign n64735 = n64616 | n64734;
  assign n47090 = ~n64733 & n64735;
  assign n47091 = x164 & x225;
  assign n47092 = n47090 & n47091;
  assign n47093 = n47090 | n47091;
  assign n47094 = ~n47092 & n47093;
  assign n64736 = n46883 & n47094;
  assign n64737 = (n47094 & n64620) | (n47094 & n64736) | (n64620 & n64736);
  assign n64738 = n46883 | n47094;
  assign n64739 = n64620 | n64738;
  assign n47097 = ~n64737 & n64739;
  assign n47098 = x163 & x226;
  assign n47099 = n47097 & n47098;
  assign n47100 = n47097 | n47098;
  assign n47101 = ~n47099 & n47100;
  assign n64740 = n46890 & n47101;
  assign n64741 = (n47101 & n64624) | (n47101 & n64740) | (n64624 & n64740);
  assign n64742 = n46890 | n47101;
  assign n64743 = n64624 | n64742;
  assign n47104 = ~n64741 & n64743;
  assign n47105 = x162 & x227;
  assign n47106 = n47104 & n47105;
  assign n47107 = n47104 | n47105;
  assign n47108 = ~n47106 & n47107;
  assign n64744 = n46897 & n47108;
  assign n64745 = (n47108 & n64628) | (n47108 & n64744) | (n64628 & n64744);
  assign n64746 = n46897 | n47108;
  assign n64747 = n64628 | n64746;
  assign n47111 = ~n64745 & n64747;
  assign n47112 = x161 & x228;
  assign n47113 = n47111 & n47112;
  assign n47114 = n47111 | n47112;
  assign n47115 = ~n47113 & n47114;
  assign n64748 = n46904 & n47115;
  assign n64749 = (n47115 & n64632) | (n47115 & n64748) | (n64632 & n64748);
  assign n64750 = n46904 | n47115;
  assign n64751 = n64632 | n64750;
  assign n47118 = ~n64749 & n64751;
  assign n47119 = x160 & x229;
  assign n47120 = n47118 & n47119;
  assign n47121 = n47118 | n47119;
  assign n47122 = ~n47120 & n47121;
  assign n64752 = n46911 & n47122;
  assign n64753 = (n47122 & n64636) | (n47122 & n64752) | (n64636 & n64752);
  assign n64754 = n46911 | n47122;
  assign n64755 = n64636 | n64754;
  assign n47125 = ~n64753 & n64755;
  assign n47126 = x159 & x230;
  assign n47127 = n47125 & n47126;
  assign n47128 = n47125 | n47126;
  assign n47129 = ~n47127 & n47128;
  assign n64756 = n46918 & n47129;
  assign n64757 = (n47129 & n64640) | (n47129 & n64756) | (n64640 & n64756);
  assign n64758 = n46918 | n47129;
  assign n64759 = n64640 | n64758;
  assign n47132 = ~n64757 & n64759;
  assign n47133 = x158 & x231;
  assign n47134 = n47132 & n47133;
  assign n47135 = n47132 | n47133;
  assign n47136 = ~n47134 & n47135;
  assign n64760 = n46925 & n47136;
  assign n64761 = (n47136 & n64644) | (n47136 & n64760) | (n64644 & n64760);
  assign n64762 = n46925 | n47136;
  assign n64763 = n64644 | n64762;
  assign n47139 = ~n64761 & n64763;
  assign n47140 = x157 & x232;
  assign n47141 = n47139 & n47140;
  assign n47142 = n47139 | n47140;
  assign n47143 = ~n47141 & n47142;
  assign n64764 = n46932 & n47143;
  assign n64765 = (n47143 & n64648) | (n47143 & n64764) | (n64648 & n64764);
  assign n64766 = n46932 | n47143;
  assign n64767 = n64648 | n64766;
  assign n47146 = ~n64765 & n64767;
  assign n47147 = x156 & x233;
  assign n47148 = n47146 & n47147;
  assign n47149 = n47146 | n47147;
  assign n47150 = ~n47148 & n47149;
  assign n64768 = n46939 & n47150;
  assign n64769 = (n47150 & n64652) | (n47150 & n64768) | (n64652 & n64768);
  assign n64770 = n46939 | n47150;
  assign n64771 = n64652 | n64770;
  assign n47153 = ~n64769 & n64771;
  assign n47154 = x155 & x234;
  assign n47155 = n47153 & n47154;
  assign n47156 = n47153 | n47154;
  assign n47157 = ~n47155 & n47156;
  assign n64772 = n46946 & n47157;
  assign n64773 = (n47157 & n64656) | (n47157 & n64772) | (n64656 & n64772);
  assign n64774 = n46946 | n47157;
  assign n64775 = n64656 | n64774;
  assign n47160 = ~n64773 & n64775;
  assign n47161 = x154 & x235;
  assign n47162 = n47160 & n47161;
  assign n47163 = n47160 | n47161;
  assign n47164 = ~n47162 & n47163;
  assign n64776 = n46953 & n47164;
  assign n64777 = (n47164 & n64660) | (n47164 & n64776) | (n64660 & n64776);
  assign n64778 = n46953 | n47164;
  assign n64779 = n64660 | n64778;
  assign n47167 = ~n64777 & n64779;
  assign n47168 = x153 & x236;
  assign n47169 = n47167 & n47168;
  assign n47170 = n47167 | n47168;
  assign n47171 = ~n47169 & n47170;
  assign n64780 = n46960 & n47171;
  assign n64781 = (n47171 & n64664) | (n47171 & n64780) | (n64664 & n64780);
  assign n64782 = n46960 | n47171;
  assign n64783 = n64664 | n64782;
  assign n47174 = ~n64781 & n64783;
  assign n47175 = x152 & x237;
  assign n47176 = n47174 & n47175;
  assign n47177 = n47174 | n47175;
  assign n47178 = ~n47176 & n47177;
  assign n64784 = n46967 & n47178;
  assign n64785 = (n47178 & n64668) | (n47178 & n64784) | (n64668 & n64784);
  assign n64786 = n46967 | n47178;
  assign n64787 = n64668 | n64786;
  assign n47181 = ~n64785 & n64787;
  assign n47182 = x151 & x238;
  assign n47183 = n47181 & n47182;
  assign n47184 = n47181 | n47182;
  assign n47185 = ~n47183 & n47184;
  assign n64788 = n46974 & n47185;
  assign n64789 = (n47185 & n64672) | (n47185 & n64788) | (n64672 & n64788);
  assign n64790 = n46974 | n47185;
  assign n64791 = n64672 | n64790;
  assign n47188 = ~n64789 & n64791;
  assign n47189 = x150 & x239;
  assign n47190 = n47188 & n47189;
  assign n47191 = n47188 | n47189;
  assign n47192 = ~n47190 & n47191;
  assign n64792 = n46981 & n47192;
  assign n64793 = (n47192 & n64676) | (n47192 & n64792) | (n64676 & n64792);
  assign n64794 = n46981 | n47192;
  assign n64795 = n64676 | n64794;
  assign n47195 = ~n64793 & n64795;
  assign n64802 = n47050 | n47052;
  assign n74125 = n46841 | n47050;
  assign n74126 = (n47050 & n47052) | (n47050 & n74125) | (n47052 & n74125);
  assign n74127 = (n64598 & n64802) | (n64598 & n74126) | (n64802 & n74126);
  assign n74128 = (n64597 & n64802) | (n64597 & n74126) | (n64802 & n74126);
  assign n74129 = (n74002 & n74127) | (n74002 & n74128) | (n74127 & n74128);
  assign n64807 = n47029 | n47031;
  assign n74130 = n46820 | n47029;
  assign n74131 = (n47029 & n47031) | (n47029 & n74130) | (n47031 & n74130);
  assign n74132 = (n64588 & n64807) | (n64588 & n74131) | (n64807 & n74131);
  assign n74133 = (n64587 & n64807) | (n64587 & n74131) | (n64807 & n74131);
  assign n74134 = (n74007 & n74132) | (n74007 & n74133) | (n74132 & n74133);
  assign n47222 = x175 & x215;
  assign n74136 = n47222 & n64694;
  assign n74137 = n47014 & n47222;
  assign n74138 = (n74064 & n74136) | (n74064 & n74137) | (n74136 & n74137);
  assign n74135 = (n47017 & n47222) | (n47017 & n74138) | (n47222 & n74138);
  assign n74139 = (n64692 & n74135) | (n64692 & n74138) | (n74135 & n74138);
  assign n74140 = (n74104 & n74135) | (n74104 & n74138) | (n74135 & n74138);
  assign n74141 = (n64453 & n74139) | (n64453 & n74140) | (n74139 & n74140);
  assign n74143 = n47222 | n64694;
  assign n74144 = n47014 | n47222;
  assign n74145 = (n74064 & n74143) | (n74064 & n74144) | (n74143 & n74144);
  assign n74142 = n47017 | n74145;
  assign n74146 = (n64692 & n74142) | (n64692 & n74145) | (n74142 & n74145);
  assign n74147 = (n74104 & n74142) | (n74104 & n74145) | (n74142 & n74145);
  assign n74148 = (n64453 & n74146) | (n64453 & n74147) | (n74146 & n74147);
  assign n47225 = ~n74141 & n74148;
  assign n64817 = n47022 & n47225;
  assign n64818 = (n47225 & n64700) | (n47225 & n64817) | (n64700 & n64817);
  assign n64819 = n47022 | n47225;
  assign n64820 = n64700 | n64819;
  assign n47228 = ~n64818 & n64820;
  assign n47229 = x174 & x216;
  assign n47230 = n47228 & n47229;
  assign n47231 = n47228 | n47229;
  assign n47232 = ~n47230 & n47231;
  assign n47233 = n74134 & n47232;
  assign n47234 = n74134 | n47232;
  assign n47235 = ~n47233 & n47234;
  assign n47236 = x173 & x217;
  assign n47237 = n47235 & n47236;
  assign n47238 = n47235 | n47236;
  assign n47239 = ~n47237 & n47238;
  assign n64804 = n47036 | n47038;
  assign n64821 = n47239 & n64804;
  assign n64822 = n47036 & n47239;
  assign n64823 = (n74102 & n64821) | (n74102 & n64822) | (n64821 & n64822);
  assign n64824 = n47239 | n64804;
  assign n64825 = n47036 | n47239;
  assign n64826 = (n74102 & n64824) | (n74102 & n64825) | (n64824 & n64825);
  assign n47242 = ~n64823 & n64826;
  assign n47243 = x172 & x218;
  assign n47244 = n47242 & n47243;
  assign n47245 = n47242 | n47243;
  assign n47246 = ~n47244 & n47245;
  assign n64827 = n47043 & n47246;
  assign n74149 = (n47246 & n64709) | (n47246 & n64827) | (n64709 & n64827);
  assign n74150 = (n47246 & n64708) | (n47246 & n64827) | (n64708 & n64827);
  assign n74151 = (n74044 & n74149) | (n74044 & n74150) | (n74149 & n74150);
  assign n64829 = n47043 | n47246;
  assign n74152 = n64709 | n64829;
  assign n74153 = n64708 | n64829;
  assign n74154 = (n74044 & n74152) | (n74044 & n74153) | (n74152 & n74153);
  assign n47249 = ~n74151 & n74154;
  assign n47250 = x171 & x219;
  assign n47251 = n47249 & n47250;
  assign n47252 = n47249 | n47250;
  assign n47253 = ~n47251 & n47252;
  assign n47254 = n74129 & n47253;
  assign n47255 = n74129 | n47253;
  assign n47256 = ~n47254 & n47255;
  assign n47257 = x170 & x220;
  assign n47258 = n47256 & n47257;
  assign n47259 = n47256 | n47257;
  assign n47260 = ~n47258 & n47259;
  assign n64799 = n47057 | n47059;
  assign n64831 = n47260 & n64799;
  assign n64832 = n47057 & n47260;
  assign n64833 = (n74097 & n64831) | (n74097 & n64832) | (n64831 & n64832);
  assign n64834 = n47260 | n64799;
  assign n64835 = n47057 | n47260;
  assign n64836 = (n74097 & n64834) | (n74097 & n64835) | (n64834 & n64835);
  assign n47263 = ~n64833 & n64836;
  assign n47264 = x169 & x221;
  assign n47265 = n47263 & n47264;
  assign n47266 = n47263 | n47264;
  assign n47267 = ~n47265 & n47266;
  assign n64837 = n47064 & n47267;
  assign n74155 = (n47267 & n64719) | (n47267 & n64837) | (n64719 & n64837);
  assign n74156 = (n47267 & n64718) | (n47267 & n64837) | (n64718 & n64837);
  assign n74157 = (n64555 & n74155) | (n64555 & n74156) | (n74155 & n74156);
  assign n64839 = n47064 | n47267;
  assign n74158 = n64719 | n64839;
  assign n74159 = n64718 | n64839;
  assign n74160 = (n64555 & n74158) | (n64555 & n74159) | (n74158 & n74159);
  assign n47270 = ~n74157 & n74160;
  assign n47271 = x168 & x222;
  assign n47272 = n47270 & n47271;
  assign n47273 = n47270 | n47271;
  assign n47274 = ~n47272 & n47273;
  assign n64797 = n47071 | n47073;
  assign n74161 = n47274 & n64797;
  assign n74123 = n46862 | n47071;
  assign n74124 = (n47071 & n47073) | (n47071 & n74123) | (n47073 & n74123);
  assign n74162 = n47274 & n74124;
  assign n74163 = (n74089 & n74161) | (n74089 & n74162) | (n74161 & n74162);
  assign n74164 = n47274 | n64797;
  assign n74165 = n47274 | n74124;
  assign n74166 = (n74089 & n74164) | (n74089 & n74165) | (n74164 & n74165);
  assign n47277 = ~n74163 & n74166;
  assign n47278 = x167 & x223;
  assign n47279 = n47277 & n47278;
  assign n47280 = n47277 | n47278;
  assign n47281 = ~n47279 & n47280;
  assign n64841 = n47078 & n47281;
  assign n74167 = (n47281 & n64728) | (n47281 & n64841) | (n64728 & n64841);
  assign n74168 = (n47080 & n47281) | (n47080 & n64841) | (n47281 & n64841);
  assign n74169 = (n64612 & n74167) | (n64612 & n74168) | (n74167 & n74168);
  assign n64843 = n47078 | n47281;
  assign n74170 = n64728 | n64843;
  assign n74171 = n47080 | n64843;
  assign n74172 = (n64612 & n74170) | (n64612 & n74171) | (n74170 & n74171);
  assign n47284 = ~n74169 & n74172;
  assign n47285 = x166 & x224;
  assign n47286 = n47284 & n47285;
  assign n47287 = n47284 | n47285;
  assign n47288 = ~n47286 & n47287;
  assign n64845 = n47085 & n47288;
  assign n64846 = (n47288 & n64733) | (n47288 & n64845) | (n64733 & n64845);
  assign n64847 = n47085 | n47288;
  assign n64848 = n64733 | n64847;
  assign n47291 = ~n64846 & n64848;
  assign n47292 = x165 & x225;
  assign n47293 = n47291 & n47292;
  assign n47294 = n47291 | n47292;
  assign n47295 = ~n47293 & n47294;
  assign n64849 = n47092 & n47295;
  assign n64850 = (n47295 & n64737) | (n47295 & n64849) | (n64737 & n64849);
  assign n64851 = n47092 | n47295;
  assign n64852 = n64737 | n64851;
  assign n47298 = ~n64850 & n64852;
  assign n47299 = x164 & x226;
  assign n47300 = n47298 & n47299;
  assign n47301 = n47298 | n47299;
  assign n47302 = ~n47300 & n47301;
  assign n64853 = n47099 & n47302;
  assign n64854 = (n47302 & n64741) | (n47302 & n64853) | (n64741 & n64853);
  assign n64855 = n47099 | n47302;
  assign n64856 = n64741 | n64855;
  assign n47305 = ~n64854 & n64856;
  assign n47306 = x163 & x227;
  assign n47307 = n47305 & n47306;
  assign n47308 = n47305 | n47306;
  assign n47309 = ~n47307 & n47308;
  assign n64857 = n47106 & n47309;
  assign n64858 = (n47309 & n64745) | (n47309 & n64857) | (n64745 & n64857);
  assign n64859 = n47106 | n47309;
  assign n64860 = n64745 | n64859;
  assign n47312 = ~n64858 & n64860;
  assign n47313 = x162 & x228;
  assign n47314 = n47312 & n47313;
  assign n47315 = n47312 | n47313;
  assign n47316 = ~n47314 & n47315;
  assign n64861 = n47113 & n47316;
  assign n64862 = (n47316 & n64749) | (n47316 & n64861) | (n64749 & n64861);
  assign n64863 = n47113 | n47316;
  assign n64864 = n64749 | n64863;
  assign n47319 = ~n64862 & n64864;
  assign n47320 = x161 & x229;
  assign n47321 = n47319 & n47320;
  assign n47322 = n47319 | n47320;
  assign n47323 = ~n47321 & n47322;
  assign n64865 = n47120 & n47323;
  assign n64866 = (n47323 & n64753) | (n47323 & n64865) | (n64753 & n64865);
  assign n64867 = n47120 | n47323;
  assign n64868 = n64753 | n64867;
  assign n47326 = ~n64866 & n64868;
  assign n47327 = x160 & x230;
  assign n47328 = n47326 & n47327;
  assign n47329 = n47326 | n47327;
  assign n47330 = ~n47328 & n47329;
  assign n64869 = n47127 & n47330;
  assign n64870 = (n47330 & n64757) | (n47330 & n64869) | (n64757 & n64869);
  assign n64871 = n47127 | n47330;
  assign n64872 = n64757 | n64871;
  assign n47333 = ~n64870 & n64872;
  assign n47334 = x159 & x231;
  assign n47335 = n47333 & n47334;
  assign n47336 = n47333 | n47334;
  assign n47337 = ~n47335 & n47336;
  assign n64873 = n47134 & n47337;
  assign n64874 = (n47337 & n64761) | (n47337 & n64873) | (n64761 & n64873);
  assign n64875 = n47134 | n47337;
  assign n64876 = n64761 | n64875;
  assign n47340 = ~n64874 & n64876;
  assign n47341 = x158 & x232;
  assign n47342 = n47340 & n47341;
  assign n47343 = n47340 | n47341;
  assign n47344 = ~n47342 & n47343;
  assign n64877 = n47141 & n47344;
  assign n64878 = (n47344 & n64765) | (n47344 & n64877) | (n64765 & n64877);
  assign n64879 = n47141 | n47344;
  assign n64880 = n64765 | n64879;
  assign n47347 = ~n64878 & n64880;
  assign n47348 = x157 & x233;
  assign n47349 = n47347 & n47348;
  assign n47350 = n47347 | n47348;
  assign n47351 = ~n47349 & n47350;
  assign n64881 = n47148 & n47351;
  assign n64882 = (n47351 & n64769) | (n47351 & n64881) | (n64769 & n64881);
  assign n64883 = n47148 | n47351;
  assign n64884 = n64769 | n64883;
  assign n47354 = ~n64882 & n64884;
  assign n47355 = x156 & x234;
  assign n47356 = n47354 & n47355;
  assign n47357 = n47354 | n47355;
  assign n47358 = ~n47356 & n47357;
  assign n64885 = n47155 & n47358;
  assign n64886 = (n47358 & n64773) | (n47358 & n64885) | (n64773 & n64885);
  assign n64887 = n47155 | n47358;
  assign n64888 = n64773 | n64887;
  assign n47361 = ~n64886 & n64888;
  assign n47362 = x155 & x235;
  assign n47363 = n47361 & n47362;
  assign n47364 = n47361 | n47362;
  assign n47365 = ~n47363 & n47364;
  assign n64889 = n47162 & n47365;
  assign n64890 = (n47365 & n64777) | (n47365 & n64889) | (n64777 & n64889);
  assign n64891 = n47162 | n47365;
  assign n64892 = n64777 | n64891;
  assign n47368 = ~n64890 & n64892;
  assign n47369 = x154 & x236;
  assign n47370 = n47368 & n47369;
  assign n47371 = n47368 | n47369;
  assign n47372 = ~n47370 & n47371;
  assign n64893 = n47169 & n47372;
  assign n64894 = (n47372 & n64781) | (n47372 & n64893) | (n64781 & n64893);
  assign n64895 = n47169 | n47372;
  assign n64896 = n64781 | n64895;
  assign n47375 = ~n64894 & n64896;
  assign n47376 = x153 & x237;
  assign n47377 = n47375 & n47376;
  assign n47378 = n47375 | n47376;
  assign n47379 = ~n47377 & n47378;
  assign n64897 = n47176 & n47379;
  assign n64898 = (n47379 & n64785) | (n47379 & n64897) | (n64785 & n64897);
  assign n64899 = n47176 | n47379;
  assign n64900 = n64785 | n64899;
  assign n47382 = ~n64898 & n64900;
  assign n47383 = x152 & x238;
  assign n47384 = n47382 & n47383;
  assign n47385 = n47382 | n47383;
  assign n47386 = ~n47384 & n47385;
  assign n64901 = n47183 & n47386;
  assign n64902 = (n47386 & n64789) | (n47386 & n64901) | (n64789 & n64901);
  assign n64903 = n47183 | n47386;
  assign n64904 = n64789 | n64903;
  assign n47389 = ~n64902 & n64904;
  assign n47390 = x151 & x239;
  assign n47391 = n47389 & n47390;
  assign n47392 = n47389 | n47390;
  assign n47393 = ~n47391 & n47392;
  assign n64905 = n47190 & n47393;
  assign n64906 = (n47393 & n64793) | (n47393 & n64905) | (n64793 & n64905);
  assign n64907 = n47190 | n47393;
  assign n64908 = n64793 | n64907;
  assign n47396 = ~n64906 & n64908;
  assign n64798 = (n74089 & n74124) | (n74089 & n64797) | (n74124 & n64797);
  assign n64912 = n47265 | n47267;
  assign n74173 = n47064 | n47265;
  assign n74174 = (n47265 & n47267) | (n47265 & n74173) | (n47267 & n74173);
  assign n74175 = (n64719 & n64912) | (n64719 & n74174) | (n64912 & n74174);
  assign n74176 = (n64718 & n64912) | (n64718 & n74174) | (n64912 & n74174);
  assign n74177 = (n64555 & n74175) | (n64555 & n74176) | (n74175 & n74176);
  assign n64917 = n47244 | n47246;
  assign n74178 = n47043 | n47244;
  assign n74179 = (n47244 & n47246) | (n47244 & n74178) | (n47246 & n74178);
  assign n74180 = (n64709 & n64917) | (n64709 & n74179) | (n64917 & n74179);
  assign n74181 = (n64708 & n64917) | (n64708 & n74179) | (n64917 & n74179);
  assign n74182 = (n74044 & n74180) | (n74044 & n74181) | (n74180 & n74181);
  assign n47422 = x175 & x216;
  assign n74183 = n47225 | n74141;
  assign n74184 = (n47022 & n74141) | (n47022 & n74183) | (n74141 & n74183);
  assign n64924 = n47422 & n74184;
  assign n74185 = n47422 & n74141;
  assign n74186 = (n47225 & n47422) | (n47225 & n74185) | (n47422 & n74185);
  assign n64926 = (n64700 & n64924) | (n64700 & n74186) | (n64924 & n74186);
  assign n64927 = n47422 | n74184;
  assign n74187 = n47422 | n74141;
  assign n74188 = n47225 | n74187;
  assign n64929 = (n64700 & n64927) | (n64700 & n74188) | (n64927 & n74188);
  assign n47425 = ~n64926 & n64929;
  assign n64931 = n47230 & n47425;
  assign n74189 = (n47232 & n47425) | (n47232 & n64931) | (n47425 & n64931);
  assign n64932 = (n74134 & n74189) | (n74134 & n64931) | (n74189 & n64931);
  assign n64934 = n47230 | n47425;
  assign n74190 = n47232 | n64934;
  assign n64935 = (n74134 & n74190) | (n74134 & n64934) | (n74190 & n64934);
  assign n47428 = ~n64932 & n64935;
  assign n47429 = x174 & x217;
  assign n47430 = n47428 & n47429;
  assign n47431 = n47428 | n47429;
  assign n47432 = ~n47430 & n47431;
  assign n64936 = n47237 & n47432;
  assign n74191 = (n47432 & n64822) | (n47432 & n64936) | (n64822 & n64936);
  assign n74192 = (n47432 & n64821) | (n47432 & n64936) | (n64821 & n64936);
  assign n74193 = (n74102 & n74191) | (n74102 & n74192) | (n74191 & n74192);
  assign n64938 = n47237 | n47432;
  assign n74194 = n64822 | n64938;
  assign n74195 = n64821 | n64938;
  assign n74196 = (n74102 & n74194) | (n74102 & n74195) | (n74194 & n74195);
  assign n47435 = ~n74193 & n74196;
  assign n47436 = x173 & x218;
  assign n47437 = n47435 & n47436;
  assign n47438 = n47435 | n47436;
  assign n47439 = ~n47437 & n47438;
  assign n47440 = n74182 & n47439;
  assign n47441 = n74182 | n47439;
  assign n47442 = ~n47440 & n47441;
  assign n47443 = x172 & x219;
  assign n47444 = n47442 & n47443;
  assign n47445 = n47442 | n47443;
  assign n47446 = ~n47444 & n47445;
  assign n64914 = n47251 | n47253;
  assign n64940 = n47446 & n64914;
  assign n64941 = n47251 & n47446;
  assign n64942 = (n74129 & n64940) | (n74129 & n64941) | (n64940 & n64941);
  assign n64943 = n47446 | n64914;
  assign n64944 = n47251 | n47446;
  assign n64945 = (n74129 & n64943) | (n74129 & n64944) | (n64943 & n64944);
  assign n47449 = ~n64942 & n64945;
  assign n47450 = x171 & x220;
  assign n47451 = n47449 & n47450;
  assign n47452 = n47449 | n47450;
  assign n47453 = ~n47451 & n47452;
  assign n64946 = n47258 & n47453;
  assign n74197 = (n47453 & n64832) | (n47453 & n64946) | (n64832 & n64946);
  assign n74198 = (n47453 & n64831) | (n47453 & n64946) | (n64831 & n64946);
  assign n74199 = (n74097 & n74197) | (n74097 & n74198) | (n74197 & n74198);
  assign n64948 = n47258 | n47453;
  assign n74200 = n64832 | n64948;
  assign n74201 = n64831 | n64948;
  assign n74202 = (n74097 & n74200) | (n74097 & n74201) | (n74200 & n74201);
  assign n47456 = ~n74199 & n74202;
  assign n47457 = x170 & x221;
  assign n47458 = n47456 & n47457;
  assign n47459 = n47456 | n47457;
  assign n47460 = ~n47458 & n47459;
  assign n47461 = n74177 & n47460;
  assign n47462 = n74177 | n47460;
  assign n47463 = ~n47461 & n47462;
  assign n47464 = x169 & x222;
  assign n47465 = n47463 & n47464;
  assign n47466 = n47463 | n47464;
  assign n47467 = ~n47465 & n47466;
  assign n64909 = n47272 | n47274;
  assign n64950 = n47467 & n64909;
  assign n64951 = n47272 & n47467;
  assign n64952 = (n64798 & n64950) | (n64798 & n64951) | (n64950 & n64951);
  assign n64953 = n47467 | n64909;
  assign n64954 = n47272 | n47467;
  assign n64955 = (n64798 & n64953) | (n64798 & n64954) | (n64953 & n64954);
  assign n47470 = ~n64952 & n64955;
  assign n47471 = x168 & x223;
  assign n47472 = n47470 & n47471;
  assign n47473 = n47470 | n47471;
  assign n47474 = ~n47472 & n47473;
  assign n64956 = n47279 & n47474;
  assign n64957 = (n47474 & n74169) | (n47474 & n64956) | (n74169 & n64956);
  assign n64958 = n47279 | n47474;
  assign n64959 = n74169 | n64958;
  assign n47477 = ~n64957 & n64959;
  assign n47478 = x167 & x224;
  assign n47479 = n47477 & n47478;
  assign n47480 = n47477 | n47478;
  assign n47481 = ~n47479 & n47480;
  assign n64960 = n47286 & n47481;
  assign n64961 = (n47481 & n64846) | (n47481 & n64960) | (n64846 & n64960);
  assign n64962 = n47286 | n47481;
  assign n64963 = n64846 | n64962;
  assign n47484 = ~n64961 & n64963;
  assign n47485 = x166 & x225;
  assign n47486 = n47484 & n47485;
  assign n47487 = n47484 | n47485;
  assign n47488 = ~n47486 & n47487;
  assign n64964 = n47293 & n47488;
  assign n64965 = (n47488 & n64850) | (n47488 & n64964) | (n64850 & n64964);
  assign n64966 = n47293 | n47488;
  assign n64967 = n64850 | n64966;
  assign n47491 = ~n64965 & n64967;
  assign n47492 = x165 & x226;
  assign n47493 = n47491 & n47492;
  assign n47494 = n47491 | n47492;
  assign n47495 = ~n47493 & n47494;
  assign n64968 = n47300 & n47495;
  assign n64969 = (n47495 & n64854) | (n47495 & n64968) | (n64854 & n64968);
  assign n64970 = n47300 | n47495;
  assign n64971 = n64854 | n64970;
  assign n47498 = ~n64969 & n64971;
  assign n47499 = x164 & x227;
  assign n47500 = n47498 & n47499;
  assign n47501 = n47498 | n47499;
  assign n47502 = ~n47500 & n47501;
  assign n64972 = n47307 & n47502;
  assign n64973 = (n47502 & n64858) | (n47502 & n64972) | (n64858 & n64972);
  assign n64974 = n47307 | n47502;
  assign n64975 = n64858 | n64974;
  assign n47505 = ~n64973 & n64975;
  assign n47506 = x163 & x228;
  assign n47507 = n47505 & n47506;
  assign n47508 = n47505 | n47506;
  assign n47509 = ~n47507 & n47508;
  assign n64976 = n47314 & n47509;
  assign n64977 = (n47509 & n64862) | (n47509 & n64976) | (n64862 & n64976);
  assign n64978 = n47314 | n47509;
  assign n64979 = n64862 | n64978;
  assign n47512 = ~n64977 & n64979;
  assign n47513 = x162 & x229;
  assign n47514 = n47512 & n47513;
  assign n47515 = n47512 | n47513;
  assign n47516 = ~n47514 & n47515;
  assign n64980 = n47321 & n47516;
  assign n64981 = (n47516 & n64866) | (n47516 & n64980) | (n64866 & n64980);
  assign n64982 = n47321 | n47516;
  assign n64983 = n64866 | n64982;
  assign n47519 = ~n64981 & n64983;
  assign n47520 = x161 & x230;
  assign n47521 = n47519 & n47520;
  assign n47522 = n47519 | n47520;
  assign n47523 = ~n47521 & n47522;
  assign n64984 = n47328 & n47523;
  assign n64985 = (n47523 & n64870) | (n47523 & n64984) | (n64870 & n64984);
  assign n64986 = n47328 | n47523;
  assign n64987 = n64870 | n64986;
  assign n47526 = ~n64985 & n64987;
  assign n47527 = x160 & x231;
  assign n47528 = n47526 & n47527;
  assign n47529 = n47526 | n47527;
  assign n47530 = ~n47528 & n47529;
  assign n64988 = n47335 & n47530;
  assign n64989 = (n47530 & n64874) | (n47530 & n64988) | (n64874 & n64988);
  assign n64990 = n47335 | n47530;
  assign n64991 = n64874 | n64990;
  assign n47533 = ~n64989 & n64991;
  assign n47534 = x159 & x232;
  assign n47535 = n47533 & n47534;
  assign n47536 = n47533 | n47534;
  assign n47537 = ~n47535 & n47536;
  assign n64992 = n47342 & n47537;
  assign n64993 = (n47537 & n64878) | (n47537 & n64992) | (n64878 & n64992);
  assign n64994 = n47342 | n47537;
  assign n64995 = n64878 | n64994;
  assign n47540 = ~n64993 & n64995;
  assign n47541 = x158 & x233;
  assign n47542 = n47540 & n47541;
  assign n47543 = n47540 | n47541;
  assign n47544 = ~n47542 & n47543;
  assign n64996 = n47349 & n47544;
  assign n64997 = (n47544 & n64882) | (n47544 & n64996) | (n64882 & n64996);
  assign n64998 = n47349 | n47544;
  assign n64999 = n64882 | n64998;
  assign n47547 = ~n64997 & n64999;
  assign n47548 = x157 & x234;
  assign n47549 = n47547 & n47548;
  assign n47550 = n47547 | n47548;
  assign n47551 = ~n47549 & n47550;
  assign n65000 = n47356 & n47551;
  assign n65001 = (n47551 & n64886) | (n47551 & n65000) | (n64886 & n65000);
  assign n65002 = n47356 | n47551;
  assign n65003 = n64886 | n65002;
  assign n47554 = ~n65001 & n65003;
  assign n47555 = x156 & x235;
  assign n47556 = n47554 & n47555;
  assign n47557 = n47554 | n47555;
  assign n47558 = ~n47556 & n47557;
  assign n65004 = n47363 & n47558;
  assign n65005 = (n47558 & n64890) | (n47558 & n65004) | (n64890 & n65004);
  assign n65006 = n47363 | n47558;
  assign n65007 = n64890 | n65006;
  assign n47561 = ~n65005 & n65007;
  assign n47562 = x155 & x236;
  assign n47563 = n47561 & n47562;
  assign n47564 = n47561 | n47562;
  assign n47565 = ~n47563 & n47564;
  assign n65008 = n47370 & n47565;
  assign n65009 = (n47565 & n64894) | (n47565 & n65008) | (n64894 & n65008);
  assign n65010 = n47370 | n47565;
  assign n65011 = n64894 | n65010;
  assign n47568 = ~n65009 & n65011;
  assign n47569 = x154 & x237;
  assign n47570 = n47568 & n47569;
  assign n47571 = n47568 | n47569;
  assign n47572 = ~n47570 & n47571;
  assign n65012 = n47377 & n47572;
  assign n65013 = (n47572 & n64898) | (n47572 & n65012) | (n64898 & n65012);
  assign n65014 = n47377 | n47572;
  assign n65015 = n64898 | n65014;
  assign n47575 = ~n65013 & n65015;
  assign n47576 = x153 & x238;
  assign n47577 = n47575 & n47576;
  assign n47578 = n47575 | n47576;
  assign n47579 = ~n47577 & n47578;
  assign n65016 = n47384 & n47579;
  assign n65017 = (n47579 & n64902) | (n47579 & n65016) | (n64902 & n65016);
  assign n65018 = n47384 | n47579;
  assign n65019 = n64902 | n65018;
  assign n47582 = ~n65017 & n65019;
  assign n47583 = x152 & x239;
  assign n47584 = n47582 & n47583;
  assign n47585 = n47582 | n47583;
  assign n47586 = ~n47584 & n47585;
  assign n65020 = n47391 & n47586;
  assign n65021 = (n47586 & n64906) | (n47586 & n65020) | (n64906 & n65020);
  assign n65022 = n47391 | n47586;
  assign n65023 = n64906 | n65022;
  assign n47589 = ~n65021 & n65023;
  assign n65030 = n47451 | n47453;
  assign n74205 = n47258 | n47451;
  assign n74206 = (n47451 & n47453) | (n47451 & n74205) | (n47453 & n74205);
  assign n74207 = (n64832 & n65030) | (n64832 & n74206) | (n65030 & n74206);
  assign n74208 = (n64831 & n65030) | (n64831 & n74206) | (n65030 & n74206);
  assign n74209 = (n74097 & n74207) | (n74097 & n74208) | (n74207 & n74208);
  assign n65035 = n47430 | n47432;
  assign n74210 = n47237 | n47430;
  assign n74211 = (n47430 & n47432) | (n47430 & n74210) | (n47432 & n74210);
  assign n74212 = (n64822 & n65035) | (n64822 & n74211) | (n65035 & n74211);
  assign n74213 = (n64821 & n65035) | (n64821 & n74211) | (n65035 & n74211);
  assign n74214 = (n74102 & n74212) | (n74102 & n74213) | (n74212 & n74213);
  assign n47614 = x175 & x217;
  assign n74215 = n47614 & n64924;
  assign n74216 = n47614 & n74186;
  assign n74217 = (n64700 & n74215) | (n64700 & n74216) | (n74215 & n74216);
  assign n74218 = (n47614 & n74189) | (n47614 & n74217) | (n74189 & n74217);
  assign n74219 = (n47614 & n64931) | (n47614 & n74217) | (n64931 & n74217);
  assign n74220 = (n74134 & n74218) | (n74134 & n74219) | (n74218 & n74219);
  assign n74221 = n47614 | n64924;
  assign n74222 = n47614 | n74186;
  assign n74223 = (n64700 & n74221) | (n64700 & n74222) | (n74221 & n74222);
  assign n74224 = n74189 | n74223;
  assign n74225 = n64931 | n74223;
  assign n74226 = (n74134 & n74224) | (n74134 & n74225) | (n74224 & n74225);
  assign n47617 = ~n74220 & n74226;
  assign n47618 = n74214 & n47617;
  assign n47619 = n74214 | n47617;
  assign n47620 = ~n47618 & n47619;
  assign n47621 = x174 & x218;
  assign n47622 = n47620 & n47621;
  assign n47623 = n47620 | n47621;
  assign n47624 = ~n47622 & n47623;
  assign n65032 = n47437 | n47439;
  assign n65041 = n47624 & n65032;
  assign n65042 = n47437 & n47624;
  assign n65043 = (n74182 & n65041) | (n74182 & n65042) | (n65041 & n65042);
  assign n65044 = n47624 | n65032;
  assign n65045 = n47437 | n47624;
  assign n65046 = (n74182 & n65044) | (n74182 & n65045) | (n65044 & n65045);
  assign n47627 = ~n65043 & n65046;
  assign n47628 = x173 & x219;
  assign n47629 = n47627 & n47628;
  assign n47630 = n47627 | n47628;
  assign n47631 = ~n47629 & n47630;
  assign n65047 = n47444 & n47631;
  assign n74227 = (n47631 & n64941) | (n47631 & n65047) | (n64941 & n65047);
  assign n74228 = (n47631 & n64940) | (n47631 & n65047) | (n64940 & n65047);
  assign n74229 = (n74129 & n74227) | (n74129 & n74228) | (n74227 & n74228);
  assign n65049 = n47444 | n47631;
  assign n74230 = n64941 | n65049;
  assign n74231 = n64940 | n65049;
  assign n74232 = (n74129 & n74230) | (n74129 & n74231) | (n74230 & n74231);
  assign n47634 = ~n74229 & n74232;
  assign n47635 = x172 & x220;
  assign n47636 = n47634 & n47635;
  assign n47637 = n47634 | n47635;
  assign n47638 = ~n47636 & n47637;
  assign n47639 = n74209 & n47638;
  assign n47640 = n74209 | n47638;
  assign n47641 = ~n47639 & n47640;
  assign n47642 = x171 & x221;
  assign n47643 = n47641 & n47642;
  assign n47644 = n47641 | n47642;
  assign n47645 = ~n47643 & n47644;
  assign n65027 = n47458 | n47460;
  assign n65051 = n47645 & n65027;
  assign n65052 = n47458 & n47645;
  assign n65053 = (n74177 & n65051) | (n74177 & n65052) | (n65051 & n65052);
  assign n65054 = n47645 | n65027;
  assign n65055 = n47458 | n47645;
  assign n65056 = (n74177 & n65054) | (n74177 & n65055) | (n65054 & n65055);
  assign n47648 = ~n65053 & n65056;
  assign n47649 = x170 & x222;
  assign n47650 = n47648 & n47649;
  assign n47651 = n47648 | n47649;
  assign n47652 = ~n47650 & n47651;
  assign n65057 = n47465 & n47652;
  assign n74233 = (n47652 & n64951) | (n47652 & n65057) | (n64951 & n65057);
  assign n74234 = (n47652 & n64950) | (n47652 & n65057) | (n64950 & n65057);
  assign n74235 = (n64798 & n74233) | (n64798 & n74234) | (n74233 & n74234);
  assign n65059 = n47465 | n47652;
  assign n74236 = n64951 | n65059;
  assign n74237 = n64950 | n65059;
  assign n74238 = (n64798 & n74236) | (n64798 & n74237) | (n74236 & n74237);
  assign n47655 = ~n74235 & n74238;
  assign n47656 = x169 & x223;
  assign n47657 = n47655 & n47656;
  assign n47658 = n47655 | n47656;
  assign n47659 = ~n47657 & n47658;
  assign n65025 = n47472 | n47474;
  assign n74239 = n47659 & n65025;
  assign n74203 = n47279 | n47472;
  assign n74204 = (n47472 & n47474) | (n47472 & n74203) | (n47474 & n74203);
  assign n74240 = n47659 & n74204;
  assign n74241 = (n74169 & n74239) | (n74169 & n74240) | (n74239 & n74240);
  assign n74242 = n47659 | n65025;
  assign n74243 = n47659 | n74204;
  assign n74244 = (n74169 & n74242) | (n74169 & n74243) | (n74242 & n74243);
  assign n47662 = ~n74241 & n74244;
  assign n47663 = x168 & x224;
  assign n47664 = n47662 & n47663;
  assign n47665 = n47662 | n47663;
  assign n47666 = ~n47664 & n47665;
  assign n65061 = n47479 & n47666;
  assign n74245 = (n47666 & n64960) | (n47666 & n65061) | (n64960 & n65061);
  assign n74246 = (n47481 & n47666) | (n47481 & n65061) | (n47666 & n65061);
  assign n74247 = (n64846 & n74245) | (n64846 & n74246) | (n74245 & n74246);
  assign n65063 = n47479 | n47666;
  assign n74248 = n64960 | n65063;
  assign n74249 = n47481 | n65063;
  assign n74250 = (n64846 & n74248) | (n64846 & n74249) | (n74248 & n74249);
  assign n47669 = ~n74247 & n74250;
  assign n47670 = x167 & x225;
  assign n47671 = n47669 & n47670;
  assign n47672 = n47669 | n47670;
  assign n47673 = ~n47671 & n47672;
  assign n65065 = n47486 & n47673;
  assign n65066 = (n47673 & n64965) | (n47673 & n65065) | (n64965 & n65065);
  assign n65067 = n47486 | n47673;
  assign n65068 = n64965 | n65067;
  assign n47676 = ~n65066 & n65068;
  assign n47677 = x166 & x226;
  assign n47678 = n47676 & n47677;
  assign n47679 = n47676 | n47677;
  assign n47680 = ~n47678 & n47679;
  assign n65069 = n47493 & n47680;
  assign n65070 = (n47680 & n64969) | (n47680 & n65069) | (n64969 & n65069);
  assign n65071 = n47493 | n47680;
  assign n65072 = n64969 | n65071;
  assign n47683 = ~n65070 & n65072;
  assign n47684 = x165 & x227;
  assign n47685 = n47683 & n47684;
  assign n47686 = n47683 | n47684;
  assign n47687 = ~n47685 & n47686;
  assign n65073 = n47500 & n47687;
  assign n65074 = (n47687 & n64973) | (n47687 & n65073) | (n64973 & n65073);
  assign n65075 = n47500 | n47687;
  assign n65076 = n64973 | n65075;
  assign n47690 = ~n65074 & n65076;
  assign n47691 = x164 & x228;
  assign n47692 = n47690 & n47691;
  assign n47693 = n47690 | n47691;
  assign n47694 = ~n47692 & n47693;
  assign n65077 = n47507 & n47694;
  assign n65078 = (n47694 & n64977) | (n47694 & n65077) | (n64977 & n65077);
  assign n65079 = n47507 | n47694;
  assign n65080 = n64977 | n65079;
  assign n47697 = ~n65078 & n65080;
  assign n47698 = x163 & x229;
  assign n47699 = n47697 & n47698;
  assign n47700 = n47697 | n47698;
  assign n47701 = ~n47699 & n47700;
  assign n65081 = n47514 & n47701;
  assign n65082 = (n47701 & n64981) | (n47701 & n65081) | (n64981 & n65081);
  assign n65083 = n47514 | n47701;
  assign n65084 = n64981 | n65083;
  assign n47704 = ~n65082 & n65084;
  assign n47705 = x162 & x230;
  assign n47706 = n47704 & n47705;
  assign n47707 = n47704 | n47705;
  assign n47708 = ~n47706 & n47707;
  assign n65085 = n47521 & n47708;
  assign n65086 = (n47708 & n64985) | (n47708 & n65085) | (n64985 & n65085);
  assign n65087 = n47521 | n47708;
  assign n65088 = n64985 | n65087;
  assign n47711 = ~n65086 & n65088;
  assign n47712 = x161 & x231;
  assign n47713 = n47711 & n47712;
  assign n47714 = n47711 | n47712;
  assign n47715 = ~n47713 & n47714;
  assign n65089 = n47528 & n47715;
  assign n65090 = (n47715 & n64989) | (n47715 & n65089) | (n64989 & n65089);
  assign n65091 = n47528 | n47715;
  assign n65092 = n64989 | n65091;
  assign n47718 = ~n65090 & n65092;
  assign n47719 = x160 & x232;
  assign n47720 = n47718 & n47719;
  assign n47721 = n47718 | n47719;
  assign n47722 = ~n47720 & n47721;
  assign n65093 = n47535 & n47722;
  assign n65094 = (n47722 & n64993) | (n47722 & n65093) | (n64993 & n65093);
  assign n65095 = n47535 | n47722;
  assign n65096 = n64993 | n65095;
  assign n47725 = ~n65094 & n65096;
  assign n47726 = x159 & x233;
  assign n47727 = n47725 & n47726;
  assign n47728 = n47725 | n47726;
  assign n47729 = ~n47727 & n47728;
  assign n65097 = n47542 & n47729;
  assign n65098 = (n47729 & n64997) | (n47729 & n65097) | (n64997 & n65097);
  assign n65099 = n47542 | n47729;
  assign n65100 = n64997 | n65099;
  assign n47732 = ~n65098 & n65100;
  assign n47733 = x158 & x234;
  assign n47734 = n47732 & n47733;
  assign n47735 = n47732 | n47733;
  assign n47736 = ~n47734 & n47735;
  assign n65101 = n47549 & n47736;
  assign n65102 = (n47736 & n65001) | (n47736 & n65101) | (n65001 & n65101);
  assign n65103 = n47549 | n47736;
  assign n65104 = n65001 | n65103;
  assign n47739 = ~n65102 & n65104;
  assign n47740 = x157 & x235;
  assign n47741 = n47739 & n47740;
  assign n47742 = n47739 | n47740;
  assign n47743 = ~n47741 & n47742;
  assign n65105 = n47556 & n47743;
  assign n65106 = (n47743 & n65005) | (n47743 & n65105) | (n65005 & n65105);
  assign n65107 = n47556 | n47743;
  assign n65108 = n65005 | n65107;
  assign n47746 = ~n65106 & n65108;
  assign n47747 = x156 & x236;
  assign n47748 = n47746 & n47747;
  assign n47749 = n47746 | n47747;
  assign n47750 = ~n47748 & n47749;
  assign n65109 = n47563 & n47750;
  assign n65110 = (n47750 & n65009) | (n47750 & n65109) | (n65009 & n65109);
  assign n65111 = n47563 | n47750;
  assign n65112 = n65009 | n65111;
  assign n47753 = ~n65110 & n65112;
  assign n47754 = x155 & x237;
  assign n47755 = n47753 & n47754;
  assign n47756 = n47753 | n47754;
  assign n47757 = ~n47755 & n47756;
  assign n65113 = n47570 & n47757;
  assign n65114 = (n47757 & n65013) | (n47757 & n65113) | (n65013 & n65113);
  assign n65115 = n47570 | n47757;
  assign n65116 = n65013 | n65115;
  assign n47760 = ~n65114 & n65116;
  assign n47761 = x154 & x238;
  assign n47762 = n47760 & n47761;
  assign n47763 = n47760 | n47761;
  assign n47764 = ~n47762 & n47763;
  assign n65117 = n47577 & n47764;
  assign n65118 = (n47764 & n65017) | (n47764 & n65117) | (n65017 & n65117);
  assign n65119 = n47577 | n47764;
  assign n65120 = n65017 | n65119;
  assign n47767 = ~n65118 & n65120;
  assign n47768 = x153 & x239;
  assign n47769 = n47767 & n47768;
  assign n47770 = n47767 | n47768;
  assign n47771 = ~n47769 & n47770;
  assign n65121 = n47584 & n47771;
  assign n65122 = (n47771 & n65021) | (n47771 & n65121) | (n65021 & n65121);
  assign n65123 = n47584 | n47771;
  assign n65124 = n65021 | n65123;
  assign n47774 = ~n65122 & n65124;
  assign n65026 = (n74169 & n74204) | (n74169 & n65025) | (n74204 & n65025);
  assign n65128 = n47650 | n47652;
  assign n74251 = n47465 | n47650;
  assign n74252 = (n47650 & n47652) | (n47650 & n74251) | (n47652 & n74251);
  assign n74253 = (n64951 & n65128) | (n64951 & n74252) | (n65128 & n74252);
  assign n74254 = (n64950 & n65128) | (n64950 & n74252) | (n65128 & n74252);
  assign n74255 = (n64798 & n74253) | (n64798 & n74254) | (n74253 & n74254);
  assign n65133 = n47629 | n47631;
  assign n74256 = n47444 | n47629;
  assign n74257 = (n47629 & n47631) | (n47629 & n74256) | (n47631 & n74256);
  assign n74258 = (n64941 & n65133) | (n64941 & n74257) | (n65133 & n74257);
  assign n74259 = (n64940 & n65133) | (n64940 & n74257) | (n65133 & n74257);
  assign n74260 = (n74129 & n74258) | (n74129 & n74259) | (n74258 & n74259);
  assign n47798 = x175 & x218;
  assign n74261 = n47798 & n74220;
  assign n74262 = (n47617 & n47798) | (n47617 & n74261) | (n47798 & n74261);
  assign n65138 = n47798 & n74220;
  assign n65139 = (n74214 & n74262) | (n74214 & n65138) | (n74262 & n65138);
  assign n74263 = n47798 | n74220;
  assign n74264 = n47617 | n74263;
  assign n65141 = n47798 | n74220;
  assign n65142 = (n74214 & n74264) | (n74214 & n65141) | (n74264 & n65141);
  assign n47801 = ~n65139 & n65142;
  assign n65143 = n47622 & n47801;
  assign n74265 = (n47801 & n65042) | (n47801 & n65143) | (n65042 & n65143);
  assign n74266 = (n47801 & n65041) | (n47801 & n65143) | (n65041 & n65143);
  assign n74267 = (n74182 & n74265) | (n74182 & n74266) | (n74265 & n74266);
  assign n65145 = n47622 | n47801;
  assign n74268 = n65042 | n65145;
  assign n74269 = n65041 | n65145;
  assign n74270 = (n74182 & n74268) | (n74182 & n74269) | (n74268 & n74269);
  assign n47804 = ~n74267 & n74270;
  assign n47805 = x174 & x219;
  assign n47806 = n47804 & n47805;
  assign n47807 = n47804 | n47805;
  assign n47808 = ~n47806 & n47807;
  assign n47809 = n74260 & n47808;
  assign n47810 = n74260 | n47808;
  assign n47811 = ~n47809 & n47810;
  assign n47812 = x173 & x220;
  assign n47813 = n47811 & n47812;
  assign n47814 = n47811 | n47812;
  assign n47815 = ~n47813 & n47814;
  assign n65130 = n47636 | n47638;
  assign n65147 = n47815 & n65130;
  assign n65148 = n47636 & n47815;
  assign n65149 = (n74209 & n65147) | (n74209 & n65148) | (n65147 & n65148);
  assign n65150 = n47815 | n65130;
  assign n65151 = n47636 | n47815;
  assign n65152 = (n74209 & n65150) | (n74209 & n65151) | (n65150 & n65151);
  assign n47818 = ~n65149 & n65152;
  assign n47819 = x172 & x221;
  assign n47820 = n47818 & n47819;
  assign n47821 = n47818 | n47819;
  assign n47822 = ~n47820 & n47821;
  assign n65153 = n47643 & n47822;
  assign n74271 = (n47822 & n65052) | (n47822 & n65153) | (n65052 & n65153);
  assign n74272 = (n47822 & n65051) | (n47822 & n65153) | (n65051 & n65153);
  assign n74273 = (n74177 & n74271) | (n74177 & n74272) | (n74271 & n74272);
  assign n65155 = n47643 | n47822;
  assign n74274 = n65052 | n65155;
  assign n74275 = n65051 | n65155;
  assign n74276 = (n74177 & n74274) | (n74177 & n74275) | (n74274 & n74275);
  assign n47825 = ~n74273 & n74276;
  assign n47826 = x171 & x222;
  assign n47827 = n47825 & n47826;
  assign n47828 = n47825 | n47826;
  assign n47829 = ~n47827 & n47828;
  assign n47830 = n74255 & n47829;
  assign n47831 = n74255 | n47829;
  assign n47832 = ~n47830 & n47831;
  assign n47833 = x170 & x223;
  assign n47834 = n47832 & n47833;
  assign n47835 = n47832 | n47833;
  assign n47836 = ~n47834 & n47835;
  assign n65125 = n47657 | n47659;
  assign n65157 = n47836 & n65125;
  assign n65158 = n47657 & n47836;
  assign n65159 = (n65026 & n65157) | (n65026 & n65158) | (n65157 & n65158);
  assign n65160 = n47836 | n65125;
  assign n65161 = n47657 | n47836;
  assign n65162 = (n65026 & n65160) | (n65026 & n65161) | (n65160 & n65161);
  assign n47839 = ~n65159 & n65162;
  assign n47840 = x169 & x224;
  assign n47841 = n47839 & n47840;
  assign n47842 = n47839 | n47840;
  assign n47843 = ~n47841 & n47842;
  assign n65163 = n47664 & n47843;
  assign n65164 = (n47843 & n74247) | (n47843 & n65163) | (n74247 & n65163);
  assign n65165 = n47664 | n47843;
  assign n65166 = n74247 | n65165;
  assign n47846 = ~n65164 & n65166;
  assign n47847 = x168 & x225;
  assign n47848 = n47846 & n47847;
  assign n47849 = n47846 | n47847;
  assign n47850 = ~n47848 & n47849;
  assign n65167 = n47671 & n47850;
  assign n65168 = (n47850 & n65066) | (n47850 & n65167) | (n65066 & n65167);
  assign n65169 = n47671 | n47850;
  assign n65170 = n65066 | n65169;
  assign n47853 = ~n65168 & n65170;
  assign n47854 = x167 & x226;
  assign n47855 = n47853 & n47854;
  assign n47856 = n47853 | n47854;
  assign n47857 = ~n47855 & n47856;
  assign n65171 = n47678 & n47857;
  assign n65172 = (n47857 & n65070) | (n47857 & n65171) | (n65070 & n65171);
  assign n65173 = n47678 | n47857;
  assign n65174 = n65070 | n65173;
  assign n47860 = ~n65172 & n65174;
  assign n47861 = x166 & x227;
  assign n47862 = n47860 & n47861;
  assign n47863 = n47860 | n47861;
  assign n47864 = ~n47862 & n47863;
  assign n65175 = n47685 & n47864;
  assign n65176 = (n47864 & n65074) | (n47864 & n65175) | (n65074 & n65175);
  assign n65177 = n47685 | n47864;
  assign n65178 = n65074 | n65177;
  assign n47867 = ~n65176 & n65178;
  assign n47868 = x165 & x228;
  assign n47869 = n47867 & n47868;
  assign n47870 = n47867 | n47868;
  assign n47871 = ~n47869 & n47870;
  assign n65179 = n47692 & n47871;
  assign n65180 = (n47871 & n65078) | (n47871 & n65179) | (n65078 & n65179);
  assign n65181 = n47692 | n47871;
  assign n65182 = n65078 | n65181;
  assign n47874 = ~n65180 & n65182;
  assign n47875 = x164 & x229;
  assign n47876 = n47874 & n47875;
  assign n47877 = n47874 | n47875;
  assign n47878 = ~n47876 & n47877;
  assign n65183 = n47699 & n47878;
  assign n65184 = (n47878 & n65082) | (n47878 & n65183) | (n65082 & n65183);
  assign n65185 = n47699 | n47878;
  assign n65186 = n65082 | n65185;
  assign n47881 = ~n65184 & n65186;
  assign n47882 = x163 & x230;
  assign n47883 = n47881 & n47882;
  assign n47884 = n47881 | n47882;
  assign n47885 = ~n47883 & n47884;
  assign n65187 = n47706 & n47885;
  assign n65188 = (n47885 & n65086) | (n47885 & n65187) | (n65086 & n65187);
  assign n65189 = n47706 | n47885;
  assign n65190 = n65086 | n65189;
  assign n47888 = ~n65188 & n65190;
  assign n47889 = x162 & x231;
  assign n47890 = n47888 & n47889;
  assign n47891 = n47888 | n47889;
  assign n47892 = ~n47890 & n47891;
  assign n65191 = n47713 & n47892;
  assign n65192 = (n47892 & n65090) | (n47892 & n65191) | (n65090 & n65191);
  assign n65193 = n47713 | n47892;
  assign n65194 = n65090 | n65193;
  assign n47895 = ~n65192 & n65194;
  assign n47896 = x161 & x232;
  assign n47897 = n47895 & n47896;
  assign n47898 = n47895 | n47896;
  assign n47899 = ~n47897 & n47898;
  assign n65195 = n47720 & n47899;
  assign n65196 = (n47899 & n65094) | (n47899 & n65195) | (n65094 & n65195);
  assign n65197 = n47720 | n47899;
  assign n65198 = n65094 | n65197;
  assign n47902 = ~n65196 & n65198;
  assign n47903 = x160 & x233;
  assign n47904 = n47902 & n47903;
  assign n47905 = n47902 | n47903;
  assign n47906 = ~n47904 & n47905;
  assign n65199 = n47727 & n47906;
  assign n65200 = (n47906 & n65098) | (n47906 & n65199) | (n65098 & n65199);
  assign n65201 = n47727 | n47906;
  assign n65202 = n65098 | n65201;
  assign n47909 = ~n65200 & n65202;
  assign n47910 = x159 & x234;
  assign n47911 = n47909 & n47910;
  assign n47912 = n47909 | n47910;
  assign n47913 = ~n47911 & n47912;
  assign n65203 = n47734 & n47913;
  assign n65204 = (n47913 & n65102) | (n47913 & n65203) | (n65102 & n65203);
  assign n65205 = n47734 | n47913;
  assign n65206 = n65102 | n65205;
  assign n47916 = ~n65204 & n65206;
  assign n47917 = x158 & x235;
  assign n47918 = n47916 & n47917;
  assign n47919 = n47916 | n47917;
  assign n47920 = ~n47918 & n47919;
  assign n65207 = n47741 & n47920;
  assign n65208 = (n47920 & n65106) | (n47920 & n65207) | (n65106 & n65207);
  assign n65209 = n47741 | n47920;
  assign n65210 = n65106 | n65209;
  assign n47923 = ~n65208 & n65210;
  assign n47924 = x157 & x236;
  assign n47925 = n47923 & n47924;
  assign n47926 = n47923 | n47924;
  assign n47927 = ~n47925 & n47926;
  assign n65211 = n47748 & n47927;
  assign n65212 = (n47927 & n65110) | (n47927 & n65211) | (n65110 & n65211);
  assign n65213 = n47748 | n47927;
  assign n65214 = n65110 | n65213;
  assign n47930 = ~n65212 & n65214;
  assign n47931 = x156 & x237;
  assign n47932 = n47930 & n47931;
  assign n47933 = n47930 | n47931;
  assign n47934 = ~n47932 & n47933;
  assign n65215 = n47755 & n47934;
  assign n65216 = (n47934 & n65114) | (n47934 & n65215) | (n65114 & n65215);
  assign n65217 = n47755 | n47934;
  assign n65218 = n65114 | n65217;
  assign n47937 = ~n65216 & n65218;
  assign n47938 = x155 & x238;
  assign n47939 = n47937 & n47938;
  assign n47940 = n47937 | n47938;
  assign n47941 = ~n47939 & n47940;
  assign n65219 = n47762 & n47941;
  assign n65220 = (n47941 & n65118) | (n47941 & n65219) | (n65118 & n65219);
  assign n65221 = n47762 | n47941;
  assign n65222 = n65118 | n65221;
  assign n47944 = ~n65220 & n65222;
  assign n47945 = x154 & x239;
  assign n47946 = n47944 & n47945;
  assign n47947 = n47944 | n47945;
  assign n47948 = ~n47946 & n47947;
  assign n65223 = n47769 & n47948;
  assign n65224 = (n47948 & n65122) | (n47948 & n65223) | (n65122 & n65223);
  assign n65225 = n47769 | n47948;
  assign n65226 = n65122 | n65225;
  assign n47951 = ~n65224 & n65226;
  assign n65233 = n47820 | n47822;
  assign n74279 = n47643 | n47820;
  assign n74280 = (n47820 & n47822) | (n47820 & n74279) | (n47822 & n74279);
  assign n74281 = (n65052 & n65233) | (n65052 & n74280) | (n65233 & n74280);
  assign n74282 = (n65051 & n65233) | (n65051 & n74280) | (n65233 & n74280);
  assign n74283 = (n74177 & n74281) | (n74177 & n74282) | (n74281 & n74282);
  assign n47974 = x175 & x219;
  assign n65238 = n47801 | n65139;
  assign n74284 = (n47622 & n65139) | (n47622 & n65238) | (n65139 & n65238);
  assign n65240 = n47974 & n74284;
  assign n74285 = n47974 & n65139;
  assign n74286 = (n47801 & n47974) | (n47801 & n74285) | (n47974 & n74285);
  assign n74287 = (n65042 & n65240) | (n65042 & n74286) | (n65240 & n74286);
  assign n74288 = (n65041 & n65240) | (n65041 & n74286) | (n65240 & n74286);
  assign n74289 = (n74182 & n74287) | (n74182 & n74288) | (n74287 & n74288);
  assign n65243 = n47974 | n74284;
  assign n74290 = n47974 | n65139;
  assign n74291 = n47801 | n74290;
  assign n74292 = (n65042 & n65243) | (n65042 & n74291) | (n65243 & n74291);
  assign n74293 = (n65041 & n65243) | (n65041 & n74291) | (n65243 & n74291);
  assign n74294 = (n74182 & n74292) | (n74182 & n74293) | (n74292 & n74293);
  assign n47977 = ~n74289 & n74294;
  assign n65247 = n47806 & n47977;
  assign n74295 = (n47808 & n47977) | (n47808 & n65247) | (n47977 & n65247);
  assign n65248 = (n74260 & n74295) | (n74260 & n65247) | (n74295 & n65247);
  assign n65250 = n47806 | n47977;
  assign n74296 = n47808 | n65250;
  assign n65251 = (n74260 & n74296) | (n74260 & n65250) | (n74296 & n65250);
  assign n47980 = ~n65248 & n65251;
  assign n47981 = x174 & x220;
  assign n47982 = n47980 & n47981;
  assign n47983 = n47980 | n47981;
  assign n47984 = ~n47982 & n47983;
  assign n65252 = n47813 & n47984;
  assign n74297 = (n47984 & n65148) | (n47984 & n65252) | (n65148 & n65252);
  assign n74298 = (n47984 & n65147) | (n47984 & n65252) | (n65147 & n65252);
  assign n74299 = (n74209 & n74297) | (n74209 & n74298) | (n74297 & n74298);
  assign n65254 = n47813 | n47984;
  assign n74300 = n65148 | n65254;
  assign n74301 = n65147 | n65254;
  assign n74302 = (n74209 & n74300) | (n74209 & n74301) | (n74300 & n74301);
  assign n47987 = ~n74299 & n74302;
  assign n47988 = x173 & x221;
  assign n47989 = n47987 & n47988;
  assign n47990 = n47987 | n47988;
  assign n47991 = ~n47989 & n47990;
  assign n47992 = n74283 & n47991;
  assign n47993 = n74283 | n47991;
  assign n47994 = ~n47992 & n47993;
  assign n47995 = x172 & x222;
  assign n47996 = n47994 & n47995;
  assign n47997 = n47994 | n47995;
  assign n47998 = ~n47996 & n47997;
  assign n65230 = n47827 | n47829;
  assign n65256 = n47998 & n65230;
  assign n65257 = n47827 & n47998;
  assign n65258 = (n74255 & n65256) | (n74255 & n65257) | (n65256 & n65257);
  assign n65259 = n47998 | n65230;
  assign n65260 = n47827 | n47998;
  assign n65261 = (n74255 & n65259) | (n74255 & n65260) | (n65259 & n65260);
  assign n48001 = ~n65258 & n65261;
  assign n48002 = x171 & x223;
  assign n48003 = n48001 & n48002;
  assign n48004 = n48001 | n48002;
  assign n48005 = ~n48003 & n48004;
  assign n65262 = n47834 & n48005;
  assign n74303 = (n48005 & n65158) | (n48005 & n65262) | (n65158 & n65262);
  assign n74304 = (n48005 & n65157) | (n48005 & n65262) | (n65157 & n65262);
  assign n74305 = (n65026 & n74303) | (n65026 & n74304) | (n74303 & n74304);
  assign n65264 = n47834 | n48005;
  assign n74306 = n65158 | n65264;
  assign n74307 = n65157 | n65264;
  assign n74308 = (n65026 & n74306) | (n65026 & n74307) | (n74306 & n74307);
  assign n48008 = ~n74305 & n74308;
  assign n48009 = x170 & x224;
  assign n48010 = n48008 & n48009;
  assign n48011 = n48008 | n48009;
  assign n48012 = ~n48010 & n48011;
  assign n65228 = n47841 | n47843;
  assign n74309 = n48012 & n65228;
  assign n74277 = n47664 | n47841;
  assign n74278 = (n47841 & n47843) | (n47841 & n74277) | (n47843 & n74277);
  assign n74310 = n48012 & n74278;
  assign n74311 = (n74247 & n74309) | (n74247 & n74310) | (n74309 & n74310);
  assign n74312 = n48012 | n65228;
  assign n74313 = n48012 | n74278;
  assign n74314 = (n74247 & n74312) | (n74247 & n74313) | (n74312 & n74313);
  assign n48015 = ~n74311 & n74314;
  assign n48016 = x169 & x225;
  assign n48017 = n48015 & n48016;
  assign n48018 = n48015 | n48016;
  assign n48019 = ~n48017 & n48018;
  assign n65266 = n47848 & n48019;
  assign n74315 = (n48019 & n65167) | (n48019 & n65266) | (n65167 & n65266);
  assign n74316 = (n47850 & n48019) | (n47850 & n65266) | (n48019 & n65266);
  assign n74317 = (n65066 & n74315) | (n65066 & n74316) | (n74315 & n74316);
  assign n65268 = n47848 | n48019;
  assign n74318 = n65167 | n65268;
  assign n74319 = n47850 | n65268;
  assign n74320 = (n65066 & n74318) | (n65066 & n74319) | (n74318 & n74319);
  assign n48022 = ~n74317 & n74320;
  assign n48023 = x168 & x226;
  assign n48024 = n48022 & n48023;
  assign n48025 = n48022 | n48023;
  assign n48026 = ~n48024 & n48025;
  assign n65270 = n47855 & n48026;
  assign n65271 = (n48026 & n65172) | (n48026 & n65270) | (n65172 & n65270);
  assign n65272 = n47855 | n48026;
  assign n65273 = n65172 | n65272;
  assign n48029 = ~n65271 & n65273;
  assign n48030 = x167 & x227;
  assign n48031 = n48029 & n48030;
  assign n48032 = n48029 | n48030;
  assign n48033 = ~n48031 & n48032;
  assign n65274 = n47862 & n48033;
  assign n65275 = (n48033 & n65176) | (n48033 & n65274) | (n65176 & n65274);
  assign n65276 = n47862 | n48033;
  assign n65277 = n65176 | n65276;
  assign n48036 = ~n65275 & n65277;
  assign n48037 = x166 & x228;
  assign n48038 = n48036 & n48037;
  assign n48039 = n48036 | n48037;
  assign n48040 = ~n48038 & n48039;
  assign n65278 = n47869 & n48040;
  assign n65279 = (n48040 & n65180) | (n48040 & n65278) | (n65180 & n65278);
  assign n65280 = n47869 | n48040;
  assign n65281 = n65180 | n65280;
  assign n48043 = ~n65279 & n65281;
  assign n48044 = x165 & x229;
  assign n48045 = n48043 & n48044;
  assign n48046 = n48043 | n48044;
  assign n48047 = ~n48045 & n48046;
  assign n65282 = n47876 & n48047;
  assign n65283 = (n48047 & n65184) | (n48047 & n65282) | (n65184 & n65282);
  assign n65284 = n47876 | n48047;
  assign n65285 = n65184 | n65284;
  assign n48050 = ~n65283 & n65285;
  assign n48051 = x164 & x230;
  assign n48052 = n48050 & n48051;
  assign n48053 = n48050 | n48051;
  assign n48054 = ~n48052 & n48053;
  assign n65286 = n47883 & n48054;
  assign n65287 = (n48054 & n65188) | (n48054 & n65286) | (n65188 & n65286);
  assign n65288 = n47883 | n48054;
  assign n65289 = n65188 | n65288;
  assign n48057 = ~n65287 & n65289;
  assign n48058 = x163 & x231;
  assign n48059 = n48057 & n48058;
  assign n48060 = n48057 | n48058;
  assign n48061 = ~n48059 & n48060;
  assign n65290 = n47890 & n48061;
  assign n65291 = (n48061 & n65192) | (n48061 & n65290) | (n65192 & n65290);
  assign n65292 = n47890 | n48061;
  assign n65293 = n65192 | n65292;
  assign n48064 = ~n65291 & n65293;
  assign n48065 = x162 & x232;
  assign n48066 = n48064 & n48065;
  assign n48067 = n48064 | n48065;
  assign n48068 = ~n48066 & n48067;
  assign n65294 = n47897 & n48068;
  assign n65295 = (n48068 & n65196) | (n48068 & n65294) | (n65196 & n65294);
  assign n65296 = n47897 | n48068;
  assign n65297 = n65196 | n65296;
  assign n48071 = ~n65295 & n65297;
  assign n48072 = x161 & x233;
  assign n48073 = n48071 & n48072;
  assign n48074 = n48071 | n48072;
  assign n48075 = ~n48073 & n48074;
  assign n65298 = n47904 & n48075;
  assign n65299 = (n48075 & n65200) | (n48075 & n65298) | (n65200 & n65298);
  assign n65300 = n47904 | n48075;
  assign n65301 = n65200 | n65300;
  assign n48078 = ~n65299 & n65301;
  assign n48079 = x160 & x234;
  assign n48080 = n48078 & n48079;
  assign n48081 = n48078 | n48079;
  assign n48082 = ~n48080 & n48081;
  assign n65302 = n47911 & n48082;
  assign n65303 = (n48082 & n65204) | (n48082 & n65302) | (n65204 & n65302);
  assign n65304 = n47911 | n48082;
  assign n65305 = n65204 | n65304;
  assign n48085 = ~n65303 & n65305;
  assign n48086 = x159 & x235;
  assign n48087 = n48085 & n48086;
  assign n48088 = n48085 | n48086;
  assign n48089 = ~n48087 & n48088;
  assign n65306 = n47918 & n48089;
  assign n65307 = (n48089 & n65208) | (n48089 & n65306) | (n65208 & n65306);
  assign n65308 = n47918 | n48089;
  assign n65309 = n65208 | n65308;
  assign n48092 = ~n65307 & n65309;
  assign n48093 = x158 & x236;
  assign n48094 = n48092 & n48093;
  assign n48095 = n48092 | n48093;
  assign n48096 = ~n48094 & n48095;
  assign n65310 = n47925 & n48096;
  assign n65311 = (n48096 & n65212) | (n48096 & n65310) | (n65212 & n65310);
  assign n65312 = n47925 | n48096;
  assign n65313 = n65212 | n65312;
  assign n48099 = ~n65311 & n65313;
  assign n48100 = x157 & x237;
  assign n48101 = n48099 & n48100;
  assign n48102 = n48099 | n48100;
  assign n48103 = ~n48101 & n48102;
  assign n65314 = n47932 & n48103;
  assign n65315 = (n48103 & n65216) | (n48103 & n65314) | (n65216 & n65314);
  assign n65316 = n47932 | n48103;
  assign n65317 = n65216 | n65316;
  assign n48106 = ~n65315 & n65317;
  assign n48107 = x156 & x238;
  assign n48108 = n48106 & n48107;
  assign n48109 = n48106 | n48107;
  assign n48110 = ~n48108 & n48109;
  assign n65318 = n47939 & n48110;
  assign n65319 = (n48110 & n65220) | (n48110 & n65318) | (n65220 & n65318);
  assign n65320 = n47939 | n48110;
  assign n65321 = n65220 | n65320;
  assign n48113 = ~n65319 & n65321;
  assign n48114 = x155 & x239;
  assign n48115 = n48113 & n48114;
  assign n48116 = n48113 | n48114;
  assign n48117 = ~n48115 & n48116;
  assign n65322 = n47946 & n48117;
  assign n65323 = (n48117 & n65224) | (n48117 & n65322) | (n65224 & n65322);
  assign n65324 = n47946 | n48117;
  assign n65325 = n65224 | n65324;
  assign n48120 = ~n65323 & n65325;
  assign n65229 = (n74247 & n74278) | (n74247 & n65228) | (n74278 & n65228);
  assign n65329 = n48003 | n48005;
  assign n74321 = n47834 | n48003;
  assign n74322 = (n48003 & n48005) | (n48003 & n74321) | (n48005 & n74321);
  assign n74323 = (n65158 & n65329) | (n65158 & n74322) | (n65329 & n74322);
  assign n74324 = (n65157 & n65329) | (n65157 & n74322) | (n65329 & n74322);
  assign n74325 = (n65026 & n74323) | (n65026 & n74324) | (n74323 & n74324);
  assign n65334 = n47982 | n47984;
  assign n74326 = n47813 | n47982;
  assign n74327 = (n47982 & n47984) | (n47982 & n74326) | (n47984 & n74326);
  assign n74328 = (n65148 & n65334) | (n65148 & n74327) | (n65334 & n74327);
  assign n74329 = (n65147 & n65334) | (n65147 & n74327) | (n65334 & n74327);
  assign n74330 = (n74209 & n74328) | (n74209 & n74329) | (n74328 & n74329);
  assign n48142 = x175 & x220;
  assign n65336 = n48142 & n74289;
  assign n74331 = (n48142 & n65336) | (n48142 & n74295) | (n65336 & n74295);
  assign n74332 = (n48142 & n65247) | (n48142 & n65336) | (n65247 & n65336);
  assign n74333 = (n74260 & n74331) | (n74260 & n74332) | (n74331 & n74332);
  assign n65338 = n48142 | n74289;
  assign n74334 = n65338 | n74295;
  assign n74335 = n65247 | n65338;
  assign n74336 = (n74260 & n74334) | (n74260 & n74335) | (n74334 & n74335);
  assign n48145 = ~n74333 & n74336;
  assign n48146 = n74330 & n48145;
  assign n48147 = n74330 | n48145;
  assign n48148 = ~n48146 & n48147;
  assign n48149 = x174 & x221;
  assign n48150 = n48148 & n48149;
  assign n48151 = n48148 | n48149;
  assign n48152 = ~n48150 & n48151;
  assign n65331 = n47989 | n47991;
  assign n65340 = n48152 & n65331;
  assign n65341 = n47989 & n48152;
  assign n65342 = (n74283 & n65340) | (n74283 & n65341) | (n65340 & n65341);
  assign n65343 = n48152 | n65331;
  assign n65344 = n47989 | n48152;
  assign n65345 = (n74283 & n65343) | (n74283 & n65344) | (n65343 & n65344);
  assign n48155 = ~n65342 & n65345;
  assign n48156 = x173 & x222;
  assign n48157 = n48155 & n48156;
  assign n48158 = n48155 | n48156;
  assign n48159 = ~n48157 & n48158;
  assign n65346 = n47996 & n48159;
  assign n74337 = (n48159 & n65257) | (n48159 & n65346) | (n65257 & n65346);
  assign n74338 = (n48159 & n65256) | (n48159 & n65346) | (n65256 & n65346);
  assign n74339 = (n74255 & n74337) | (n74255 & n74338) | (n74337 & n74338);
  assign n65348 = n47996 | n48159;
  assign n74340 = n65257 | n65348;
  assign n74341 = n65256 | n65348;
  assign n74342 = (n74255 & n74340) | (n74255 & n74341) | (n74340 & n74341);
  assign n48162 = ~n74339 & n74342;
  assign n48163 = x172 & x223;
  assign n48164 = n48162 & n48163;
  assign n48165 = n48162 | n48163;
  assign n48166 = ~n48164 & n48165;
  assign n48167 = n74325 & n48166;
  assign n48168 = n74325 | n48166;
  assign n48169 = ~n48167 & n48168;
  assign n48170 = x171 & x224;
  assign n48171 = n48169 & n48170;
  assign n48172 = n48169 | n48170;
  assign n48173 = ~n48171 & n48172;
  assign n65326 = n48010 | n48012;
  assign n65350 = n48173 & n65326;
  assign n65351 = n48010 & n48173;
  assign n65352 = (n65229 & n65350) | (n65229 & n65351) | (n65350 & n65351);
  assign n65353 = n48173 | n65326;
  assign n65354 = n48010 | n48173;
  assign n65355 = (n65229 & n65353) | (n65229 & n65354) | (n65353 & n65354);
  assign n48176 = ~n65352 & n65355;
  assign n48177 = x170 & x225;
  assign n48178 = n48176 & n48177;
  assign n48179 = n48176 | n48177;
  assign n48180 = ~n48178 & n48179;
  assign n65356 = n48017 & n48180;
  assign n65357 = (n48180 & n74317) | (n48180 & n65356) | (n74317 & n65356);
  assign n65358 = n48017 | n48180;
  assign n65359 = n74317 | n65358;
  assign n48183 = ~n65357 & n65359;
  assign n48184 = x169 & x226;
  assign n48185 = n48183 & n48184;
  assign n48186 = n48183 | n48184;
  assign n48187 = ~n48185 & n48186;
  assign n65360 = n48024 & n48187;
  assign n65361 = (n48187 & n65271) | (n48187 & n65360) | (n65271 & n65360);
  assign n65362 = n48024 | n48187;
  assign n65363 = n65271 | n65362;
  assign n48190 = ~n65361 & n65363;
  assign n48191 = x168 & x227;
  assign n48192 = n48190 & n48191;
  assign n48193 = n48190 | n48191;
  assign n48194 = ~n48192 & n48193;
  assign n65364 = n48031 & n48194;
  assign n65365 = (n48194 & n65275) | (n48194 & n65364) | (n65275 & n65364);
  assign n65366 = n48031 | n48194;
  assign n65367 = n65275 | n65366;
  assign n48197 = ~n65365 & n65367;
  assign n48198 = x167 & x228;
  assign n48199 = n48197 & n48198;
  assign n48200 = n48197 | n48198;
  assign n48201 = ~n48199 & n48200;
  assign n65368 = n48038 & n48201;
  assign n65369 = (n48201 & n65279) | (n48201 & n65368) | (n65279 & n65368);
  assign n65370 = n48038 | n48201;
  assign n65371 = n65279 | n65370;
  assign n48204 = ~n65369 & n65371;
  assign n48205 = x166 & x229;
  assign n48206 = n48204 & n48205;
  assign n48207 = n48204 | n48205;
  assign n48208 = ~n48206 & n48207;
  assign n65372 = n48045 & n48208;
  assign n65373 = (n48208 & n65283) | (n48208 & n65372) | (n65283 & n65372);
  assign n65374 = n48045 | n48208;
  assign n65375 = n65283 | n65374;
  assign n48211 = ~n65373 & n65375;
  assign n48212 = x165 & x230;
  assign n48213 = n48211 & n48212;
  assign n48214 = n48211 | n48212;
  assign n48215 = ~n48213 & n48214;
  assign n65376 = n48052 & n48215;
  assign n65377 = (n48215 & n65287) | (n48215 & n65376) | (n65287 & n65376);
  assign n65378 = n48052 | n48215;
  assign n65379 = n65287 | n65378;
  assign n48218 = ~n65377 & n65379;
  assign n48219 = x164 & x231;
  assign n48220 = n48218 & n48219;
  assign n48221 = n48218 | n48219;
  assign n48222 = ~n48220 & n48221;
  assign n65380 = n48059 & n48222;
  assign n65381 = (n48222 & n65291) | (n48222 & n65380) | (n65291 & n65380);
  assign n65382 = n48059 | n48222;
  assign n65383 = n65291 | n65382;
  assign n48225 = ~n65381 & n65383;
  assign n48226 = x163 & x232;
  assign n48227 = n48225 & n48226;
  assign n48228 = n48225 | n48226;
  assign n48229 = ~n48227 & n48228;
  assign n65384 = n48066 & n48229;
  assign n65385 = (n48229 & n65295) | (n48229 & n65384) | (n65295 & n65384);
  assign n65386 = n48066 | n48229;
  assign n65387 = n65295 | n65386;
  assign n48232 = ~n65385 & n65387;
  assign n48233 = x162 & x233;
  assign n48234 = n48232 & n48233;
  assign n48235 = n48232 | n48233;
  assign n48236 = ~n48234 & n48235;
  assign n65388 = n48073 & n48236;
  assign n65389 = (n48236 & n65299) | (n48236 & n65388) | (n65299 & n65388);
  assign n65390 = n48073 | n48236;
  assign n65391 = n65299 | n65390;
  assign n48239 = ~n65389 & n65391;
  assign n48240 = x161 & x234;
  assign n48241 = n48239 & n48240;
  assign n48242 = n48239 | n48240;
  assign n48243 = ~n48241 & n48242;
  assign n65392 = n48080 & n48243;
  assign n65393 = (n48243 & n65303) | (n48243 & n65392) | (n65303 & n65392);
  assign n65394 = n48080 | n48243;
  assign n65395 = n65303 | n65394;
  assign n48246 = ~n65393 & n65395;
  assign n48247 = x160 & x235;
  assign n48248 = n48246 & n48247;
  assign n48249 = n48246 | n48247;
  assign n48250 = ~n48248 & n48249;
  assign n65396 = n48087 & n48250;
  assign n65397 = (n48250 & n65307) | (n48250 & n65396) | (n65307 & n65396);
  assign n65398 = n48087 | n48250;
  assign n65399 = n65307 | n65398;
  assign n48253 = ~n65397 & n65399;
  assign n48254 = x159 & x236;
  assign n48255 = n48253 & n48254;
  assign n48256 = n48253 | n48254;
  assign n48257 = ~n48255 & n48256;
  assign n65400 = n48094 & n48257;
  assign n65401 = (n48257 & n65311) | (n48257 & n65400) | (n65311 & n65400);
  assign n65402 = n48094 | n48257;
  assign n65403 = n65311 | n65402;
  assign n48260 = ~n65401 & n65403;
  assign n48261 = x158 & x237;
  assign n48262 = n48260 & n48261;
  assign n48263 = n48260 | n48261;
  assign n48264 = ~n48262 & n48263;
  assign n65404 = n48101 & n48264;
  assign n65405 = (n48264 & n65315) | (n48264 & n65404) | (n65315 & n65404);
  assign n65406 = n48101 | n48264;
  assign n65407 = n65315 | n65406;
  assign n48267 = ~n65405 & n65407;
  assign n48268 = x157 & x238;
  assign n48269 = n48267 & n48268;
  assign n48270 = n48267 | n48268;
  assign n48271 = ~n48269 & n48270;
  assign n65408 = n48108 & n48271;
  assign n65409 = (n48271 & n65319) | (n48271 & n65408) | (n65319 & n65408);
  assign n65410 = n48108 | n48271;
  assign n65411 = n65319 | n65410;
  assign n48274 = ~n65409 & n65411;
  assign n48275 = x156 & x239;
  assign n48276 = n48274 & n48275;
  assign n48277 = n48274 | n48275;
  assign n48278 = ~n48276 & n48277;
  assign n65412 = n48115 & n48278;
  assign n65413 = (n48278 & n65323) | (n48278 & n65412) | (n65323 & n65412);
  assign n65414 = n48115 | n48278;
  assign n65415 = n65323 | n65414;
  assign n48281 = ~n65413 & n65415;
  assign n65422 = n48157 | n48159;
  assign n74345 = n47996 | n48157;
  assign n74346 = (n48157 & n48159) | (n48157 & n74345) | (n48159 & n74345);
  assign n74347 = (n65257 & n65422) | (n65257 & n74346) | (n65422 & n74346);
  assign n74348 = (n65256 & n65422) | (n65256 & n74346) | (n65422 & n74346);
  assign n74349 = (n74255 & n74347) | (n74255 & n74348) | (n74347 & n74348);
  assign n48302 = x175 & x221;
  assign n74350 = n48302 & n74333;
  assign n74351 = (n48145 & n48302) | (n48145 & n74350) | (n48302 & n74350);
  assign n74352 = n48302 & n74331;
  assign n74353 = n48302 & n74332;
  assign n74354 = (n74260 & n74352) | (n74260 & n74353) | (n74352 & n74353);
  assign n65428 = (n74330 & n74351) | (n74330 & n74354) | (n74351 & n74354);
  assign n74355 = n48302 | n74333;
  assign n74356 = n48145 | n74355;
  assign n74357 = n48302 | n74331;
  assign n74358 = n48302 | n74332;
  assign n74359 = (n74260 & n74357) | (n74260 & n74358) | (n74357 & n74358);
  assign n65431 = (n74330 & n74356) | (n74330 & n74359) | (n74356 & n74359);
  assign n48305 = ~n65428 & n65431;
  assign n65432 = n48150 & n48305;
  assign n74360 = (n48305 & n65341) | (n48305 & n65432) | (n65341 & n65432);
  assign n74361 = (n48305 & n65340) | (n48305 & n65432) | (n65340 & n65432);
  assign n74362 = (n74283 & n74360) | (n74283 & n74361) | (n74360 & n74361);
  assign n65434 = n48150 | n48305;
  assign n74363 = n65341 | n65434;
  assign n74364 = n65340 | n65434;
  assign n74365 = (n74283 & n74363) | (n74283 & n74364) | (n74363 & n74364);
  assign n48308 = ~n74362 & n74365;
  assign n48309 = x174 & x222;
  assign n48310 = n48308 & n48309;
  assign n48311 = n48308 | n48309;
  assign n48312 = ~n48310 & n48311;
  assign n48313 = n74349 & n48312;
  assign n48314 = n74349 | n48312;
  assign n48315 = ~n48313 & n48314;
  assign n48316 = x173 & x223;
  assign n48317 = n48315 & n48316;
  assign n48318 = n48315 | n48316;
  assign n48319 = ~n48317 & n48318;
  assign n65419 = n48164 | n48166;
  assign n65436 = n48319 & n65419;
  assign n65437 = n48164 & n48319;
  assign n65438 = (n74325 & n65436) | (n74325 & n65437) | (n65436 & n65437);
  assign n65439 = n48319 | n65419;
  assign n65440 = n48164 | n48319;
  assign n65441 = (n74325 & n65439) | (n74325 & n65440) | (n65439 & n65440);
  assign n48322 = ~n65438 & n65441;
  assign n48323 = x172 & x224;
  assign n48324 = n48322 & n48323;
  assign n48325 = n48322 | n48323;
  assign n48326 = ~n48324 & n48325;
  assign n65442 = n48171 & n48326;
  assign n74366 = (n48326 & n65351) | (n48326 & n65442) | (n65351 & n65442);
  assign n74367 = (n48326 & n65350) | (n48326 & n65442) | (n65350 & n65442);
  assign n74368 = (n65229 & n74366) | (n65229 & n74367) | (n74366 & n74367);
  assign n65444 = n48171 | n48326;
  assign n74369 = n65351 | n65444;
  assign n74370 = n65350 | n65444;
  assign n74371 = (n65229 & n74369) | (n65229 & n74370) | (n74369 & n74370);
  assign n48329 = ~n74368 & n74371;
  assign n48330 = x171 & x225;
  assign n48331 = n48329 & n48330;
  assign n48332 = n48329 | n48330;
  assign n48333 = ~n48331 & n48332;
  assign n65417 = n48178 | n48180;
  assign n74372 = n48333 & n65417;
  assign n74343 = n48017 | n48178;
  assign n74344 = (n48178 & n48180) | (n48178 & n74343) | (n48180 & n74343);
  assign n74373 = n48333 & n74344;
  assign n74374 = (n74317 & n74372) | (n74317 & n74373) | (n74372 & n74373);
  assign n74375 = n48333 | n65417;
  assign n74376 = n48333 | n74344;
  assign n74377 = (n74317 & n74375) | (n74317 & n74376) | (n74375 & n74376);
  assign n48336 = ~n74374 & n74377;
  assign n48337 = x170 & x226;
  assign n48338 = n48336 & n48337;
  assign n48339 = n48336 | n48337;
  assign n48340 = ~n48338 & n48339;
  assign n65446 = n48185 & n48340;
  assign n74378 = (n48340 & n65360) | (n48340 & n65446) | (n65360 & n65446);
  assign n74379 = (n48187 & n48340) | (n48187 & n65446) | (n48340 & n65446);
  assign n74380 = (n65271 & n74378) | (n65271 & n74379) | (n74378 & n74379);
  assign n65448 = n48185 | n48340;
  assign n74381 = n65360 | n65448;
  assign n74382 = n48187 | n65448;
  assign n74383 = (n65271 & n74381) | (n65271 & n74382) | (n74381 & n74382);
  assign n48343 = ~n74380 & n74383;
  assign n48344 = x169 & x227;
  assign n48345 = n48343 & n48344;
  assign n48346 = n48343 | n48344;
  assign n48347 = ~n48345 & n48346;
  assign n65450 = n48192 & n48347;
  assign n65451 = (n48347 & n65365) | (n48347 & n65450) | (n65365 & n65450);
  assign n65452 = n48192 | n48347;
  assign n65453 = n65365 | n65452;
  assign n48350 = ~n65451 & n65453;
  assign n48351 = x168 & x228;
  assign n48352 = n48350 & n48351;
  assign n48353 = n48350 | n48351;
  assign n48354 = ~n48352 & n48353;
  assign n65454 = n48199 & n48354;
  assign n65455 = (n48354 & n65369) | (n48354 & n65454) | (n65369 & n65454);
  assign n65456 = n48199 | n48354;
  assign n65457 = n65369 | n65456;
  assign n48357 = ~n65455 & n65457;
  assign n48358 = x167 & x229;
  assign n48359 = n48357 & n48358;
  assign n48360 = n48357 | n48358;
  assign n48361 = ~n48359 & n48360;
  assign n65458 = n48206 & n48361;
  assign n65459 = (n48361 & n65373) | (n48361 & n65458) | (n65373 & n65458);
  assign n65460 = n48206 | n48361;
  assign n65461 = n65373 | n65460;
  assign n48364 = ~n65459 & n65461;
  assign n48365 = x166 & x230;
  assign n48366 = n48364 & n48365;
  assign n48367 = n48364 | n48365;
  assign n48368 = ~n48366 & n48367;
  assign n65462 = n48213 & n48368;
  assign n65463 = (n48368 & n65377) | (n48368 & n65462) | (n65377 & n65462);
  assign n65464 = n48213 | n48368;
  assign n65465 = n65377 | n65464;
  assign n48371 = ~n65463 & n65465;
  assign n48372 = x165 & x231;
  assign n48373 = n48371 & n48372;
  assign n48374 = n48371 | n48372;
  assign n48375 = ~n48373 & n48374;
  assign n65466 = n48220 & n48375;
  assign n65467 = (n48375 & n65381) | (n48375 & n65466) | (n65381 & n65466);
  assign n65468 = n48220 | n48375;
  assign n65469 = n65381 | n65468;
  assign n48378 = ~n65467 & n65469;
  assign n48379 = x164 & x232;
  assign n48380 = n48378 & n48379;
  assign n48381 = n48378 | n48379;
  assign n48382 = ~n48380 & n48381;
  assign n65470 = n48227 & n48382;
  assign n65471 = (n48382 & n65385) | (n48382 & n65470) | (n65385 & n65470);
  assign n65472 = n48227 | n48382;
  assign n65473 = n65385 | n65472;
  assign n48385 = ~n65471 & n65473;
  assign n48386 = x163 & x233;
  assign n48387 = n48385 & n48386;
  assign n48388 = n48385 | n48386;
  assign n48389 = ~n48387 & n48388;
  assign n65474 = n48234 & n48389;
  assign n65475 = (n48389 & n65389) | (n48389 & n65474) | (n65389 & n65474);
  assign n65476 = n48234 | n48389;
  assign n65477 = n65389 | n65476;
  assign n48392 = ~n65475 & n65477;
  assign n48393 = x162 & x234;
  assign n48394 = n48392 & n48393;
  assign n48395 = n48392 | n48393;
  assign n48396 = ~n48394 & n48395;
  assign n65478 = n48241 & n48396;
  assign n65479 = (n48396 & n65393) | (n48396 & n65478) | (n65393 & n65478);
  assign n65480 = n48241 | n48396;
  assign n65481 = n65393 | n65480;
  assign n48399 = ~n65479 & n65481;
  assign n48400 = x161 & x235;
  assign n48401 = n48399 & n48400;
  assign n48402 = n48399 | n48400;
  assign n48403 = ~n48401 & n48402;
  assign n65482 = n48248 & n48403;
  assign n65483 = (n48403 & n65397) | (n48403 & n65482) | (n65397 & n65482);
  assign n65484 = n48248 | n48403;
  assign n65485 = n65397 | n65484;
  assign n48406 = ~n65483 & n65485;
  assign n48407 = x160 & x236;
  assign n48408 = n48406 & n48407;
  assign n48409 = n48406 | n48407;
  assign n48410 = ~n48408 & n48409;
  assign n65486 = n48255 & n48410;
  assign n65487 = (n48410 & n65401) | (n48410 & n65486) | (n65401 & n65486);
  assign n65488 = n48255 | n48410;
  assign n65489 = n65401 | n65488;
  assign n48413 = ~n65487 & n65489;
  assign n48414 = x159 & x237;
  assign n48415 = n48413 & n48414;
  assign n48416 = n48413 | n48414;
  assign n48417 = ~n48415 & n48416;
  assign n65490 = n48262 & n48417;
  assign n65491 = (n48417 & n65405) | (n48417 & n65490) | (n65405 & n65490);
  assign n65492 = n48262 | n48417;
  assign n65493 = n65405 | n65492;
  assign n48420 = ~n65491 & n65493;
  assign n48421 = x158 & x238;
  assign n48422 = n48420 & n48421;
  assign n48423 = n48420 | n48421;
  assign n48424 = ~n48422 & n48423;
  assign n65494 = n48269 & n48424;
  assign n65495 = (n48424 & n65409) | (n48424 & n65494) | (n65409 & n65494);
  assign n65496 = n48269 | n48424;
  assign n65497 = n65409 | n65496;
  assign n48427 = ~n65495 & n65497;
  assign n48428 = x157 & x239;
  assign n48429 = n48427 & n48428;
  assign n48430 = n48427 | n48428;
  assign n48431 = ~n48429 & n48430;
  assign n65498 = n48276 & n48431;
  assign n65499 = (n48431 & n65413) | (n48431 & n65498) | (n65413 & n65498);
  assign n65500 = n48276 | n48431;
  assign n65501 = n65413 | n65500;
  assign n48434 = ~n65499 & n65501;
  assign n65418 = (n74317 & n74344) | (n74317 & n65417) | (n74344 & n65417);
  assign n65505 = n48324 | n48326;
  assign n74384 = n48171 | n48324;
  assign n74385 = (n48324 & n48326) | (n48324 & n74384) | (n48326 & n74384);
  assign n74386 = (n65351 & n65505) | (n65351 & n74385) | (n65505 & n74385);
  assign n74387 = (n65350 & n65505) | (n65350 & n74385) | (n65505 & n74385);
  assign n74388 = (n65229 & n74386) | (n65229 & n74387) | (n74386 & n74387);
  assign n48454 = x175 & x222;
  assign n65510 = n48305 | n65428;
  assign n74389 = (n48150 & n65428) | (n48150 & n65510) | (n65428 & n65510);
  assign n65512 = n48454 & n74389;
  assign n74390 = n48454 & n65428;
  assign n74391 = (n48305 & n48454) | (n48305 & n74390) | (n48454 & n74390);
  assign n74392 = (n65341 & n65512) | (n65341 & n74391) | (n65512 & n74391);
  assign n74393 = (n65340 & n65512) | (n65340 & n74391) | (n65512 & n74391);
  assign n74394 = (n74283 & n74392) | (n74283 & n74393) | (n74392 & n74393);
  assign n65515 = n48454 | n74389;
  assign n74395 = n48454 | n65428;
  assign n74396 = n48305 | n74395;
  assign n74397 = (n65341 & n65515) | (n65341 & n74396) | (n65515 & n74396);
  assign n74398 = (n65340 & n65515) | (n65340 & n74396) | (n65515 & n74396);
  assign n74399 = (n74283 & n74397) | (n74283 & n74398) | (n74397 & n74398);
  assign n48457 = ~n74394 & n74399;
  assign n65519 = n48310 & n48457;
  assign n74400 = (n48312 & n48457) | (n48312 & n65519) | (n48457 & n65519);
  assign n65520 = (n74349 & n74400) | (n74349 & n65519) | (n74400 & n65519);
  assign n65522 = n48310 | n48457;
  assign n74401 = n48312 | n65522;
  assign n65523 = (n74349 & n74401) | (n74349 & n65522) | (n74401 & n65522);
  assign n48460 = ~n65520 & n65523;
  assign n48461 = x174 & x223;
  assign n48462 = n48460 & n48461;
  assign n48463 = n48460 | n48461;
  assign n48464 = ~n48462 & n48463;
  assign n65524 = n48317 & n48464;
  assign n74402 = (n48464 & n65437) | (n48464 & n65524) | (n65437 & n65524);
  assign n74403 = (n48464 & n65436) | (n48464 & n65524) | (n65436 & n65524);
  assign n74404 = (n74325 & n74402) | (n74325 & n74403) | (n74402 & n74403);
  assign n65526 = n48317 | n48464;
  assign n74405 = n65437 | n65526;
  assign n74406 = n65436 | n65526;
  assign n74407 = (n74325 & n74405) | (n74325 & n74406) | (n74405 & n74406);
  assign n48467 = ~n74404 & n74407;
  assign n48468 = x173 & x224;
  assign n48469 = n48467 & n48468;
  assign n48470 = n48467 | n48468;
  assign n48471 = ~n48469 & n48470;
  assign n48472 = n74388 & n48471;
  assign n48473 = n74388 | n48471;
  assign n48474 = ~n48472 & n48473;
  assign n48475 = x172 & x225;
  assign n48476 = n48474 & n48475;
  assign n48477 = n48474 | n48475;
  assign n48478 = ~n48476 & n48477;
  assign n65502 = n48331 | n48333;
  assign n65528 = n48478 & n65502;
  assign n65529 = n48331 & n48478;
  assign n65530 = (n65418 & n65528) | (n65418 & n65529) | (n65528 & n65529);
  assign n65531 = n48478 | n65502;
  assign n65532 = n48331 | n48478;
  assign n65533 = (n65418 & n65531) | (n65418 & n65532) | (n65531 & n65532);
  assign n48481 = ~n65530 & n65533;
  assign n48482 = x171 & x226;
  assign n48483 = n48481 & n48482;
  assign n48484 = n48481 | n48482;
  assign n48485 = ~n48483 & n48484;
  assign n65534 = n48338 & n48485;
  assign n65535 = (n48485 & n74380) | (n48485 & n65534) | (n74380 & n65534);
  assign n65536 = n48338 | n48485;
  assign n65537 = n74380 | n65536;
  assign n48488 = ~n65535 & n65537;
  assign n48489 = x170 & x227;
  assign n48490 = n48488 & n48489;
  assign n48491 = n48488 | n48489;
  assign n48492 = ~n48490 & n48491;
  assign n65538 = n48345 & n48492;
  assign n65539 = (n48492 & n65451) | (n48492 & n65538) | (n65451 & n65538);
  assign n65540 = n48345 | n48492;
  assign n65541 = n65451 | n65540;
  assign n48495 = ~n65539 & n65541;
  assign n48496 = x169 & x228;
  assign n48497 = n48495 & n48496;
  assign n48498 = n48495 | n48496;
  assign n48499 = ~n48497 & n48498;
  assign n65542 = n48352 & n48499;
  assign n65543 = (n48499 & n65455) | (n48499 & n65542) | (n65455 & n65542);
  assign n65544 = n48352 | n48499;
  assign n65545 = n65455 | n65544;
  assign n48502 = ~n65543 & n65545;
  assign n48503 = x168 & x229;
  assign n48504 = n48502 & n48503;
  assign n48505 = n48502 | n48503;
  assign n48506 = ~n48504 & n48505;
  assign n65546 = n48359 & n48506;
  assign n65547 = (n48506 & n65459) | (n48506 & n65546) | (n65459 & n65546);
  assign n65548 = n48359 | n48506;
  assign n65549 = n65459 | n65548;
  assign n48509 = ~n65547 & n65549;
  assign n48510 = x167 & x230;
  assign n48511 = n48509 & n48510;
  assign n48512 = n48509 | n48510;
  assign n48513 = ~n48511 & n48512;
  assign n65550 = n48366 & n48513;
  assign n65551 = (n48513 & n65463) | (n48513 & n65550) | (n65463 & n65550);
  assign n65552 = n48366 | n48513;
  assign n65553 = n65463 | n65552;
  assign n48516 = ~n65551 & n65553;
  assign n48517 = x166 & x231;
  assign n48518 = n48516 & n48517;
  assign n48519 = n48516 | n48517;
  assign n48520 = ~n48518 & n48519;
  assign n65554 = n48373 & n48520;
  assign n65555 = (n48520 & n65467) | (n48520 & n65554) | (n65467 & n65554);
  assign n65556 = n48373 | n48520;
  assign n65557 = n65467 | n65556;
  assign n48523 = ~n65555 & n65557;
  assign n48524 = x165 & x232;
  assign n48525 = n48523 & n48524;
  assign n48526 = n48523 | n48524;
  assign n48527 = ~n48525 & n48526;
  assign n65558 = n48380 & n48527;
  assign n65559 = (n48527 & n65471) | (n48527 & n65558) | (n65471 & n65558);
  assign n65560 = n48380 | n48527;
  assign n65561 = n65471 | n65560;
  assign n48530 = ~n65559 & n65561;
  assign n48531 = x164 & x233;
  assign n48532 = n48530 & n48531;
  assign n48533 = n48530 | n48531;
  assign n48534 = ~n48532 & n48533;
  assign n65562 = n48387 & n48534;
  assign n65563 = (n48534 & n65475) | (n48534 & n65562) | (n65475 & n65562);
  assign n65564 = n48387 | n48534;
  assign n65565 = n65475 | n65564;
  assign n48537 = ~n65563 & n65565;
  assign n48538 = x163 & x234;
  assign n48539 = n48537 & n48538;
  assign n48540 = n48537 | n48538;
  assign n48541 = ~n48539 & n48540;
  assign n65566 = n48394 & n48541;
  assign n65567 = (n48541 & n65479) | (n48541 & n65566) | (n65479 & n65566);
  assign n65568 = n48394 | n48541;
  assign n65569 = n65479 | n65568;
  assign n48544 = ~n65567 & n65569;
  assign n48545 = x162 & x235;
  assign n48546 = n48544 & n48545;
  assign n48547 = n48544 | n48545;
  assign n48548 = ~n48546 & n48547;
  assign n65570 = n48401 & n48548;
  assign n65571 = (n48548 & n65483) | (n48548 & n65570) | (n65483 & n65570);
  assign n65572 = n48401 | n48548;
  assign n65573 = n65483 | n65572;
  assign n48551 = ~n65571 & n65573;
  assign n48552 = x161 & x236;
  assign n48553 = n48551 & n48552;
  assign n48554 = n48551 | n48552;
  assign n48555 = ~n48553 & n48554;
  assign n65574 = n48408 & n48555;
  assign n65575 = (n48555 & n65487) | (n48555 & n65574) | (n65487 & n65574);
  assign n65576 = n48408 | n48555;
  assign n65577 = n65487 | n65576;
  assign n48558 = ~n65575 & n65577;
  assign n48559 = x160 & x237;
  assign n48560 = n48558 & n48559;
  assign n48561 = n48558 | n48559;
  assign n48562 = ~n48560 & n48561;
  assign n65578 = n48415 & n48562;
  assign n65579 = (n48562 & n65491) | (n48562 & n65578) | (n65491 & n65578);
  assign n65580 = n48415 | n48562;
  assign n65581 = n65491 | n65580;
  assign n48565 = ~n65579 & n65581;
  assign n48566 = x159 & x238;
  assign n48567 = n48565 & n48566;
  assign n48568 = n48565 | n48566;
  assign n48569 = ~n48567 & n48568;
  assign n65582 = n48422 & n48569;
  assign n65583 = (n48569 & n65495) | (n48569 & n65582) | (n65495 & n65582);
  assign n65584 = n48422 | n48569;
  assign n65585 = n65495 | n65584;
  assign n48572 = ~n65583 & n65585;
  assign n48573 = x158 & x239;
  assign n48574 = n48572 & n48573;
  assign n48575 = n48572 | n48573;
  assign n48576 = ~n48574 & n48575;
  assign n65586 = n48429 & n48576;
  assign n65587 = (n48576 & n65499) | (n48576 & n65586) | (n65499 & n65586);
  assign n65588 = n48429 | n48576;
  assign n65589 = n65499 | n65588;
  assign n48579 = ~n65587 & n65589;
  assign n65596 = n48462 | n48464;
  assign n74410 = n48317 | n48462;
  assign n74411 = (n48462 & n48464) | (n48462 & n74410) | (n48464 & n74410);
  assign n74412 = (n65437 & n65596) | (n65437 & n74411) | (n65596 & n74411);
  assign n74413 = (n65436 & n65596) | (n65436 & n74411) | (n65596 & n74411);
  assign n74414 = (n74325 & n74412) | (n74325 & n74413) | (n74412 & n74413);
  assign n48598 = x175 & x223;
  assign n65598 = n48598 & n74394;
  assign n74415 = (n48598 & n65598) | (n48598 & n74400) | (n65598 & n74400);
  assign n74416 = (n48598 & n65519) | (n48598 & n65598) | (n65519 & n65598);
  assign n74417 = (n74349 & n74415) | (n74349 & n74416) | (n74415 & n74416);
  assign n65600 = n48598 | n74394;
  assign n74418 = n65600 | n74400;
  assign n74419 = n65519 | n65600;
  assign n74420 = (n74349 & n74418) | (n74349 & n74419) | (n74418 & n74419);
  assign n48601 = ~n74417 & n74420;
  assign n48602 = n74414 & n48601;
  assign n48603 = n74414 | n48601;
  assign n48604 = ~n48602 & n48603;
  assign n48605 = x174 & x224;
  assign n48606 = n48604 & n48605;
  assign n48607 = n48604 | n48605;
  assign n48608 = ~n48606 & n48607;
  assign n65593 = n48469 | n48471;
  assign n65602 = n48608 & n65593;
  assign n65603 = n48469 & n48608;
  assign n65604 = (n74388 & n65602) | (n74388 & n65603) | (n65602 & n65603);
  assign n65605 = n48608 | n65593;
  assign n65606 = n48469 | n48608;
  assign n65607 = (n74388 & n65605) | (n74388 & n65606) | (n65605 & n65606);
  assign n48611 = ~n65604 & n65607;
  assign n48612 = x173 & x225;
  assign n48613 = n48611 & n48612;
  assign n48614 = n48611 | n48612;
  assign n48615 = ~n48613 & n48614;
  assign n65608 = n48476 & n48615;
  assign n74421 = (n48615 & n65529) | (n48615 & n65608) | (n65529 & n65608);
  assign n74422 = (n48615 & n65528) | (n48615 & n65608) | (n65528 & n65608);
  assign n74423 = (n65418 & n74421) | (n65418 & n74422) | (n74421 & n74422);
  assign n65610 = n48476 | n48615;
  assign n74424 = n65529 | n65610;
  assign n74425 = n65528 | n65610;
  assign n74426 = (n65418 & n74424) | (n65418 & n74425) | (n74424 & n74425);
  assign n48618 = ~n74423 & n74426;
  assign n48619 = x172 & x226;
  assign n48620 = n48618 & n48619;
  assign n48621 = n48618 | n48619;
  assign n48622 = ~n48620 & n48621;
  assign n65591 = n48483 | n48485;
  assign n74427 = n48622 & n65591;
  assign n74408 = n48338 | n48483;
  assign n74409 = (n48483 & n48485) | (n48483 & n74408) | (n48485 & n74408);
  assign n74428 = n48622 & n74409;
  assign n74429 = (n74380 & n74427) | (n74380 & n74428) | (n74427 & n74428);
  assign n74430 = n48622 | n65591;
  assign n74431 = n48622 | n74409;
  assign n74432 = (n74380 & n74430) | (n74380 & n74431) | (n74430 & n74431);
  assign n48625 = ~n74429 & n74432;
  assign n48626 = x171 & x227;
  assign n48627 = n48625 & n48626;
  assign n48628 = n48625 | n48626;
  assign n48629 = ~n48627 & n48628;
  assign n65612 = n48490 & n48629;
  assign n74433 = (n48629 & n65538) | (n48629 & n65612) | (n65538 & n65612);
  assign n74434 = (n48492 & n48629) | (n48492 & n65612) | (n48629 & n65612);
  assign n74435 = (n65451 & n74433) | (n65451 & n74434) | (n74433 & n74434);
  assign n65614 = n48490 | n48629;
  assign n74436 = n65538 | n65614;
  assign n74437 = n48492 | n65614;
  assign n74438 = (n65451 & n74436) | (n65451 & n74437) | (n74436 & n74437);
  assign n48632 = ~n74435 & n74438;
  assign n48633 = x170 & x228;
  assign n48634 = n48632 & n48633;
  assign n48635 = n48632 | n48633;
  assign n48636 = ~n48634 & n48635;
  assign n65616 = n48497 & n48636;
  assign n65617 = (n48636 & n65543) | (n48636 & n65616) | (n65543 & n65616);
  assign n65618 = n48497 | n48636;
  assign n65619 = n65543 | n65618;
  assign n48639 = ~n65617 & n65619;
  assign n48640 = x169 & x229;
  assign n48641 = n48639 & n48640;
  assign n48642 = n48639 | n48640;
  assign n48643 = ~n48641 & n48642;
  assign n65620 = n48504 & n48643;
  assign n65621 = (n48643 & n65547) | (n48643 & n65620) | (n65547 & n65620);
  assign n65622 = n48504 | n48643;
  assign n65623 = n65547 | n65622;
  assign n48646 = ~n65621 & n65623;
  assign n48647 = x168 & x230;
  assign n48648 = n48646 & n48647;
  assign n48649 = n48646 | n48647;
  assign n48650 = ~n48648 & n48649;
  assign n65624 = n48511 & n48650;
  assign n65625 = (n48650 & n65551) | (n48650 & n65624) | (n65551 & n65624);
  assign n65626 = n48511 | n48650;
  assign n65627 = n65551 | n65626;
  assign n48653 = ~n65625 & n65627;
  assign n48654 = x167 & x231;
  assign n48655 = n48653 & n48654;
  assign n48656 = n48653 | n48654;
  assign n48657 = ~n48655 & n48656;
  assign n65628 = n48518 & n48657;
  assign n65629 = (n48657 & n65555) | (n48657 & n65628) | (n65555 & n65628);
  assign n65630 = n48518 | n48657;
  assign n65631 = n65555 | n65630;
  assign n48660 = ~n65629 & n65631;
  assign n48661 = x166 & x232;
  assign n48662 = n48660 & n48661;
  assign n48663 = n48660 | n48661;
  assign n48664 = ~n48662 & n48663;
  assign n65632 = n48525 & n48664;
  assign n65633 = (n48664 & n65559) | (n48664 & n65632) | (n65559 & n65632);
  assign n65634 = n48525 | n48664;
  assign n65635 = n65559 | n65634;
  assign n48667 = ~n65633 & n65635;
  assign n48668 = x165 & x233;
  assign n48669 = n48667 & n48668;
  assign n48670 = n48667 | n48668;
  assign n48671 = ~n48669 & n48670;
  assign n65636 = n48532 & n48671;
  assign n65637 = (n48671 & n65563) | (n48671 & n65636) | (n65563 & n65636);
  assign n65638 = n48532 | n48671;
  assign n65639 = n65563 | n65638;
  assign n48674 = ~n65637 & n65639;
  assign n48675 = x164 & x234;
  assign n48676 = n48674 & n48675;
  assign n48677 = n48674 | n48675;
  assign n48678 = ~n48676 & n48677;
  assign n65640 = n48539 & n48678;
  assign n65641 = (n48678 & n65567) | (n48678 & n65640) | (n65567 & n65640);
  assign n65642 = n48539 | n48678;
  assign n65643 = n65567 | n65642;
  assign n48681 = ~n65641 & n65643;
  assign n48682 = x163 & x235;
  assign n48683 = n48681 & n48682;
  assign n48684 = n48681 | n48682;
  assign n48685 = ~n48683 & n48684;
  assign n65644 = n48546 & n48685;
  assign n65645 = (n48685 & n65571) | (n48685 & n65644) | (n65571 & n65644);
  assign n65646 = n48546 | n48685;
  assign n65647 = n65571 | n65646;
  assign n48688 = ~n65645 & n65647;
  assign n48689 = x162 & x236;
  assign n48690 = n48688 & n48689;
  assign n48691 = n48688 | n48689;
  assign n48692 = ~n48690 & n48691;
  assign n65648 = n48553 & n48692;
  assign n65649 = (n48692 & n65575) | (n48692 & n65648) | (n65575 & n65648);
  assign n65650 = n48553 | n48692;
  assign n65651 = n65575 | n65650;
  assign n48695 = ~n65649 & n65651;
  assign n48696 = x161 & x237;
  assign n48697 = n48695 & n48696;
  assign n48698 = n48695 | n48696;
  assign n48699 = ~n48697 & n48698;
  assign n65652 = n48560 & n48699;
  assign n65653 = (n48699 & n65579) | (n48699 & n65652) | (n65579 & n65652);
  assign n65654 = n48560 | n48699;
  assign n65655 = n65579 | n65654;
  assign n48702 = ~n65653 & n65655;
  assign n48703 = x160 & x238;
  assign n48704 = n48702 & n48703;
  assign n48705 = n48702 | n48703;
  assign n48706 = ~n48704 & n48705;
  assign n65656 = n48567 & n48706;
  assign n65657 = (n48706 & n65583) | (n48706 & n65656) | (n65583 & n65656);
  assign n65658 = n48567 | n48706;
  assign n65659 = n65583 | n65658;
  assign n48709 = ~n65657 & n65659;
  assign n48710 = x159 & x239;
  assign n48711 = n48709 & n48710;
  assign n48712 = n48709 | n48710;
  assign n48713 = ~n48711 & n48712;
  assign n65660 = n48574 & n48713;
  assign n65661 = (n48713 & n65587) | (n48713 & n65660) | (n65587 & n65660);
  assign n65662 = n48574 | n48713;
  assign n65663 = n65587 | n65662;
  assign n48716 = ~n65661 & n65663;
  assign n65592 = (n74380 & n74409) | (n74380 & n65591) | (n74409 & n65591);
  assign n65667 = n48613 | n48615;
  assign n74439 = n48476 | n48613;
  assign n74440 = (n48613 & n48615) | (n48613 & n74439) | (n48615 & n74439);
  assign n74441 = (n65529 & n65667) | (n65529 & n74440) | (n65667 & n74440);
  assign n74442 = (n65528 & n65667) | (n65528 & n74440) | (n65667 & n74440);
  assign n74443 = (n65418 & n74441) | (n65418 & n74442) | (n74441 & n74442);
  assign n48734 = x175 & x224;
  assign n74444 = n48734 & n74417;
  assign n74445 = (n48601 & n48734) | (n48601 & n74444) | (n48734 & n74444);
  assign n74446 = n48734 & n74415;
  assign n74447 = n48734 & n74416;
  assign n74448 = (n74349 & n74446) | (n74349 & n74447) | (n74446 & n74447);
  assign n65673 = (n74414 & n74445) | (n74414 & n74448) | (n74445 & n74448);
  assign n74449 = n48734 | n74417;
  assign n74450 = n48601 | n74449;
  assign n74451 = n48734 | n74415;
  assign n74452 = n48734 | n74416;
  assign n74453 = (n74349 & n74451) | (n74349 & n74452) | (n74451 & n74452);
  assign n65676 = (n74414 & n74450) | (n74414 & n74453) | (n74450 & n74453);
  assign n48737 = ~n65673 & n65676;
  assign n65677 = n48606 & n48737;
  assign n74454 = (n48737 & n65603) | (n48737 & n65677) | (n65603 & n65677);
  assign n74455 = (n48737 & n65602) | (n48737 & n65677) | (n65602 & n65677);
  assign n74456 = (n74388 & n74454) | (n74388 & n74455) | (n74454 & n74455);
  assign n65679 = n48606 | n48737;
  assign n74457 = n65603 | n65679;
  assign n74458 = n65602 | n65679;
  assign n74459 = (n74388 & n74457) | (n74388 & n74458) | (n74457 & n74458);
  assign n48740 = ~n74456 & n74459;
  assign n48741 = x174 & x225;
  assign n48742 = n48740 & n48741;
  assign n48743 = n48740 | n48741;
  assign n48744 = ~n48742 & n48743;
  assign n48745 = n74443 & n48744;
  assign n48746 = n74443 | n48744;
  assign n48747 = ~n48745 & n48746;
  assign n48748 = x173 & x226;
  assign n48749 = n48747 & n48748;
  assign n48750 = n48747 | n48748;
  assign n48751 = ~n48749 & n48750;
  assign n65664 = n48620 | n48622;
  assign n65681 = n48751 & n65664;
  assign n65682 = n48620 & n48751;
  assign n65683 = (n65592 & n65681) | (n65592 & n65682) | (n65681 & n65682);
  assign n65684 = n48751 | n65664;
  assign n65685 = n48620 | n48751;
  assign n65686 = (n65592 & n65684) | (n65592 & n65685) | (n65684 & n65685);
  assign n48754 = ~n65683 & n65686;
  assign n48755 = x172 & x227;
  assign n48756 = n48754 & n48755;
  assign n48757 = n48754 | n48755;
  assign n48758 = ~n48756 & n48757;
  assign n65687 = n48627 & n48758;
  assign n65688 = (n48758 & n74435) | (n48758 & n65687) | (n74435 & n65687);
  assign n65689 = n48627 | n48758;
  assign n65690 = n74435 | n65689;
  assign n48761 = ~n65688 & n65690;
  assign n48762 = x171 & x228;
  assign n48763 = n48761 & n48762;
  assign n48764 = n48761 | n48762;
  assign n48765 = ~n48763 & n48764;
  assign n65691 = n48634 & n48765;
  assign n65692 = (n48765 & n65617) | (n48765 & n65691) | (n65617 & n65691);
  assign n65693 = n48634 | n48765;
  assign n65694 = n65617 | n65693;
  assign n48768 = ~n65692 & n65694;
  assign n48769 = x170 & x229;
  assign n48770 = n48768 & n48769;
  assign n48771 = n48768 | n48769;
  assign n48772 = ~n48770 & n48771;
  assign n65695 = n48641 & n48772;
  assign n65696 = (n48772 & n65621) | (n48772 & n65695) | (n65621 & n65695);
  assign n65697 = n48641 | n48772;
  assign n65698 = n65621 | n65697;
  assign n48775 = ~n65696 & n65698;
  assign n48776 = x169 & x230;
  assign n48777 = n48775 & n48776;
  assign n48778 = n48775 | n48776;
  assign n48779 = ~n48777 & n48778;
  assign n65699 = n48648 & n48779;
  assign n65700 = (n48779 & n65625) | (n48779 & n65699) | (n65625 & n65699);
  assign n65701 = n48648 | n48779;
  assign n65702 = n65625 | n65701;
  assign n48782 = ~n65700 & n65702;
  assign n48783 = x168 & x231;
  assign n48784 = n48782 & n48783;
  assign n48785 = n48782 | n48783;
  assign n48786 = ~n48784 & n48785;
  assign n65703 = n48655 & n48786;
  assign n65704 = (n48786 & n65629) | (n48786 & n65703) | (n65629 & n65703);
  assign n65705 = n48655 | n48786;
  assign n65706 = n65629 | n65705;
  assign n48789 = ~n65704 & n65706;
  assign n48790 = x167 & x232;
  assign n48791 = n48789 & n48790;
  assign n48792 = n48789 | n48790;
  assign n48793 = ~n48791 & n48792;
  assign n65707 = n48662 & n48793;
  assign n65708 = (n48793 & n65633) | (n48793 & n65707) | (n65633 & n65707);
  assign n65709 = n48662 | n48793;
  assign n65710 = n65633 | n65709;
  assign n48796 = ~n65708 & n65710;
  assign n48797 = x166 & x233;
  assign n48798 = n48796 & n48797;
  assign n48799 = n48796 | n48797;
  assign n48800 = ~n48798 & n48799;
  assign n65711 = n48669 & n48800;
  assign n65712 = (n48800 & n65637) | (n48800 & n65711) | (n65637 & n65711);
  assign n65713 = n48669 | n48800;
  assign n65714 = n65637 | n65713;
  assign n48803 = ~n65712 & n65714;
  assign n48804 = x165 & x234;
  assign n48805 = n48803 & n48804;
  assign n48806 = n48803 | n48804;
  assign n48807 = ~n48805 & n48806;
  assign n65715 = n48676 & n48807;
  assign n65716 = (n48807 & n65641) | (n48807 & n65715) | (n65641 & n65715);
  assign n65717 = n48676 | n48807;
  assign n65718 = n65641 | n65717;
  assign n48810 = ~n65716 & n65718;
  assign n48811 = x164 & x235;
  assign n48812 = n48810 & n48811;
  assign n48813 = n48810 | n48811;
  assign n48814 = ~n48812 & n48813;
  assign n65719 = n48683 & n48814;
  assign n65720 = (n48814 & n65645) | (n48814 & n65719) | (n65645 & n65719);
  assign n65721 = n48683 | n48814;
  assign n65722 = n65645 | n65721;
  assign n48817 = ~n65720 & n65722;
  assign n48818 = x163 & x236;
  assign n48819 = n48817 & n48818;
  assign n48820 = n48817 | n48818;
  assign n48821 = ~n48819 & n48820;
  assign n65723 = n48690 & n48821;
  assign n65724 = (n48821 & n65649) | (n48821 & n65723) | (n65649 & n65723);
  assign n65725 = n48690 | n48821;
  assign n65726 = n65649 | n65725;
  assign n48824 = ~n65724 & n65726;
  assign n48825 = x162 & x237;
  assign n48826 = n48824 & n48825;
  assign n48827 = n48824 | n48825;
  assign n48828 = ~n48826 & n48827;
  assign n65727 = n48697 & n48828;
  assign n65728 = (n48828 & n65653) | (n48828 & n65727) | (n65653 & n65727);
  assign n65729 = n48697 | n48828;
  assign n65730 = n65653 | n65729;
  assign n48831 = ~n65728 & n65730;
  assign n48832 = x161 & x238;
  assign n48833 = n48831 & n48832;
  assign n48834 = n48831 | n48832;
  assign n48835 = ~n48833 & n48834;
  assign n65731 = n48704 & n48835;
  assign n65732 = (n48835 & n65657) | (n48835 & n65731) | (n65657 & n65731);
  assign n65733 = n48704 | n48835;
  assign n65734 = n65657 | n65733;
  assign n48838 = ~n65732 & n65734;
  assign n48839 = x160 & x239;
  assign n48840 = n48838 & n48839;
  assign n48841 = n48838 | n48839;
  assign n48842 = ~n48840 & n48841;
  assign n65735 = n48711 & n48842;
  assign n65736 = (n48842 & n65661) | (n48842 & n65735) | (n65661 & n65735);
  assign n65737 = n48711 | n48842;
  assign n65738 = n65661 | n65737;
  assign n48845 = ~n65736 & n65738;
  assign n48862 = x175 & x225;
  assign n65745 = n48737 | n65673;
  assign n74462 = (n48606 & n65673) | (n48606 & n65745) | (n65673 & n65745);
  assign n65747 = n48862 & n74462;
  assign n74463 = n48862 & n65673;
  assign n74464 = (n48737 & n48862) | (n48737 & n74463) | (n48862 & n74463);
  assign n74465 = (n65603 & n65747) | (n65603 & n74464) | (n65747 & n74464);
  assign n74466 = (n65602 & n65747) | (n65602 & n74464) | (n65747 & n74464);
  assign n74467 = (n74388 & n74465) | (n74388 & n74466) | (n74465 & n74466);
  assign n65750 = n48862 | n74462;
  assign n74468 = n48862 | n65673;
  assign n74469 = n48737 | n74468;
  assign n74470 = (n65603 & n65750) | (n65603 & n74469) | (n65750 & n74469);
  assign n74471 = (n65602 & n65750) | (n65602 & n74469) | (n65750 & n74469);
  assign n74472 = (n74388 & n74470) | (n74388 & n74471) | (n74470 & n74471);
  assign n48865 = ~n74467 & n74472;
  assign n65754 = n48742 & n48865;
  assign n74473 = (n48744 & n48865) | (n48744 & n65754) | (n48865 & n65754);
  assign n65755 = (n74443 & n74473) | (n74443 & n65754) | (n74473 & n65754);
  assign n65757 = n48742 | n48865;
  assign n74474 = n48744 | n65757;
  assign n65758 = (n74443 & n74474) | (n74443 & n65757) | (n74474 & n65757);
  assign n48868 = ~n65755 & n65758;
  assign n48869 = x174 & x226;
  assign n48870 = n48868 & n48869;
  assign n48871 = n48868 | n48869;
  assign n48872 = ~n48870 & n48871;
  assign n65759 = n48749 & n48872;
  assign n74475 = (n48872 & n65682) | (n48872 & n65759) | (n65682 & n65759);
  assign n74476 = (n48872 & n65681) | (n48872 & n65759) | (n65681 & n65759);
  assign n74477 = (n65592 & n74475) | (n65592 & n74476) | (n74475 & n74476);
  assign n65761 = n48749 | n48872;
  assign n74478 = n65682 | n65761;
  assign n74479 = n65681 | n65761;
  assign n74480 = (n65592 & n74478) | (n65592 & n74479) | (n74478 & n74479);
  assign n48875 = ~n74477 & n74480;
  assign n48876 = x173 & x227;
  assign n48877 = n48875 & n48876;
  assign n48878 = n48875 | n48876;
  assign n48879 = ~n48877 & n48878;
  assign n65740 = n48756 | n48758;
  assign n74481 = n48879 & n65740;
  assign n74460 = n48627 | n48756;
  assign n74461 = (n48756 & n48758) | (n48756 & n74460) | (n48758 & n74460);
  assign n74482 = n48879 & n74461;
  assign n74483 = (n74435 & n74481) | (n74435 & n74482) | (n74481 & n74482);
  assign n74484 = n48879 | n65740;
  assign n74485 = n48879 | n74461;
  assign n74486 = (n74435 & n74484) | (n74435 & n74485) | (n74484 & n74485);
  assign n48882 = ~n74483 & n74486;
  assign n48883 = x172 & x228;
  assign n48884 = n48882 & n48883;
  assign n48885 = n48882 | n48883;
  assign n48886 = ~n48884 & n48885;
  assign n65763 = n48763 & n48886;
  assign n74487 = (n48886 & n65691) | (n48886 & n65763) | (n65691 & n65763);
  assign n74488 = (n48765 & n48886) | (n48765 & n65763) | (n48886 & n65763);
  assign n74489 = (n65617 & n74487) | (n65617 & n74488) | (n74487 & n74488);
  assign n65765 = n48763 | n48886;
  assign n74490 = n65691 | n65765;
  assign n74491 = n48765 | n65765;
  assign n74492 = (n65617 & n74490) | (n65617 & n74491) | (n74490 & n74491);
  assign n48889 = ~n74489 & n74492;
  assign n48890 = x171 & x229;
  assign n48891 = n48889 & n48890;
  assign n48892 = n48889 | n48890;
  assign n48893 = ~n48891 & n48892;
  assign n65767 = n48770 & n48893;
  assign n65768 = (n48893 & n65696) | (n48893 & n65767) | (n65696 & n65767);
  assign n65769 = n48770 | n48893;
  assign n65770 = n65696 | n65769;
  assign n48896 = ~n65768 & n65770;
  assign n48897 = x170 & x230;
  assign n48898 = n48896 & n48897;
  assign n48899 = n48896 | n48897;
  assign n48900 = ~n48898 & n48899;
  assign n65771 = n48777 & n48900;
  assign n65772 = (n48900 & n65700) | (n48900 & n65771) | (n65700 & n65771);
  assign n65773 = n48777 | n48900;
  assign n65774 = n65700 | n65773;
  assign n48903 = ~n65772 & n65774;
  assign n48904 = x169 & x231;
  assign n48905 = n48903 & n48904;
  assign n48906 = n48903 | n48904;
  assign n48907 = ~n48905 & n48906;
  assign n65775 = n48784 & n48907;
  assign n65776 = (n48907 & n65704) | (n48907 & n65775) | (n65704 & n65775);
  assign n65777 = n48784 | n48907;
  assign n65778 = n65704 | n65777;
  assign n48910 = ~n65776 & n65778;
  assign n48911 = x168 & x232;
  assign n48912 = n48910 & n48911;
  assign n48913 = n48910 | n48911;
  assign n48914 = ~n48912 & n48913;
  assign n65779 = n48791 & n48914;
  assign n65780 = (n48914 & n65708) | (n48914 & n65779) | (n65708 & n65779);
  assign n65781 = n48791 | n48914;
  assign n65782 = n65708 | n65781;
  assign n48917 = ~n65780 & n65782;
  assign n48918 = x167 & x233;
  assign n48919 = n48917 & n48918;
  assign n48920 = n48917 | n48918;
  assign n48921 = ~n48919 & n48920;
  assign n65783 = n48798 & n48921;
  assign n65784 = (n48921 & n65712) | (n48921 & n65783) | (n65712 & n65783);
  assign n65785 = n48798 | n48921;
  assign n65786 = n65712 | n65785;
  assign n48924 = ~n65784 & n65786;
  assign n48925 = x166 & x234;
  assign n48926 = n48924 & n48925;
  assign n48927 = n48924 | n48925;
  assign n48928 = ~n48926 & n48927;
  assign n65787 = n48805 & n48928;
  assign n65788 = (n48928 & n65716) | (n48928 & n65787) | (n65716 & n65787);
  assign n65789 = n48805 | n48928;
  assign n65790 = n65716 | n65789;
  assign n48931 = ~n65788 & n65790;
  assign n48932 = x165 & x235;
  assign n48933 = n48931 & n48932;
  assign n48934 = n48931 | n48932;
  assign n48935 = ~n48933 & n48934;
  assign n65791 = n48812 & n48935;
  assign n65792 = (n48935 & n65720) | (n48935 & n65791) | (n65720 & n65791);
  assign n65793 = n48812 | n48935;
  assign n65794 = n65720 | n65793;
  assign n48938 = ~n65792 & n65794;
  assign n48939 = x164 & x236;
  assign n48940 = n48938 & n48939;
  assign n48941 = n48938 | n48939;
  assign n48942 = ~n48940 & n48941;
  assign n65795 = n48819 & n48942;
  assign n65796 = (n48942 & n65724) | (n48942 & n65795) | (n65724 & n65795);
  assign n65797 = n48819 | n48942;
  assign n65798 = n65724 | n65797;
  assign n48945 = ~n65796 & n65798;
  assign n48946 = x163 & x237;
  assign n48947 = n48945 & n48946;
  assign n48948 = n48945 | n48946;
  assign n48949 = ~n48947 & n48948;
  assign n65799 = n48826 & n48949;
  assign n65800 = (n48949 & n65728) | (n48949 & n65799) | (n65728 & n65799);
  assign n65801 = n48826 | n48949;
  assign n65802 = n65728 | n65801;
  assign n48952 = ~n65800 & n65802;
  assign n48953 = x162 & x238;
  assign n48954 = n48952 & n48953;
  assign n48955 = n48952 | n48953;
  assign n48956 = ~n48954 & n48955;
  assign n65803 = n48833 & n48956;
  assign n65804 = (n48956 & n65732) | (n48956 & n65803) | (n65732 & n65803);
  assign n65805 = n48833 | n48956;
  assign n65806 = n65732 | n65805;
  assign n48959 = ~n65804 & n65806;
  assign n48960 = x161 & x239;
  assign n48961 = n48959 & n48960;
  assign n48962 = n48959 | n48960;
  assign n48963 = ~n48961 & n48962;
  assign n65807 = n48840 & n48963;
  assign n65808 = (n48963 & n65736) | (n48963 & n65807) | (n65736 & n65807);
  assign n65809 = n48840 | n48963;
  assign n65810 = n65736 | n65809;
  assign n48966 = ~n65808 & n65810;
  assign n65741 = (n74435 & n74461) | (n74435 & n65740) | (n74461 & n65740);
  assign n65814 = n48870 | n48872;
  assign n74493 = n48749 | n48870;
  assign n74494 = (n48870 & n48872) | (n48870 & n74493) | (n48872 & n74493);
  assign n74495 = (n65682 & n65814) | (n65682 & n74494) | (n65814 & n74494);
  assign n74496 = (n65681 & n65814) | (n65681 & n74494) | (n65814 & n74494);
  assign n74497 = (n65592 & n74495) | (n65592 & n74496) | (n74495 & n74496);
  assign n48982 = x175 & x226;
  assign n65816 = n48982 & n74467;
  assign n74498 = (n48982 & n65816) | (n48982 & n74473) | (n65816 & n74473);
  assign n74499 = (n48982 & n65754) | (n48982 & n65816) | (n65754 & n65816);
  assign n74500 = (n74443 & n74498) | (n74443 & n74499) | (n74498 & n74499);
  assign n65818 = n48982 | n74467;
  assign n74501 = n65818 | n74473;
  assign n74502 = n65754 | n65818;
  assign n74503 = (n74443 & n74501) | (n74443 & n74502) | (n74501 & n74502);
  assign n48985 = ~n74500 & n74503;
  assign n48986 = n74497 & n48985;
  assign n48987 = n74497 | n48985;
  assign n48988 = ~n48986 & n48987;
  assign n48989 = x174 & x227;
  assign n48990 = n48988 & n48989;
  assign n48991 = n48988 | n48989;
  assign n48992 = ~n48990 & n48991;
  assign n65811 = n48877 | n48879;
  assign n65820 = n48992 & n65811;
  assign n65821 = n48877 & n48992;
  assign n65822 = (n65741 & n65820) | (n65741 & n65821) | (n65820 & n65821);
  assign n65823 = n48992 | n65811;
  assign n65824 = n48877 | n48992;
  assign n65825 = (n65741 & n65823) | (n65741 & n65824) | (n65823 & n65824);
  assign n48995 = ~n65822 & n65825;
  assign n48996 = x173 & x228;
  assign n48997 = n48995 & n48996;
  assign n48998 = n48995 | n48996;
  assign n48999 = ~n48997 & n48998;
  assign n65826 = n48884 & n48999;
  assign n65827 = (n48999 & n74489) | (n48999 & n65826) | (n74489 & n65826);
  assign n65828 = n48884 | n48999;
  assign n65829 = n74489 | n65828;
  assign n49002 = ~n65827 & n65829;
  assign n49003 = x172 & x229;
  assign n49004 = n49002 & n49003;
  assign n49005 = n49002 | n49003;
  assign n49006 = ~n49004 & n49005;
  assign n65830 = n48891 & n49006;
  assign n65831 = (n49006 & n65768) | (n49006 & n65830) | (n65768 & n65830);
  assign n65832 = n48891 | n49006;
  assign n65833 = n65768 | n65832;
  assign n49009 = ~n65831 & n65833;
  assign n49010 = x171 & x230;
  assign n49011 = n49009 & n49010;
  assign n49012 = n49009 | n49010;
  assign n49013 = ~n49011 & n49012;
  assign n65834 = n48898 & n49013;
  assign n65835 = (n49013 & n65772) | (n49013 & n65834) | (n65772 & n65834);
  assign n65836 = n48898 | n49013;
  assign n65837 = n65772 | n65836;
  assign n49016 = ~n65835 & n65837;
  assign n49017 = x170 & x231;
  assign n49018 = n49016 & n49017;
  assign n49019 = n49016 | n49017;
  assign n49020 = ~n49018 & n49019;
  assign n65838 = n48905 & n49020;
  assign n65839 = (n49020 & n65776) | (n49020 & n65838) | (n65776 & n65838);
  assign n65840 = n48905 | n49020;
  assign n65841 = n65776 | n65840;
  assign n49023 = ~n65839 & n65841;
  assign n49024 = x169 & x232;
  assign n49025 = n49023 & n49024;
  assign n49026 = n49023 | n49024;
  assign n49027 = ~n49025 & n49026;
  assign n65842 = n48912 & n49027;
  assign n65843 = (n49027 & n65780) | (n49027 & n65842) | (n65780 & n65842);
  assign n65844 = n48912 | n49027;
  assign n65845 = n65780 | n65844;
  assign n49030 = ~n65843 & n65845;
  assign n49031 = x168 & x233;
  assign n49032 = n49030 & n49031;
  assign n49033 = n49030 | n49031;
  assign n49034 = ~n49032 & n49033;
  assign n65846 = n48919 & n49034;
  assign n65847 = (n49034 & n65784) | (n49034 & n65846) | (n65784 & n65846);
  assign n65848 = n48919 | n49034;
  assign n65849 = n65784 | n65848;
  assign n49037 = ~n65847 & n65849;
  assign n49038 = x167 & x234;
  assign n49039 = n49037 & n49038;
  assign n49040 = n49037 | n49038;
  assign n49041 = ~n49039 & n49040;
  assign n65850 = n48926 & n49041;
  assign n65851 = (n49041 & n65788) | (n49041 & n65850) | (n65788 & n65850);
  assign n65852 = n48926 | n49041;
  assign n65853 = n65788 | n65852;
  assign n49044 = ~n65851 & n65853;
  assign n49045 = x166 & x235;
  assign n49046 = n49044 & n49045;
  assign n49047 = n49044 | n49045;
  assign n49048 = ~n49046 & n49047;
  assign n65854 = n48933 & n49048;
  assign n65855 = (n49048 & n65792) | (n49048 & n65854) | (n65792 & n65854);
  assign n65856 = n48933 | n49048;
  assign n65857 = n65792 | n65856;
  assign n49051 = ~n65855 & n65857;
  assign n49052 = x165 & x236;
  assign n49053 = n49051 & n49052;
  assign n49054 = n49051 | n49052;
  assign n49055 = ~n49053 & n49054;
  assign n65858 = n48940 & n49055;
  assign n65859 = (n49055 & n65796) | (n49055 & n65858) | (n65796 & n65858);
  assign n65860 = n48940 | n49055;
  assign n65861 = n65796 | n65860;
  assign n49058 = ~n65859 & n65861;
  assign n49059 = x164 & x237;
  assign n49060 = n49058 & n49059;
  assign n49061 = n49058 | n49059;
  assign n49062 = ~n49060 & n49061;
  assign n65862 = n48947 & n49062;
  assign n65863 = (n49062 & n65800) | (n49062 & n65862) | (n65800 & n65862);
  assign n65864 = n48947 | n49062;
  assign n65865 = n65800 | n65864;
  assign n49065 = ~n65863 & n65865;
  assign n49066 = x163 & x238;
  assign n49067 = n49065 & n49066;
  assign n49068 = n49065 | n49066;
  assign n49069 = ~n49067 & n49068;
  assign n65866 = n48954 & n49069;
  assign n65867 = (n49069 & n65804) | (n49069 & n65866) | (n65804 & n65866);
  assign n65868 = n48954 | n49069;
  assign n65869 = n65804 | n65868;
  assign n49072 = ~n65867 & n65869;
  assign n49073 = x162 & x239;
  assign n49074 = n49072 & n49073;
  assign n49075 = n49072 | n49073;
  assign n49076 = ~n49074 & n49075;
  assign n65870 = n48961 & n49076;
  assign n65871 = (n49076 & n65808) | (n49076 & n65870) | (n65808 & n65870);
  assign n65872 = n48961 | n49076;
  assign n65873 = n65808 | n65872;
  assign n49079 = ~n65871 & n65873;
  assign n49094 = x175 & x227;
  assign n74506 = n49094 & n74500;
  assign n74507 = (n48985 & n49094) | (n48985 & n74506) | (n49094 & n74506);
  assign n74508 = n49094 & n74498;
  assign n74509 = n49094 & n74499;
  assign n74510 = (n74443 & n74508) | (n74443 & n74509) | (n74508 & n74509);
  assign n65881 = (n74497 & n74507) | (n74497 & n74510) | (n74507 & n74510);
  assign n74511 = n49094 | n74500;
  assign n74512 = n48985 | n74511;
  assign n74513 = n49094 | n74498;
  assign n74514 = n49094 | n74499;
  assign n74515 = (n74443 & n74513) | (n74443 & n74514) | (n74513 & n74514);
  assign n65884 = (n74497 & n74512) | (n74497 & n74515) | (n74512 & n74515);
  assign n49097 = ~n65881 & n65884;
  assign n65885 = n48990 & n49097;
  assign n74516 = (n49097 & n65821) | (n49097 & n65885) | (n65821 & n65885);
  assign n74517 = (n49097 & n65820) | (n49097 & n65885) | (n65820 & n65885);
  assign n74518 = (n65741 & n74516) | (n65741 & n74517) | (n74516 & n74517);
  assign n65887 = n48990 | n49097;
  assign n74519 = n65821 | n65887;
  assign n74520 = n65820 | n65887;
  assign n74521 = (n65741 & n74519) | (n65741 & n74520) | (n74519 & n74520);
  assign n49100 = ~n74518 & n74521;
  assign n49101 = x174 & x228;
  assign n49102 = n49100 & n49101;
  assign n49103 = n49100 | n49101;
  assign n49104 = ~n49102 & n49103;
  assign n65875 = n48997 | n48999;
  assign n74522 = n49104 & n65875;
  assign n74504 = n48884 | n48997;
  assign n74505 = (n48997 & n48999) | (n48997 & n74504) | (n48999 & n74504);
  assign n74523 = n49104 & n74505;
  assign n74524 = (n74489 & n74522) | (n74489 & n74523) | (n74522 & n74523);
  assign n74525 = n49104 | n65875;
  assign n74526 = n49104 | n74505;
  assign n74527 = (n74489 & n74525) | (n74489 & n74526) | (n74525 & n74526);
  assign n49107 = ~n74524 & n74527;
  assign n49108 = x173 & x229;
  assign n49109 = n49107 & n49108;
  assign n49110 = n49107 | n49108;
  assign n49111 = ~n49109 & n49110;
  assign n65889 = n49004 & n49111;
  assign n74528 = (n49111 & n65830) | (n49111 & n65889) | (n65830 & n65889);
  assign n74529 = (n49006 & n49111) | (n49006 & n65889) | (n49111 & n65889);
  assign n74530 = (n65768 & n74528) | (n65768 & n74529) | (n74528 & n74529);
  assign n65891 = n49004 | n49111;
  assign n74531 = n65830 | n65891;
  assign n74532 = n49006 | n65891;
  assign n74533 = (n65768 & n74531) | (n65768 & n74532) | (n74531 & n74532);
  assign n49114 = ~n74530 & n74533;
  assign n49115 = x172 & x230;
  assign n49116 = n49114 & n49115;
  assign n49117 = n49114 | n49115;
  assign n49118 = ~n49116 & n49117;
  assign n65893 = n49011 & n49118;
  assign n65894 = (n49118 & n65835) | (n49118 & n65893) | (n65835 & n65893);
  assign n65895 = n49011 | n49118;
  assign n65896 = n65835 | n65895;
  assign n49121 = ~n65894 & n65896;
  assign n49122 = x171 & x231;
  assign n49123 = n49121 & n49122;
  assign n49124 = n49121 | n49122;
  assign n49125 = ~n49123 & n49124;
  assign n65897 = n49018 & n49125;
  assign n65898 = (n49125 & n65839) | (n49125 & n65897) | (n65839 & n65897);
  assign n65899 = n49018 | n49125;
  assign n65900 = n65839 | n65899;
  assign n49128 = ~n65898 & n65900;
  assign n49129 = x170 & x232;
  assign n49130 = n49128 & n49129;
  assign n49131 = n49128 | n49129;
  assign n49132 = ~n49130 & n49131;
  assign n65901 = n49025 & n49132;
  assign n65902 = (n49132 & n65843) | (n49132 & n65901) | (n65843 & n65901);
  assign n65903 = n49025 | n49132;
  assign n65904 = n65843 | n65903;
  assign n49135 = ~n65902 & n65904;
  assign n49136 = x169 & x233;
  assign n49137 = n49135 & n49136;
  assign n49138 = n49135 | n49136;
  assign n49139 = ~n49137 & n49138;
  assign n65905 = n49032 & n49139;
  assign n65906 = (n49139 & n65847) | (n49139 & n65905) | (n65847 & n65905);
  assign n65907 = n49032 | n49139;
  assign n65908 = n65847 | n65907;
  assign n49142 = ~n65906 & n65908;
  assign n49143 = x168 & x234;
  assign n49144 = n49142 & n49143;
  assign n49145 = n49142 | n49143;
  assign n49146 = ~n49144 & n49145;
  assign n65909 = n49039 & n49146;
  assign n65910 = (n49146 & n65851) | (n49146 & n65909) | (n65851 & n65909);
  assign n65911 = n49039 | n49146;
  assign n65912 = n65851 | n65911;
  assign n49149 = ~n65910 & n65912;
  assign n49150 = x167 & x235;
  assign n49151 = n49149 & n49150;
  assign n49152 = n49149 | n49150;
  assign n49153 = ~n49151 & n49152;
  assign n65913 = n49046 & n49153;
  assign n65914 = (n49153 & n65855) | (n49153 & n65913) | (n65855 & n65913);
  assign n65915 = n49046 | n49153;
  assign n65916 = n65855 | n65915;
  assign n49156 = ~n65914 & n65916;
  assign n49157 = x166 & x236;
  assign n49158 = n49156 & n49157;
  assign n49159 = n49156 | n49157;
  assign n49160 = ~n49158 & n49159;
  assign n65917 = n49053 & n49160;
  assign n65918 = (n49160 & n65859) | (n49160 & n65917) | (n65859 & n65917);
  assign n65919 = n49053 | n49160;
  assign n65920 = n65859 | n65919;
  assign n49163 = ~n65918 & n65920;
  assign n49164 = x165 & x237;
  assign n49165 = n49163 & n49164;
  assign n49166 = n49163 | n49164;
  assign n49167 = ~n49165 & n49166;
  assign n65921 = n49060 & n49167;
  assign n65922 = (n49167 & n65863) | (n49167 & n65921) | (n65863 & n65921);
  assign n65923 = n49060 | n49167;
  assign n65924 = n65863 | n65923;
  assign n49170 = ~n65922 & n65924;
  assign n49171 = x164 & x238;
  assign n49172 = n49170 & n49171;
  assign n49173 = n49170 | n49171;
  assign n49174 = ~n49172 & n49173;
  assign n65925 = n49067 & n49174;
  assign n65926 = (n49174 & n65867) | (n49174 & n65925) | (n65867 & n65925);
  assign n65927 = n49067 | n49174;
  assign n65928 = n65867 | n65927;
  assign n49177 = ~n65926 & n65928;
  assign n49178 = x163 & x239;
  assign n49179 = n49177 & n49178;
  assign n49180 = n49177 | n49178;
  assign n49181 = ~n49179 & n49180;
  assign n65929 = n49074 & n49181;
  assign n65930 = (n49181 & n65871) | (n49181 & n65929) | (n65871 & n65929);
  assign n65931 = n49074 | n49181;
  assign n65932 = n65871 | n65931;
  assign n49184 = ~n65930 & n65932;
  assign n49198 = x175 & x228;
  assign n65936 = n49097 | n65881;
  assign n74534 = (n48990 & n65881) | (n48990 & n65936) | (n65881 & n65936);
  assign n65938 = n49198 & n74534;
  assign n74535 = n49198 & n65881;
  assign n74536 = (n49097 & n49198) | (n49097 & n74535) | (n49198 & n74535);
  assign n74537 = (n65821 & n65938) | (n65821 & n74536) | (n65938 & n74536);
  assign n74538 = (n65820 & n65938) | (n65820 & n74536) | (n65938 & n74536);
  assign n74539 = (n65741 & n74537) | (n65741 & n74538) | (n74537 & n74538);
  assign n65941 = n49198 | n74534;
  assign n74540 = n49198 | n65881;
  assign n74541 = n49097 | n74540;
  assign n74542 = (n65821 & n65941) | (n65821 & n74541) | (n65941 & n74541);
  assign n74543 = (n65820 & n65941) | (n65820 & n74541) | (n65941 & n74541);
  assign n74544 = (n65741 & n74542) | (n65741 & n74543) | (n74542 & n74543);
  assign n49201 = ~n74539 & n74544;
  assign n65945 = n49102 & n49201;
  assign n74545 = (n49104 & n49201) | (n49104 & n65945) | (n49201 & n65945);
  assign n74546 = (n65875 & n65945) | (n65875 & n74545) | (n65945 & n74545);
  assign n74547 = (n65945 & n74505) | (n65945 & n74545) | (n74505 & n74545);
  assign n74548 = (n74489 & n74546) | (n74489 & n74547) | (n74546 & n74547);
  assign n65948 = n49102 | n49201;
  assign n74549 = n49104 | n65948;
  assign n74550 = (n65875 & n65948) | (n65875 & n74549) | (n65948 & n74549);
  assign n74551 = (n65948 & n74505) | (n65948 & n74549) | (n74505 & n74549);
  assign n74552 = (n74489 & n74550) | (n74489 & n74551) | (n74550 & n74551);
  assign n49204 = ~n74548 & n74552;
  assign n49205 = x174 & x229;
  assign n49206 = n49204 & n49205;
  assign n49207 = n49204 | n49205;
  assign n49208 = ~n49206 & n49207;
  assign n65950 = n49109 & n49208;
  assign n65951 = (n49208 & n74530) | (n49208 & n65950) | (n74530 & n65950);
  assign n65952 = n49109 | n49208;
  assign n65953 = n74530 | n65952;
  assign n49211 = ~n65951 & n65953;
  assign n49212 = x173 & x230;
  assign n49213 = n49211 & n49212;
  assign n49214 = n49211 | n49212;
  assign n49215 = ~n49213 & n49214;
  assign n65954 = n49116 & n49215;
  assign n65955 = (n49215 & n65894) | (n49215 & n65954) | (n65894 & n65954);
  assign n65956 = n49116 | n49215;
  assign n65957 = n65894 | n65956;
  assign n49218 = ~n65955 & n65957;
  assign n49219 = x172 & x231;
  assign n49220 = n49218 & n49219;
  assign n49221 = n49218 | n49219;
  assign n49222 = ~n49220 & n49221;
  assign n65958 = n49123 & n49222;
  assign n65959 = (n49222 & n65898) | (n49222 & n65958) | (n65898 & n65958);
  assign n65960 = n49123 | n49222;
  assign n65961 = n65898 | n65960;
  assign n49225 = ~n65959 & n65961;
  assign n49226 = x171 & x232;
  assign n49227 = n49225 & n49226;
  assign n49228 = n49225 | n49226;
  assign n49229 = ~n49227 & n49228;
  assign n65962 = n49130 & n49229;
  assign n65963 = (n49229 & n65902) | (n49229 & n65962) | (n65902 & n65962);
  assign n65964 = n49130 | n49229;
  assign n65965 = n65902 | n65964;
  assign n49232 = ~n65963 & n65965;
  assign n49233 = x170 & x233;
  assign n49234 = n49232 & n49233;
  assign n49235 = n49232 | n49233;
  assign n49236 = ~n49234 & n49235;
  assign n65966 = n49137 & n49236;
  assign n65967 = (n49236 & n65906) | (n49236 & n65966) | (n65906 & n65966);
  assign n65968 = n49137 | n49236;
  assign n65969 = n65906 | n65968;
  assign n49239 = ~n65967 & n65969;
  assign n49240 = x169 & x234;
  assign n49241 = n49239 & n49240;
  assign n49242 = n49239 | n49240;
  assign n49243 = ~n49241 & n49242;
  assign n65970 = n49144 & n49243;
  assign n65971 = (n49243 & n65910) | (n49243 & n65970) | (n65910 & n65970);
  assign n65972 = n49144 | n49243;
  assign n65973 = n65910 | n65972;
  assign n49246 = ~n65971 & n65973;
  assign n49247 = x168 & x235;
  assign n49248 = n49246 & n49247;
  assign n49249 = n49246 | n49247;
  assign n49250 = ~n49248 & n49249;
  assign n65974 = n49151 & n49250;
  assign n65975 = (n49250 & n65914) | (n49250 & n65974) | (n65914 & n65974);
  assign n65976 = n49151 | n49250;
  assign n65977 = n65914 | n65976;
  assign n49253 = ~n65975 & n65977;
  assign n49254 = x167 & x236;
  assign n49255 = n49253 & n49254;
  assign n49256 = n49253 | n49254;
  assign n49257 = ~n49255 & n49256;
  assign n65978 = n49158 & n49257;
  assign n65979 = (n49257 & n65918) | (n49257 & n65978) | (n65918 & n65978);
  assign n65980 = n49158 | n49257;
  assign n65981 = n65918 | n65980;
  assign n49260 = ~n65979 & n65981;
  assign n49261 = x166 & x237;
  assign n49262 = n49260 & n49261;
  assign n49263 = n49260 | n49261;
  assign n49264 = ~n49262 & n49263;
  assign n65982 = n49165 & n49264;
  assign n65983 = (n49264 & n65922) | (n49264 & n65982) | (n65922 & n65982);
  assign n65984 = n49165 | n49264;
  assign n65985 = n65922 | n65984;
  assign n49267 = ~n65983 & n65985;
  assign n49268 = x165 & x238;
  assign n49269 = n49267 & n49268;
  assign n49270 = n49267 | n49268;
  assign n49271 = ~n49269 & n49270;
  assign n65986 = n49172 & n49271;
  assign n65987 = (n49271 & n65926) | (n49271 & n65986) | (n65926 & n65986);
  assign n65988 = n49172 | n49271;
  assign n65989 = n65926 | n65988;
  assign n49274 = ~n65987 & n65989;
  assign n49275 = x164 & x239;
  assign n49276 = n49274 & n49275;
  assign n49277 = n49274 | n49275;
  assign n49278 = ~n49276 & n49277;
  assign n65990 = n49179 & n49278;
  assign n65991 = (n49278 & n65930) | (n49278 & n65990) | (n65930 & n65990);
  assign n65992 = n49179 | n49278;
  assign n65993 = n65930 | n65992;
  assign n49281 = ~n65991 & n65993;
  assign n49294 = x175 & x229;
  assign n65997 = n49294 & n74539;
  assign n65998 = (n49294 & n74548) | (n49294 & n65997) | (n74548 & n65997);
  assign n65999 = n49294 | n74539;
  assign n66000 = n74548 | n65999;
  assign n49297 = ~n65998 & n66000;
  assign n65995 = n49206 | n49208;
  assign n74555 = n49297 & n65995;
  assign n74553 = n49109 | n49206;
  assign n74554 = (n49206 & n49208) | (n49206 & n74553) | (n49208 & n74553);
  assign n74556 = n49297 & n74554;
  assign n74557 = (n74530 & n74555) | (n74530 & n74556) | (n74555 & n74556);
  assign n74558 = n49297 | n65995;
  assign n74559 = n49297 | n74554;
  assign n74560 = (n74530 & n74558) | (n74530 & n74559) | (n74558 & n74559);
  assign n49300 = ~n74557 & n74560;
  assign n49301 = x174 & x230;
  assign n49302 = n49300 & n49301;
  assign n49303 = n49300 | n49301;
  assign n49304 = ~n49302 & n49303;
  assign n66001 = n49213 & n49304;
  assign n74561 = (n49304 & n65954) | (n49304 & n66001) | (n65954 & n66001);
  assign n74562 = (n49215 & n49304) | (n49215 & n66001) | (n49304 & n66001);
  assign n74563 = (n65894 & n74561) | (n65894 & n74562) | (n74561 & n74562);
  assign n66003 = n49213 | n49304;
  assign n74564 = n65954 | n66003;
  assign n74565 = n49215 | n66003;
  assign n74566 = (n65894 & n74564) | (n65894 & n74565) | (n74564 & n74565);
  assign n49307 = ~n74563 & n74566;
  assign n49308 = x173 & x231;
  assign n49309 = n49307 & n49308;
  assign n49310 = n49307 | n49308;
  assign n49311 = ~n49309 & n49310;
  assign n66005 = n49220 & n49311;
  assign n66006 = (n49311 & n65959) | (n49311 & n66005) | (n65959 & n66005);
  assign n66007 = n49220 | n49311;
  assign n66008 = n65959 | n66007;
  assign n49314 = ~n66006 & n66008;
  assign n49315 = x172 & x232;
  assign n49316 = n49314 & n49315;
  assign n49317 = n49314 | n49315;
  assign n49318 = ~n49316 & n49317;
  assign n66009 = n49227 & n49318;
  assign n66010 = (n49318 & n65963) | (n49318 & n66009) | (n65963 & n66009);
  assign n66011 = n49227 | n49318;
  assign n66012 = n65963 | n66011;
  assign n49321 = ~n66010 & n66012;
  assign n49322 = x171 & x233;
  assign n49323 = n49321 & n49322;
  assign n49324 = n49321 | n49322;
  assign n49325 = ~n49323 & n49324;
  assign n66013 = n49234 & n49325;
  assign n66014 = (n49325 & n65967) | (n49325 & n66013) | (n65967 & n66013);
  assign n66015 = n49234 | n49325;
  assign n66016 = n65967 | n66015;
  assign n49328 = ~n66014 & n66016;
  assign n49329 = x170 & x234;
  assign n49330 = n49328 & n49329;
  assign n49331 = n49328 | n49329;
  assign n49332 = ~n49330 & n49331;
  assign n66017 = n49241 & n49332;
  assign n66018 = (n49332 & n65971) | (n49332 & n66017) | (n65971 & n66017);
  assign n66019 = n49241 | n49332;
  assign n66020 = n65971 | n66019;
  assign n49335 = ~n66018 & n66020;
  assign n49336 = x169 & x235;
  assign n49337 = n49335 & n49336;
  assign n49338 = n49335 | n49336;
  assign n49339 = ~n49337 & n49338;
  assign n66021 = n49248 & n49339;
  assign n66022 = (n49339 & n65975) | (n49339 & n66021) | (n65975 & n66021);
  assign n66023 = n49248 | n49339;
  assign n66024 = n65975 | n66023;
  assign n49342 = ~n66022 & n66024;
  assign n49343 = x168 & x236;
  assign n49344 = n49342 & n49343;
  assign n49345 = n49342 | n49343;
  assign n49346 = ~n49344 & n49345;
  assign n66025 = n49255 & n49346;
  assign n66026 = (n49346 & n65979) | (n49346 & n66025) | (n65979 & n66025);
  assign n66027 = n49255 | n49346;
  assign n66028 = n65979 | n66027;
  assign n49349 = ~n66026 & n66028;
  assign n49350 = x167 & x237;
  assign n49351 = n49349 & n49350;
  assign n49352 = n49349 | n49350;
  assign n49353 = ~n49351 & n49352;
  assign n66029 = n49262 & n49353;
  assign n66030 = (n49353 & n65983) | (n49353 & n66029) | (n65983 & n66029);
  assign n66031 = n49262 | n49353;
  assign n66032 = n65983 | n66031;
  assign n49356 = ~n66030 & n66032;
  assign n49357 = x166 & x238;
  assign n49358 = n49356 & n49357;
  assign n49359 = n49356 | n49357;
  assign n49360 = ~n49358 & n49359;
  assign n66033 = n49269 & n49360;
  assign n66034 = (n49360 & n65987) | (n49360 & n66033) | (n65987 & n66033);
  assign n66035 = n49269 | n49360;
  assign n66036 = n65987 | n66035;
  assign n49363 = ~n66034 & n66036;
  assign n49364 = x165 & x239;
  assign n49365 = n49363 & n49364;
  assign n49366 = n49363 | n49364;
  assign n49367 = ~n49365 & n49366;
  assign n66037 = n49276 & n49367;
  assign n66038 = (n49367 & n65991) | (n49367 & n66037) | (n65991 & n66037);
  assign n66039 = n49276 | n49367;
  assign n66040 = n65991 | n66039;
  assign n49370 = ~n66038 & n66040;
  assign n49382 = x175 & x230;
  assign n74568 = n49382 & n65997;
  assign n74569 = n49294 & n49382;
  assign n74570 = (n74548 & n74568) | (n74548 & n74569) | (n74568 & n74569);
  assign n74567 = (n49297 & n49382) | (n49297 & n74570) | (n49382 & n74570);
  assign n74571 = (n65995 & n74567) | (n65995 & n74570) | (n74567 & n74570);
  assign n74572 = (n74554 & n74567) | (n74554 & n74570) | (n74567 & n74570);
  assign n74573 = (n74530 & n74571) | (n74530 & n74572) | (n74571 & n74572);
  assign n74575 = n49382 | n65997;
  assign n74576 = n49294 | n49382;
  assign n74577 = (n74548 & n74575) | (n74548 & n74576) | (n74575 & n74576);
  assign n74574 = n49297 | n74577;
  assign n74578 = (n65995 & n74574) | (n65995 & n74577) | (n74574 & n74577);
  assign n74579 = (n74554 & n74574) | (n74554 & n74577) | (n74574 & n74577);
  assign n74580 = (n74530 & n74578) | (n74530 & n74579) | (n74578 & n74579);
  assign n49385 = ~n74573 & n74580;
  assign n66049 = n49302 & n49385;
  assign n66050 = (n49385 & n74563) | (n49385 & n66049) | (n74563 & n66049);
  assign n66051 = n49302 | n49385;
  assign n66052 = n74563 | n66051;
  assign n49388 = ~n66050 & n66052;
  assign n49389 = x174 & x231;
  assign n49390 = n49388 & n49389;
  assign n49391 = n49388 | n49389;
  assign n49392 = ~n49390 & n49391;
  assign n66053 = n49309 & n49392;
  assign n66054 = (n49392 & n66006) | (n49392 & n66053) | (n66006 & n66053);
  assign n66055 = n49309 | n49392;
  assign n66056 = n66006 | n66055;
  assign n49395 = ~n66054 & n66056;
  assign n49396 = x173 & x232;
  assign n49397 = n49395 & n49396;
  assign n49398 = n49395 | n49396;
  assign n49399 = ~n49397 & n49398;
  assign n66057 = n49316 & n49399;
  assign n66058 = (n49399 & n66010) | (n49399 & n66057) | (n66010 & n66057);
  assign n66059 = n49316 | n49399;
  assign n66060 = n66010 | n66059;
  assign n49402 = ~n66058 & n66060;
  assign n49403 = x172 & x233;
  assign n49404 = n49402 & n49403;
  assign n49405 = n49402 | n49403;
  assign n49406 = ~n49404 & n49405;
  assign n66061 = n49323 & n49406;
  assign n66062 = (n49406 & n66014) | (n49406 & n66061) | (n66014 & n66061);
  assign n66063 = n49323 | n49406;
  assign n66064 = n66014 | n66063;
  assign n49409 = ~n66062 & n66064;
  assign n49410 = x171 & x234;
  assign n49411 = n49409 & n49410;
  assign n49412 = n49409 | n49410;
  assign n49413 = ~n49411 & n49412;
  assign n66065 = n49330 & n49413;
  assign n66066 = (n49413 & n66018) | (n49413 & n66065) | (n66018 & n66065);
  assign n66067 = n49330 | n49413;
  assign n66068 = n66018 | n66067;
  assign n49416 = ~n66066 & n66068;
  assign n49417 = x170 & x235;
  assign n49418 = n49416 & n49417;
  assign n49419 = n49416 | n49417;
  assign n49420 = ~n49418 & n49419;
  assign n66069 = n49337 & n49420;
  assign n66070 = (n49420 & n66022) | (n49420 & n66069) | (n66022 & n66069);
  assign n66071 = n49337 | n49420;
  assign n66072 = n66022 | n66071;
  assign n49423 = ~n66070 & n66072;
  assign n49424 = x169 & x236;
  assign n49425 = n49423 & n49424;
  assign n49426 = n49423 | n49424;
  assign n49427 = ~n49425 & n49426;
  assign n66073 = n49344 & n49427;
  assign n66074 = (n49427 & n66026) | (n49427 & n66073) | (n66026 & n66073);
  assign n66075 = n49344 | n49427;
  assign n66076 = n66026 | n66075;
  assign n49430 = ~n66074 & n66076;
  assign n49431 = x168 & x237;
  assign n49432 = n49430 & n49431;
  assign n49433 = n49430 | n49431;
  assign n49434 = ~n49432 & n49433;
  assign n66077 = n49351 & n49434;
  assign n66078 = (n49434 & n66030) | (n49434 & n66077) | (n66030 & n66077);
  assign n66079 = n49351 | n49434;
  assign n66080 = n66030 | n66079;
  assign n49437 = ~n66078 & n66080;
  assign n49438 = x167 & x238;
  assign n49439 = n49437 & n49438;
  assign n49440 = n49437 | n49438;
  assign n49441 = ~n49439 & n49440;
  assign n66081 = n49358 & n49441;
  assign n66082 = (n49441 & n66034) | (n49441 & n66081) | (n66034 & n66081);
  assign n66083 = n49358 | n49441;
  assign n66084 = n66034 | n66083;
  assign n49444 = ~n66082 & n66084;
  assign n49445 = x166 & x239;
  assign n49446 = n49444 & n49445;
  assign n49447 = n49444 | n49445;
  assign n49448 = ~n49446 & n49447;
  assign n66085 = n49365 & n49448;
  assign n66086 = (n49448 & n66038) | (n49448 & n66085) | (n66038 & n66085);
  assign n66087 = n49365 | n49448;
  assign n66088 = n66038 | n66087;
  assign n49451 = ~n66086 & n66088;
  assign n49462 = x175 & x231;
  assign n74581 = n49385 | n74573;
  assign n74582 = (n49302 & n74573) | (n49302 & n74581) | (n74573 & n74581);
  assign n66092 = n49462 & n74582;
  assign n74583 = n49462 & n74573;
  assign n74584 = (n49385 & n49462) | (n49385 & n74583) | (n49462 & n74583);
  assign n66094 = (n74563 & n66092) | (n74563 & n74584) | (n66092 & n74584);
  assign n66095 = n49462 | n74582;
  assign n74585 = n49462 | n74573;
  assign n74586 = n49385 | n74585;
  assign n66097 = (n74563 & n66095) | (n74563 & n74586) | (n66095 & n74586);
  assign n49465 = ~n66094 & n66097;
  assign n66098 = n49390 & n49465;
  assign n74587 = (n49465 & n66053) | (n49465 & n66098) | (n66053 & n66098);
  assign n74588 = (n49392 & n49465) | (n49392 & n66098) | (n49465 & n66098);
  assign n74589 = (n66006 & n74587) | (n66006 & n74588) | (n74587 & n74588);
  assign n66100 = n49390 | n49465;
  assign n74590 = n66053 | n66100;
  assign n74591 = n49392 | n66100;
  assign n74592 = (n66006 & n74590) | (n66006 & n74591) | (n74590 & n74591);
  assign n49468 = ~n74589 & n74592;
  assign n49469 = x174 & x232;
  assign n49470 = n49468 & n49469;
  assign n49471 = n49468 | n49469;
  assign n49472 = ~n49470 & n49471;
  assign n66102 = n49397 & n49472;
  assign n66103 = (n49472 & n66058) | (n49472 & n66102) | (n66058 & n66102);
  assign n66104 = n49397 | n49472;
  assign n66105 = n66058 | n66104;
  assign n49475 = ~n66103 & n66105;
  assign n49476 = x173 & x233;
  assign n49477 = n49475 & n49476;
  assign n49478 = n49475 | n49476;
  assign n49479 = ~n49477 & n49478;
  assign n66106 = n49404 & n49479;
  assign n66107 = (n49479 & n66062) | (n49479 & n66106) | (n66062 & n66106);
  assign n66108 = n49404 | n49479;
  assign n66109 = n66062 | n66108;
  assign n49482 = ~n66107 & n66109;
  assign n49483 = x172 & x234;
  assign n49484 = n49482 & n49483;
  assign n49485 = n49482 | n49483;
  assign n49486 = ~n49484 & n49485;
  assign n66110 = n49411 & n49486;
  assign n66111 = (n49486 & n66066) | (n49486 & n66110) | (n66066 & n66110);
  assign n66112 = n49411 | n49486;
  assign n66113 = n66066 | n66112;
  assign n49489 = ~n66111 & n66113;
  assign n49490 = x171 & x235;
  assign n49491 = n49489 & n49490;
  assign n49492 = n49489 | n49490;
  assign n49493 = ~n49491 & n49492;
  assign n66114 = n49418 & n49493;
  assign n66115 = (n49493 & n66070) | (n49493 & n66114) | (n66070 & n66114);
  assign n66116 = n49418 | n49493;
  assign n66117 = n66070 | n66116;
  assign n49496 = ~n66115 & n66117;
  assign n49497 = x170 & x236;
  assign n49498 = n49496 & n49497;
  assign n49499 = n49496 | n49497;
  assign n49500 = ~n49498 & n49499;
  assign n66118 = n49425 & n49500;
  assign n66119 = (n49500 & n66074) | (n49500 & n66118) | (n66074 & n66118);
  assign n66120 = n49425 | n49500;
  assign n66121 = n66074 | n66120;
  assign n49503 = ~n66119 & n66121;
  assign n49504 = x169 & x237;
  assign n49505 = n49503 & n49504;
  assign n49506 = n49503 | n49504;
  assign n49507 = ~n49505 & n49506;
  assign n66122 = n49432 & n49507;
  assign n66123 = (n49507 & n66078) | (n49507 & n66122) | (n66078 & n66122);
  assign n66124 = n49432 | n49507;
  assign n66125 = n66078 | n66124;
  assign n49510 = ~n66123 & n66125;
  assign n49511 = x168 & x238;
  assign n49512 = n49510 & n49511;
  assign n49513 = n49510 | n49511;
  assign n49514 = ~n49512 & n49513;
  assign n66126 = n49439 & n49514;
  assign n66127 = (n49514 & n66082) | (n49514 & n66126) | (n66082 & n66126);
  assign n66128 = n49439 | n49514;
  assign n66129 = n66082 | n66128;
  assign n49517 = ~n66127 & n66129;
  assign n49518 = x167 & x239;
  assign n49519 = n49517 & n49518;
  assign n49520 = n49517 | n49518;
  assign n49521 = ~n49519 & n49520;
  assign n66130 = n49446 & n49521;
  assign n66131 = (n49521 & n66086) | (n49521 & n66130) | (n66086 & n66130);
  assign n66132 = n49446 | n49521;
  assign n66133 = n66086 | n66132;
  assign n49524 = ~n66131 & n66133;
  assign n49534 = x175 & x232;
  assign n66135 = n49465 | n66094;
  assign n74593 = (n49390 & n66094) | (n49390 & n66135) | (n66094 & n66135);
  assign n66137 = n49534 & n74593;
  assign n74594 = n49534 & n66094;
  assign n74595 = (n49465 & n49534) | (n49465 & n74594) | (n49534 & n74594);
  assign n74596 = (n66053 & n66137) | (n66053 & n74595) | (n66137 & n74595);
  assign n74597 = (n49392 & n66137) | (n49392 & n74595) | (n66137 & n74595);
  assign n74598 = (n66006 & n74596) | (n66006 & n74597) | (n74596 & n74597);
  assign n66140 = n49534 | n74593;
  assign n74599 = n49534 | n66094;
  assign n74600 = n49465 | n74599;
  assign n74601 = (n66053 & n66140) | (n66053 & n74600) | (n66140 & n74600);
  assign n74602 = (n49392 & n66140) | (n49392 & n74600) | (n66140 & n74600);
  assign n74603 = (n66006 & n74601) | (n66006 & n74602) | (n74601 & n74602);
  assign n49537 = ~n74598 & n74603;
  assign n66143 = n49470 & n49537;
  assign n74604 = (n49537 & n66102) | (n49537 & n66143) | (n66102 & n66143);
  assign n74605 = (n49472 & n49537) | (n49472 & n66143) | (n49537 & n66143);
  assign n74606 = (n66058 & n74604) | (n66058 & n74605) | (n74604 & n74605);
  assign n66145 = n49470 | n49537;
  assign n74607 = n66102 | n66145;
  assign n74608 = n49472 | n66145;
  assign n74609 = (n66058 & n74607) | (n66058 & n74608) | (n74607 & n74608);
  assign n49540 = ~n74606 & n74609;
  assign n49541 = x174 & x233;
  assign n49542 = n49540 & n49541;
  assign n49543 = n49540 | n49541;
  assign n49544 = ~n49542 & n49543;
  assign n66147 = n49477 & n49544;
  assign n66148 = (n49544 & n66107) | (n49544 & n66147) | (n66107 & n66147);
  assign n66149 = n49477 | n49544;
  assign n66150 = n66107 | n66149;
  assign n49547 = ~n66148 & n66150;
  assign n49548 = x173 & x234;
  assign n49549 = n49547 & n49548;
  assign n49550 = n49547 | n49548;
  assign n49551 = ~n49549 & n49550;
  assign n66151 = n49484 & n49551;
  assign n66152 = (n49551 & n66111) | (n49551 & n66151) | (n66111 & n66151);
  assign n66153 = n49484 | n49551;
  assign n66154 = n66111 | n66153;
  assign n49554 = ~n66152 & n66154;
  assign n49555 = x172 & x235;
  assign n49556 = n49554 & n49555;
  assign n49557 = n49554 | n49555;
  assign n49558 = ~n49556 & n49557;
  assign n66155 = n49491 & n49558;
  assign n66156 = (n49558 & n66115) | (n49558 & n66155) | (n66115 & n66155);
  assign n66157 = n49491 | n49558;
  assign n66158 = n66115 | n66157;
  assign n49561 = ~n66156 & n66158;
  assign n49562 = x171 & x236;
  assign n49563 = n49561 & n49562;
  assign n49564 = n49561 | n49562;
  assign n49565 = ~n49563 & n49564;
  assign n66159 = n49498 & n49565;
  assign n66160 = (n49565 & n66119) | (n49565 & n66159) | (n66119 & n66159);
  assign n66161 = n49498 | n49565;
  assign n66162 = n66119 | n66161;
  assign n49568 = ~n66160 & n66162;
  assign n49569 = x170 & x237;
  assign n49570 = n49568 & n49569;
  assign n49571 = n49568 | n49569;
  assign n49572 = ~n49570 & n49571;
  assign n66163 = n49505 & n49572;
  assign n66164 = (n49572 & n66123) | (n49572 & n66163) | (n66123 & n66163);
  assign n66165 = n49505 | n49572;
  assign n66166 = n66123 | n66165;
  assign n49575 = ~n66164 & n66166;
  assign n49576 = x169 & x238;
  assign n49577 = n49575 & n49576;
  assign n49578 = n49575 | n49576;
  assign n49579 = ~n49577 & n49578;
  assign n66167 = n49512 & n49579;
  assign n66168 = (n49579 & n66127) | (n49579 & n66167) | (n66127 & n66167);
  assign n66169 = n49512 | n49579;
  assign n66170 = n66127 | n66169;
  assign n49582 = ~n66168 & n66170;
  assign n49583 = x168 & x239;
  assign n49584 = n49582 & n49583;
  assign n49585 = n49582 | n49583;
  assign n49586 = ~n49584 & n49585;
  assign n66171 = n49519 & n49586;
  assign n66172 = (n49586 & n66131) | (n49586 & n66171) | (n66131 & n66171);
  assign n66173 = n49519 | n49586;
  assign n66174 = n66131 | n66173;
  assign n49589 = ~n66172 & n66174;
  assign n49598 = x175 & x233;
  assign n74610 = n49537 | n74598;
  assign n74611 = (n49470 & n74598) | (n49470 & n74610) | (n74598 & n74610);
  assign n66178 = n49598 & n74611;
  assign n74612 = n49598 & n74598;
  assign n74613 = (n49537 & n49598) | (n49537 & n74612) | (n49598 & n74612);
  assign n74614 = (n66102 & n66178) | (n66102 & n74613) | (n66178 & n74613);
  assign n74615 = (n49472 & n66178) | (n49472 & n74613) | (n66178 & n74613);
  assign n74616 = (n66058 & n74614) | (n66058 & n74615) | (n74614 & n74615);
  assign n66181 = n49598 | n74611;
  assign n74617 = n49598 | n74598;
  assign n74618 = n49537 | n74617;
  assign n74619 = (n66102 & n66181) | (n66102 & n74618) | (n66181 & n74618);
  assign n74620 = (n49472 & n66181) | (n49472 & n74618) | (n66181 & n74618);
  assign n74621 = (n66058 & n74619) | (n66058 & n74620) | (n74619 & n74620);
  assign n49601 = ~n74616 & n74621;
  assign n66184 = n49542 & n49601;
  assign n74622 = (n49601 & n66147) | (n49601 & n66184) | (n66147 & n66184);
  assign n74623 = (n49544 & n49601) | (n49544 & n66184) | (n49601 & n66184);
  assign n74624 = (n66107 & n74622) | (n66107 & n74623) | (n74622 & n74623);
  assign n66186 = n49542 | n49601;
  assign n74625 = n66147 | n66186;
  assign n74626 = n49544 | n66186;
  assign n74627 = (n66107 & n74625) | (n66107 & n74626) | (n74625 & n74626);
  assign n49604 = ~n74624 & n74627;
  assign n49605 = x174 & x234;
  assign n49606 = n49604 & n49605;
  assign n49607 = n49604 | n49605;
  assign n49608 = ~n49606 & n49607;
  assign n66188 = n49549 & n49608;
  assign n66189 = (n49608 & n66152) | (n49608 & n66188) | (n66152 & n66188);
  assign n66190 = n49549 | n49608;
  assign n66191 = n66152 | n66190;
  assign n49611 = ~n66189 & n66191;
  assign n49612 = x173 & x235;
  assign n49613 = n49611 & n49612;
  assign n49614 = n49611 | n49612;
  assign n49615 = ~n49613 & n49614;
  assign n66192 = n49556 & n49615;
  assign n66193 = (n49615 & n66156) | (n49615 & n66192) | (n66156 & n66192);
  assign n66194 = n49556 | n49615;
  assign n66195 = n66156 | n66194;
  assign n49618 = ~n66193 & n66195;
  assign n49619 = x172 & x236;
  assign n49620 = n49618 & n49619;
  assign n49621 = n49618 | n49619;
  assign n49622 = ~n49620 & n49621;
  assign n66196 = n49563 & n49622;
  assign n66197 = (n49622 & n66160) | (n49622 & n66196) | (n66160 & n66196);
  assign n66198 = n49563 | n49622;
  assign n66199 = n66160 | n66198;
  assign n49625 = ~n66197 & n66199;
  assign n49626 = x171 & x237;
  assign n49627 = n49625 & n49626;
  assign n49628 = n49625 | n49626;
  assign n49629 = ~n49627 & n49628;
  assign n66200 = n49570 & n49629;
  assign n66201 = (n49629 & n66164) | (n49629 & n66200) | (n66164 & n66200);
  assign n66202 = n49570 | n49629;
  assign n66203 = n66164 | n66202;
  assign n49632 = ~n66201 & n66203;
  assign n49633 = x170 & x238;
  assign n49634 = n49632 & n49633;
  assign n49635 = n49632 | n49633;
  assign n49636 = ~n49634 & n49635;
  assign n66204 = n49577 & n49636;
  assign n66205 = (n49636 & n66168) | (n49636 & n66204) | (n66168 & n66204);
  assign n66206 = n49577 | n49636;
  assign n66207 = n66168 | n66206;
  assign n49639 = ~n66205 & n66207;
  assign n49640 = x169 & x239;
  assign n49641 = n49639 & n49640;
  assign n49642 = n49639 | n49640;
  assign n49643 = ~n49641 & n49642;
  assign n66208 = n49584 & n49643;
  assign n66209 = (n49643 & n66172) | (n49643 & n66208) | (n66172 & n66208);
  assign n66210 = n49584 | n49643;
  assign n66211 = n66172 | n66210;
  assign n49646 = ~n66209 & n66211;
  assign n49654 = x175 & x234;
  assign n74628 = n49601 | n74616;
  assign n74629 = (n49542 & n74616) | (n49542 & n74628) | (n74616 & n74628);
  assign n66215 = n49654 & n74629;
  assign n74630 = n49654 & n74616;
  assign n74631 = (n49601 & n49654) | (n49601 & n74630) | (n49654 & n74630);
  assign n74632 = (n66147 & n66215) | (n66147 & n74631) | (n66215 & n74631);
  assign n74633 = (n49544 & n66215) | (n49544 & n74631) | (n66215 & n74631);
  assign n74634 = (n66107 & n74632) | (n66107 & n74633) | (n74632 & n74633);
  assign n66218 = n49654 | n74629;
  assign n74635 = n49654 | n74616;
  assign n74636 = n49601 | n74635;
  assign n74637 = (n66147 & n66218) | (n66147 & n74636) | (n66218 & n74636);
  assign n74638 = (n49544 & n66218) | (n49544 & n74636) | (n66218 & n74636);
  assign n74639 = (n66107 & n74637) | (n66107 & n74638) | (n74637 & n74638);
  assign n49657 = ~n74634 & n74639;
  assign n66221 = n49606 & n49657;
  assign n74640 = (n49657 & n66188) | (n49657 & n66221) | (n66188 & n66221);
  assign n74641 = (n49608 & n49657) | (n49608 & n66221) | (n49657 & n66221);
  assign n74642 = (n66152 & n74640) | (n66152 & n74641) | (n74640 & n74641);
  assign n66223 = n49606 | n49657;
  assign n74643 = n66188 | n66223;
  assign n74644 = n49608 | n66223;
  assign n74645 = (n66152 & n74643) | (n66152 & n74644) | (n74643 & n74644);
  assign n49660 = ~n74642 & n74645;
  assign n49661 = x174 & x235;
  assign n49662 = n49660 & n49661;
  assign n49663 = n49660 | n49661;
  assign n49664 = ~n49662 & n49663;
  assign n66225 = n49613 & n49664;
  assign n66226 = (n49664 & n66193) | (n49664 & n66225) | (n66193 & n66225);
  assign n66227 = n49613 | n49664;
  assign n66228 = n66193 | n66227;
  assign n49667 = ~n66226 & n66228;
  assign n49668 = x173 & x236;
  assign n49669 = n49667 & n49668;
  assign n49670 = n49667 | n49668;
  assign n49671 = ~n49669 & n49670;
  assign n66229 = n49620 & n49671;
  assign n66230 = (n49671 & n66197) | (n49671 & n66229) | (n66197 & n66229);
  assign n66231 = n49620 | n49671;
  assign n66232 = n66197 | n66231;
  assign n49674 = ~n66230 & n66232;
  assign n49675 = x172 & x237;
  assign n49676 = n49674 & n49675;
  assign n49677 = n49674 | n49675;
  assign n49678 = ~n49676 & n49677;
  assign n66233 = n49627 & n49678;
  assign n66234 = (n49678 & n66201) | (n49678 & n66233) | (n66201 & n66233);
  assign n66235 = n49627 | n49678;
  assign n66236 = n66201 | n66235;
  assign n49681 = ~n66234 & n66236;
  assign n49682 = x171 & x238;
  assign n49683 = n49681 & n49682;
  assign n49684 = n49681 | n49682;
  assign n49685 = ~n49683 & n49684;
  assign n66237 = n49634 & n49685;
  assign n66238 = (n49685 & n66205) | (n49685 & n66237) | (n66205 & n66237);
  assign n66239 = n49634 | n49685;
  assign n66240 = n66205 | n66239;
  assign n49688 = ~n66238 & n66240;
  assign n49689 = x170 & x239;
  assign n49690 = n49688 & n49689;
  assign n49691 = n49688 | n49689;
  assign n49692 = ~n49690 & n49691;
  assign n66241 = n49641 & n49692;
  assign n66242 = (n49692 & n66209) | (n49692 & n66241) | (n66209 & n66241);
  assign n66243 = n49641 | n49692;
  assign n66244 = n66209 | n66243;
  assign n49695 = ~n66242 & n66244;
  assign n49702 = x175 & x235;
  assign n74646 = n49657 | n74634;
  assign n74647 = (n49606 & n74634) | (n49606 & n74646) | (n74634 & n74646);
  assign n66248 = n49702 & n74647;
  assign n74648 = n49702 & n74634;
  assign n74649 = (n49657 & n49702) | (n49657 & n74648) | (n49702 & n74648);
  assign n74650 = (n66188 & n66248) | (n66188 & n74649) | (n66248 & n74649);
  assign n74651 = (n49608 & n66248) | (n49608 & n74649) | (n66248 & n74649);
  assign n74652 = (n66152 & n74650) | (n66152 & n74651) | (n74650 & n74651);
  assign n66251 = n49702 | n74647;
  assign n74653 = n49702 | n74634;
  assign n74654 = n49657 | n74653;
  assign n74655 = (n66188 & n66251) | (n66188 & n74654) | (n66251 & n74654);
  assign n74656 = (n49608 & n66251) | (n49608 & n74654) | (n66251 & n74654);
  assign n74657 = (n66152 & n74655) | (n66152 & n74656) | (n74655 & n74656);
  assign n49705 = ~n74652 & n74657;
  assign n66254 = n49662 & n49705;
  assign n74658 = (n49705 & n66225) | (n49705 & n66254) | (n66225 & n66254);
  assign n74659 = (n49664 & n49705) | (n49664 & n66254) | (n49705 & n66254);
  assign n74660 = (n66193 & n74658) | (n66193 & n74659) | (n74658 & n74659);
  assign n66256 = n49662 | n49705;
  assign n74661 = n66225 | n66256;
  assign n74662 = n49664 | n66256;
  assign n74663 = (n66193 & n74661) | (n66193 & n74662) | (n74661 & n74662);
  assign n49708 = ~n74660 & n74663;
  assign n49709 = x174 & x236;
  assign n49710 = n49708 & n49709;
  assign n49711 = n49708 | n49709;
  assign n49712 = ~n49710 & n49711;
  assign n66258 = n49669 & n49712;
  assign n66259 = (n49712 & n66230) | (n49712 & n66258) | (n66230 & n66258);
  assign n66260 = n49669 | n49712;
  assign n66261 = n66230 | n66260;
  assign n49715 = ~n66259 & n66261;
  assign n49716 = x173 & x237;
  assign n49717 = n49715 & n49716;
  assign n49718 = n49715 | n49716;
  assign n49719 = ~n49717 & n49718;
  assign n66262 = n49676 & n49719;
  assign n66263 = (n49719 & n66234) | (n49719 & n66262) | (n66234 & n66262);
  assign n66264 = n49676 | n49719;
  assign n66265 = n66234 | n66264;
  assign n49722 = ~n66263 & n66265;
  assign n49723 = x172 & x238;
  assign n49724 = n49722 & n49723;
  assign n49725 = n49722 | n49723;
  assign n49726 = ~n49724 & n49725;
  assign n66266 = n49683 & n49726;
  assign n66267 = (n49726 & n66238) | (n49726 & n66266) | (n66238 & n66266);
  assign n66268 = n49683 | n49726;
  assign n66269 = n66238 | n66268;
  assign n49729 = ~n66267 & n66269;
  assign n49730 = x171 & x239;
  assign n49731 = n49729 & n49730;
  assign n49732 = n49729 | n49730;
  assign n49733 = ~n49731 & n49732;
  assign n66270 = n49690 & n49733;
  assign n66271 = (n49733 & n66242) | (n49733 & n66270) | (n66242 & n66270);
  assign n66272 = n49690 | n49733;
  assign n66273 = n66242 | n66272;
  assign n49736 = ~n66271 & n66273;
  assign n49742 = x175 & x236;
  assign n74664 = n49705 | n74652;
  assign n74665 = (n49662 & n74652) | (n49662 & n74664) | (n74652 & n74664);
  assign n66277 = n49742 & n74665;
  assign n74666 = n49742 & n74652;
  assign n74667 = (n49705 & n49742) | (n49705 & n74666) | (n49742 & n74666);
  assign n74668 = (n66225 & n66277) | (n66225 & n74667) | (n66277 & n74667);
  assign n74669 = (n49664 & n66277) | (n49664 & n74667) | (n66277 & n74667);
  assign n74670 = (n66193 & n74668) | (n66193 & n74669) | (n74668 & n74669);
  assign n66280 = n49742 | n74665;
  assign n74671 = n49742 | n74652;
  assign n74672 = n49705 | n74671;
  assign n74673 = (n66225 & n66280) | (n66225 & n74672) | (n66280 & n74672);
  assign n74674 = (n49664 & n66280) | (n49664 & n74672) | (n66280 & n74672);
  assign n74675 = (n66193 & n74673) | (n66193 & n74674) | (n74673 & n74674);
  assign n49745 = ~n74670 & n74675;
  assign n66283 = n49710 & n49745;
  assign n74676 = (n49745 & n66258) | (n49745 & n66283) | (n66258 & n66283);
  assign n74677 = (n49712 & n49745) | (n49712 & n66283) | (n49745 & n66283);
  assign n74678 = (n66230 & n74676) | (n66230 & n74677) | (n74676 & n74677);
  assign n66285 = n49710 | n49745;
  assign n74679 = n66258 | n66285;
  assign n74680 = n49712 | n66285;
  assign n74681 = (n66230 & n74679) | (n66230 & n74680) | (n74679 & n74680);
  assign n49748 = ~n74678 & n74681;
  assign n49749 = x174 & x237;
  assign n49750 = n49748 & n49749;
  assign n49751 = n49748 | n49749;
  assign n49752 = ~n49750 & n49751;
  assign n66287 = n49717 & n49752;
  assign n66288 = (n49752 & n66263) | (n49752 & n66287) | (n66263 & n66287);
  assign n66289 = n49717 | n49752;
  assign n66290 = n66263 | n66289;
  assign n49755 = ~n66288 & n66290;
  assign n49756 = x173 & x238;
  assign n49757 = n49755 & n49756;
  assign n49758 = n49755 | n49756;
  assign n49759 = ~n49757 & n49758;
  assign n66291 = n49724 & n49759;
  assign n66292 = (n49759 & n66267) | (n49759 & n66291) | (n66267 & n66291);
  assign n66293 = n49724 | n49759;
  assign n66294 = n66267 | n66293;
  assign n49762 = ~n66292 & n66294;
  assign n49763 = x172 & x239;
  assign n49764 = n49762 & n49763;
  assign n49765 = n49762 | n49763;
  assign n49766 = ~n49764 & n49765;
  assign n66295 = n49731 & n49766;
  assign n66296 = (n49766 & n66271) | (n49766 & n66295) | (n66271 & n66295);
  assign n66297 = n49731 | n49766;
  assign n66298 = n66271 | n66297;
  assign n49769 = ~n66296 & n66298;
  assign n49774 = x175 & x237;
  assign n74682 = n49745 | n74670;
  assign n74683 = (n49710 & n74670) | (n49710 & n74682) | (n74670 & n74682);
  assign n66302 = n49774 & n74683;
  assign n74684 = n49774 & n74670;
  assign n74685 = (n49745 & n49774) | (n49745 & n74684) | (n49774 & n74684);
  assign n74686 = (n66258 & n66302) | (n66258 & n74685) | (n66302 & n74685);
  assign n74687 = (n49712 & n66302) | (n49712 & n74685) | (n66302 & n74685);
  assign n74688 = (n66230 & n74686) | (n66230 & n74687) | (n74686 & n74687);
  assign n66305 = n49774 | n74683;
  assign n74689 = n49774 | n74670;
  assign n74690 = n49745 | n74689;
  assign n74691 = (n66258 & n66305) | (n66258 & n74690) | (n66305 & n74690);
  assign n74692 = (n49712 & n66305) | (n49712 & n74690) | (n66305 & n74690);
  assign n74693 = (n66230 & n74691) | (n66230 & n74692) | (n74691 & n74692);
  assign n49777 = ~n74688 & n74693;
  assign n66308 = n49750 & n49777;
  assign n74694 = (n49777 & n66287) | (n49777 & n66308) | (n66287 & n66308);
  assign n74695 = (n49752 & n49777) | (n49752 & n66308) | (n49777 & n66308);
  assign n74696 = (n66263 & n74694) | (n66263 & n74695) | (n74694 & n74695);
  assign n66310 = n49750 | n49777;
  assign n74697 = n66287 | n66310;
  assign n74698 = n49752 | n66310;
  assign n74699 = (n66263 & n74697) | (n66263 & n74698) | (n74697 & n74698);
  assign n49780 = ~n74696 & n74699;
  assign n49781 = x174 & x238;
  assign n49782 = n49780 & n49781;
  assign n49783 = n49780 | n49781;
  assign n49784 = ~n49782 & n49783;
  assign n66312 = n49757 & n49784;
  assign n66313 = (n49784 & n66292) | (n49784 & n66312) | (n66292 & n66312);
  assign n66314 = n49757 | n49784;
  assign n66315 = n66292 | n66314;
  assign n49787 = ~n66313 & n66315;
  assign n49788 = x173 & x239;
  assign n49789 = n49787 & n49788;
  assign n49790 = n49787 | n49788;
  assign n49791 = ~n49789 & n49790;
  assign n66316 = n49764 & n49791;
  assign n66317 = (n49791 & n66296) | (n49791 & n66316) | (n66296 & n66316);
  assign n66318 = n49764 | n49791;
  assign n66319 = n66296 | n66318;
  assign n49794 = ~n66317 & n66319;
  assign n49798 = x175 & x238;
  assign n74700 = n49777 | n74688;
  assign n74701 = (n49750 & n74688) | (n49750 & n74700) | (n74688 & n74700);
  assign n66323 = n49798 & n74701;
  assign n74702 = n49798 & n74688;
  assign n74703 = (n49777 & n49798) | (n49777 & n74702) | (n49798 & n74702);
  assign n74704 = (n66287 & n66323) | (n66287 & n74703) | (n66323 & n74703);
  assign n74705 = (n49752 & n66323) | (n49752 & n74703) | (n66323 & n74703);
  assign n74706 = (n66263 & n74704) | (n66263 & n74705) | (n74704 & n74705);
  assign n66326 = n49798 | n74701;
  assign n74707 = n49798 | n74688;
  assign n74708 = n49777 | n74707;
  assign n74709 = (n66287 & n66326) | (n66287 & n74708) | (n66326 & n74708);
  assign n74710 = (n49752 & n66326) | (n49752 & n74708) | (n66326 & n74708);
  assign n74711 = (n66263 & n74709) | (n66263 & n74710) | (n74709 & n74710);
  assign n49801 = ~n74706 & n74711;
  assign n66329 = n49782 & n49801;
  assign n74712 = (n49801 & n66312) | (n49801 & n66329) | (n66312 & n66329);
  assign n74713 = (n49784 & n49801) | (n49784 & n66329) | (n49801 & n66329);
  assign n74714 = (n66292 & n74712) | (n66292 & n74713) | (n74712 & n74713);
  assign n66331 = n49782 | n49801;
  assign n74715 = n66312 | n66331;
  assign n74716 = n49784 | n66331;
  assign n74717 = (n66292 & n74715) | (n66292 & n74716) | (n74715 & n74716);
  assign n49804 = ~n74714 & n74717;
  assign n49805 = x174 & x239;
  assign n49806 = n49804 & n49805;
  assign n49807 = n49804 | n49805;
  assign n49808 = ~n49806 & n49807;
  assign n66333 = n49789 & n49808;
  assign n66334 = (n49808 & n66317) | (n49808 & n66333) | (n66317 & n66333);
  assign n66335 = n49789 | n49808;
  assign n66336 = n66317 | n66335;
  assign n49811 = ~n66334 & n66336;
  assign n49814 = x175 & x239;
  assign n74718 = n49801 | n74706;
  assign n74719 = (n49782 & n74706) | (n49782 & n74718) | (n74706 & n74718);
  assign n66340 = n49814 & n74719;
  assign n74720 = n49814 & n74706;
  assign n74721 = (n49801 & n49814) | (n49801 & n74720) | (n49814 & n74720);
  assign n74722 = (n66312 & n66340) | (n66312 & n74721) | (n66340 & n74721);
  assign n74723 = (n49784 & n66340) | (n49784 & n74721) | (n66340 & n74721);
  assign n74724 = (n66292 & n74722) | (n66292 & n74723) | (n74722 & n74723);
  assign n66343 = n49814 | n74719;
  assign n74725 = n49814 | n74706;
  assign n74726 = n49801 | n74725;
  assign n74727 = (n66312 & n66343) | (n66312 & n74726) | (n66343 & n74726);
  assign n74728 = (n49784 & n66343) | (n49784 & n74726) | (n66343 & n74726);
  assign n74729 = (n66292 & n74727) | (n66292 & n74728) | (n74727 & n74728);
  assign n49817 = ~n74724 & n74729;
  assign n66346 = n49806 & n49817;
  assign n74730 = (n49817 & n66333) | (n49817 & n66346) | (n66333 & n66346);
  assign n74731 = (n49808 & n49817) | (n49808 & n66346) | (n49817 & n66346);
  assign n74732 = (n66317 & n74730) | (n66317 & n74731) | (n74730 & n74731);
  assign n66348 = n49806 | n49817;
  assign n74733 = n66333 | n66348;
  assign n74734 = n49808 | n66348;
  assign n74735 = (n66317 & n74733) | (n66317 & n74734) | (n74733 & n74734);
  assign n49820 = ~n74732 & n74735;
  assign n66351 = n49817 | n74724;
  assign n74736 = n49817 | n74724;
  assign n74737 = (n49806 & n74724) | (n49806 & n74736) | (n74724 & n74736);
  assign n74738 = (n66333 & n66351) | (n66333 & n74737) | (n66351 & n74737);
  assign n74739 = (n49808 & n66351) | (n49808 & n74737) | (n66351 & n74737);
  assign n74740 = (n66317 & n74738) | (n66317 & n74739) | (n74738 & n74739);
  assign y0 = n17;
  assign y1 = n22;
  assign y2 = n34;
  assign y3 = n54;
  assign y4 = n82;
  assign y5 = n118;
  assign y6 = n162;
  assign y7 = n214;
  assign y8 = n266;
  assign y9 = n314;
  assign y10 = n355;
  assign y11 = n388;
  assign y12 = n413;
  assign y13 = n430;
  assign y14 = n439;
  assign y15 = n723;
  assign y16 = n756;
  assign y17 = n761;
  assign y18 = n773;
  assign y19 = n793;
  assign y20 = n821;
  assign y21 = n857;
  assign y22 = n901;
  assign y23 = n953;
  assign y24 = n1013;
  assign y25 = n1081;
  assign y26 = n1157;
  assign y27 = n1241;
  assign y28 = n1333;
  assign y29 = n1433;
  assign y30 = n1541;
  assign y31 = n1657;
  assign y32 = n1773;
  assign y33 = n1885;
  assign y34 = n1990;
  assign y35 = n2087;
  assign y36 = n2176;
  assign y37 = n2257;
  assign y38 = n2330;
  assign y39 = n2395;
  assign y40 = n2452;
  assign y41 = n2501;
  assign y42 = n2542;
  assign y43 = n2575;
  assign y44 = n2600;
  assign y45 = n2617;
  assign y46 = n2626;
  assign y47 = n3882;
  assign y48 = n3947;
  assign y49 = n3952;
  assign y50 = n3964;
  assign y51 = n3984;
  assign y52 = n4012;
  assign y53 = n4048;
  assign y54 = n4092;
  assign y55 = n4144;
  assign y56 = n4204;
  assign y57 = n4272;
  assign y58 = n4348;
  assign y59 = n4432;
  assign y60 = n4524;
  assign y61 = n4624;
  assign y62 = n4732;
  assign y63 = n4848;
  assign y64 = n4972;
  assign y65 = n5104;
  assign y66 = n5244;
  assign y67 = n5392;
  assign y68 = n5548;
  assign y69 = n5712;
  assign y70 = n5884;
  assign y71 = n6064;
  assign y72 = n6252;
  assign y73 = n6448;
  assign y74 = n6652;
  assign y75 = n6864;
  assign y76 = n7084;
  assign y77 = n7312;
  assign y78 = n7548;
  assign y79 = n7792;
  assign y80 = n8036;
  assign y81 = n8276;
  assign y82 = n8509;
  assign y83 = n8734;
  assign y84 = n8951;
  assign y85 = n9160;
  assign y86 = n9361;
  assign y87 = n9554;
  assign y88 = n9739;
  assign y89 = n9916;
  assign y90 = n10085;
  assign y91 = n10246;
  assign y92 = n10399;
  assign y93 = n10544;
  assign y94 = n10681;
  assign y95 = n10810;
  assign y96 = n10931;
  assign y97 = n11044;
  assign y98 = n11149;
  assign y99 = n11246;
  assign y100 = n11335;
  assign y101 = n11416;
  assign y102 = n11489;
  assign y103 = n11554;
  assign y104 = n11611;
  assign y105 = n11660;
  assign y106 = n11701;
  assign y107 = n11734;
  assign y108 = n11759;
  assign y109 = n11776;
  assign y110 = n11785;
  assign y111 = n17629;
  assign y112 = n17758;
  assign y113 = n17763;
  assign y114 = n17775;
  assign y115 = n17795;
  assign y116 = n17823;
  assign y117 = n17859;
  assign y118 = n17903;
  assign y119 = n17955;
  assign y120 = n18015;
  assign y121 = n18083;
  assign y122 = n18159;
  assign y123 = n18243;
  assign y124 = n18335;
  assign y125 = n18435;
  assign y126 = n18543;
  assign y127 = n18659;
  assign y128 = n18783;
  assign y129 = n18915;
  assign y130 = n19055;
  assign y131 = n19203;
  assign y132 = n19359;
  assign y133 = n19523;
  assign y134 = n19695;
  assign y135 = n19875;
  assign y136 = n20063;
  assign y137 = n20259;
  assign y138 = n20463;
  assign y139 = n20675;
  assign y140 = n20895;
  assign y141 = n21123;
  assign y142 = n21359;
  assign y143 = n21603;
  assign y144 = n21855;
  assign y145 = n22115;
  assign y146 = n22383;
  assign y147 = n22659;
  assign y148 = n22943;
  assign y149 = n23235;
  assign y150 = n23535;
  assign y151 = n23843;
  assign y152 = n24159;
  assign y153 = n24483;
  assign y154 = n24815;
  assign y155 = n25155;
  assign y156 = n25503;
  assign y157 = n25859;
  assign y158 = n26223;
  assign y159 = n26595;
  assign y160 = n26975;
  assign y161 = n27363;
  assign y162 = n27759;
  assign y163 = n28163;
  assign y164 = n28575;
  assign y165 = n28995;
  assign y166 = n29423;
  assign y167 = n29859;
  assign y168 = n30303;
  assign y169 = n30755;
  assign y170 = n31215;
  assign y171 = n31683;
  assign y172 = n32159;
  assign y173 = n32643;
  assign y174 = n33135;
  assign y175 = n33635;
  assign y176 = n34135;
  assign y177 = n34631;
  assign y178 = n35120;
  assign y179 = n35601;
  assign y180 = n36074;
  assign y181 = n36539;
  assign y182 = n36996;
  assign y183 = n37445;
  assign y184 = n37886;
  assign y185 = n38319;
  assign y186 = n38744;
  assign y187 = n39161;
  assign y188 = n39570;
  assign y189 = n39971;
  assign y190 = n40364;
  assign y191 = n40749;
  assign y192 = n41126;
  assign y193 = n41495;
  assign y194 = n41856;
  assign y195 = n42209;
  assign y196 = n42554;
  assign y197 = n42891;
  assign y198 = n43220;
  assign y199 = n43541;
  assign y200 = n43854;
  assign y201 = n44159;
  assign y202 = n44456;
  assign y203 = n44745;
  assign y204 = n45026;
  assign y205 = n45299;
  assign y206 = n45564;
  assign y207 = n45821;
  assign y208 = n46070;
  assign y209 = n46311;
  assign y210 = n46544;
  assign y211 = n46769;
  assign y212 = n46986;
  assign y213 = n47195;
  assign y214 = n47396;
  assign y215 = n47589;
  assign y216 = n47774;
  assign y217 = n47951;
  assign y218 = n48120;
  assign y219 = n48281;
  assign y220 = n48434;
  assign y221 = n48579;
  assign y222 = n48716;
  assign y223 = n48845;
  assign y224 = n48966;
  assign y225 = n49079;
  assign y226 = n49184;
  assign y227 = n49281;
  assign y228 = n49370;
  assign y229 = n49451;
  assign y230 = n49524;
  assign y231 = n49589;
  assign y232 = n49646;
  assign y233 = n49695;
  assign y234 = n49736;
  assign y235 = n49769;
  assign y236 = n49794;
  assign y237 = n49811;
  assign y238 = n49820;
  assign y239 = n74740;
endmodule

